magic
tech EFS8A
magscale 1 2
timestamp 1604399536
<< locali >>
rect 2973 23035 3007 23205
rect 13277 22423 13311 22525
rect 8585 21879 8619 22049
rect 6837 16031 6871 16133
rect 17325 12631 17359 12801
rect 8125 11543 8159 11645
<< viali >>
rect 7941 25381 7975 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 3065 25313 3099 25347
rect 4721 25313 4755 25347
rect 4813 25245 4847 25279
rect 4997 25245 5031 25279
rect 6929 25245 6963 25279
rect 2421 25177 2455 25211
rect 4353 25177 4387 25211
rect 1593 25109 1627 25143
rect 2697 25109 2731 25143
rect 8401 25109 8435 25143
rect 12909 25109 12943 25143
rect 1869 24837 1903 24871
rect 2329 24837 2363 24871
rect 3065 24769 3099 24803
rect 4629 24769 4663 24803
rect 5089 24769 5123 24803
rect 6837 24769 6871 24803
rect 7757 24769 7791 24803
rect 8309 24769 8343 24803
rect 8401 24769 8435 24803
rect 12265 24769 12299 24803
rect 12909 24769 12943 24803
rect 13093 24769 13127 24803
rect 1409 24701 1443 24735
rect 2789 24701 2823 24735
rect 3525 24701 3559 24735
rect 4353 24701 4387 24735
rect 5365 24701 5399 24735
rect 5549 24701 5583 24735
rect 6193 24701 6227 24735
rect 9597 24701 9631 24735
rect 2881 24633 2915 24667
rect 3893 24633 3927 24667
rect 7389 24633 7423 24667
rect 9137 24633 9171 24667
rect 9842 24633 9876 24667
rect 11805 24633 11839 24667
rect 12817 24633 12851 24667
rect 1593 24565 1627 24599
rect 2421 24565 2455 24599
rect 3985 24565 4019 24599
rect 4445 24565 4479 24599
rect 5733 24565 5767 24599
rect 7849 24565 7883 24599
rect 8217 24565 8251 24599
rect 9413 24565 9447 24599
rect 10977 24565 11011 24599
rect 12449 24565 12483 24599
rect 2605 24361 2639 24395
rect 8033 24361 8067 24395
rect 10149 24361 10183 24395
rect 15669 24361 15703 24395
rect 17325 24361 17359 24395
rect 21833 24361 21867 24395
rect 23489 24361 23523 24395
rect 2145 24293 2179 24327
rect 2697 24293 2731 24327
rect 3249 24293 3283 24327
rect 3893 24293 3927 24327
rect 11682 24293 11716 24327
rect 5080 24225 5114 24259
rect 7941 24225 7975 24259
rect 10057 24225 10091 24259
rect 15485 24225 15519 24259
rect 17141 24225 17175 24259
rect 21649 24225 21683 24259
rect 23305 24225 23339 24259
rect 2789 24157 2823 24191
rect 4813 24157 4847 24191
rect 8217 24157 8251 24191
rect 10333 24157 10367 24191
rect 11437 24157 11471 24191
rect 6929 24089 6963 24123
rect 7573 24089 7607 24123
rect 1685 24021 1719 24055
rect 2237 24021 2271 24055
rect 4445 24021 4479 24055
rect 6193 24021 6227 24055
rect 7297 24021 7331 24055
rect 9689 24021 9723 24055
rect 10793 24021 10827 24055
rect 12817 24021 12851 24055
rect 13921 24021 13955 24055
rect 4445 23817 4479 23851
rect 4997 23817 5031 23851
rect 6469 23817 6503 23851
rect 7021 23817 7055 23851
rect 9321 23817 9355 23851
rect 9781 23817 9815 23851
rect 16497 23817 16531 23851
rect 18429 23817 18463 23851
rect 19533 23817 19567 23851
rect 20637 23817 20671 23851
rect 21741 23817 21775 23851
rect 23857 23817 23891 23851
rect 24961 23817 24995 23851
rect 8217 23749 8251 23783
rect 5641 23681 5675 23715
rect 7757 23681 7791 23715
rect 9873 23681 9907 23715
rect 2329 23613 2363 23647
rect 4905 23613 4939 23647
rect 5457 23613 5491 23647
rect 7573 23613 7607 23647
rect 7665 23613 7699 23647
rect 8585 23613 8619 23647
rect 8861 23613 8895 23647
rect 13829 23613 13863 23647
rect 16313 23613 16347 23647
rect 18245 23613 18279 23647
rect 18797 23613 18831 23647
rect 19349 23613 19383 23647
rect 20453 23613 20487 23647
rect 21005 23613 21039 23647
rect 21557 23613 21591 23647
rect 22109 23613 22143 23647
rect 23673 23613 23707 23647
rect 24777 23613 24811 23647
rect 25329 23613 25363 23647
rect 2574 23545 2608 23579
rect 5365 23545 5399 23579
rect 10140 23545 10174 23579
rect 12173 23545 12207 23579
rect 14074 23545 14108 23579
rect 15761 23545 15795 23579
rect 19901 23545 19935 23579
rect 22477 23545 22511 23579
rect 1777 23477 1811 23511
rect 2237 23477 2271 23511
rect 3709 23477 3743 23511
rect 6009 23477 6043 23511
rect 7205 23477 7239 23511
rect 11253 23477 11287 23511
rect 11805 23477 11839 23511
rect 12817 23477 12851 23511
rect 13645 23477 13679 23511
rect 15209 23477 15243 23511
rect 16129 23477 16163 23511
rect 17141 23477 17175 23511
rect 23305 23477 23339 23511
rect 24225 23477 24259 23511
rect 2513 23273 2547 23307
rect 3433 23273 3467 23307
rect 4537 23273 4571 23307
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 9505 23273 9539 23307
rect 10057 23273 10091 23307
rect 10149 23273 10183 23307
rect 13369 23273 13403 23307
rect 15485 23273 15519 23307
rect 16773 23273 16807 23307
rect 19073 23273 19107 23307
rect 21097 23273 21131 23307
rect 22385 23273 22419 23307
rect 24041 23273 24075 23307
rect 2421 23205 2455 23239
rect 2973 23205 3007 23239
rect 10701 23205 10735 23239
rect 12256 23205 12290 23239
rect 1961 23137 1995 23171
rect 2605 23069 2639 23103
rect 4629 23137 4663 23171
rect 4885 23137 4919 23171
rect 7369 23137 7403 23171
rect 11989 23137 12023 23171
rect 15301 23137 15335 23171
rect 16589 23137 16623 23171
rect 17877 23137 17911 23171
rect 18889 23137 18923 23171
rect 20913 23137 20947 23171
rect 22201 23137 22235 23171
rect 23857 23137 23891 23171
rect 7113 23069 7147 23103
rect 10241 23069 10275 23103
rect 2973 23001 3007 23035
rect 3157 23001 3191 23035
rect 18061 23001 18095 23035
rect 2053 22933 2087 22967
rect 6009 22933 6043 22967
rect 6653 22933 6687 22967
rect 9689 22933 9723 22967
rect 11069 22933 11103 22967
rect 11437 22933 11471 22967
rect 3525 22729 3559 22763
rect 4261 22729 4295 22763
rect 4629 22729 4663 22763
rect 6653 22729 6687 22763
rect 9689 22729 9723 22763
rect 11713 22729 11747 22763
rect 16497 22729 16531 22763
rect 7113 22661 7147 22695
rect 7573 22661 7607 22695
rect 11989 22661 12023 22695
rect 22753 22661 22787 22695
rect 23857 22661 23891 22695
rect 5089 22593 5123 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 7757 22593 7791 22627
rect 11069 22593 11103 22627
rect 2145 22525 2179 22559
rect 5549 22525 5583 22559
rect 10977 22525 11011 22559
rect 13277 22525 13311 22559
rect 13553 22525 13587 22559
rect 16313 22525 16347 22559
rect 16773 22525 16807 22559
rect 22569 22525 22603 22559
rect 23029 22525 23063 22559
rect 2390 22457 2424 22491
rect 8002 22457 8036 22491
rect 10425 22457 10459 22491
rect 10885 22457 10919 22491
rect 12449 22457 12483 22491
rect 13093 22457 13127 22491
rect 13820 22457 13854 22491
rect 18245 22457 18279 22491
rect 1685 22389 1719 22423
rect 2053 22389 2087 22423
rect 5181 22389 5215 22423
rect 6285 22389 6319 22423
rect 9137 22389 9171 22423
rect 10517 22389 10551 22423
rect 13277 22389 13311 22423
rect 13369 22389 13403 22423
rect 14933 22389 14967 22423
rect 15577 22389 15611 22423
rect 17233 22389 17267 22423
rect 18889 22389 18923 22423
rect 20913 22389 20947 22423
rect 22201 22389 22235 22423
rect 1685 22185 1719 22219
rect 2145 22185 2179 22219
rect 2237 22185 2271 22219
rect 4077 22185 4111 22219
rect 4721 22185 4755 22219
rect 5089 22185 5123 22219
rect 7021 22185 7055 22219
rect 7757 22185 7791 22219
rect 8033 22185 8067 22219
rect 9781 22185 9815 22219
rect 10793 22185 10827 22219
rect 13001 22185 13035 22219
rect 5457 22117 5491 22151
rect 10609 22117 10643 22151
rect 11161 22117 11195 22151
rect 2881 22049 2915 22083
rect 8217 22049 8251 22083
rect 8585 22049 8619 22083
rect 9505 22049 9539 22083
rect 11253 22049 11287 22083
rect 12173 22049 12207 22083
rect 13093 22049 13127 22083
rect 2421 21981 2455 22015
rect 5549 21981 5583 22015
rect 5733 21981 5767 22015
rect 7113 21981 7147 22015
rect 7205 21981 7239 22015
rect 3709 21913 3743 21947
rect 6561 21913 6595 21947
rect 9137 21981 9171 22015
rect 11345 21981 11379 22015
rect 12449 21981 12483 22015
rect 13277 21981 13311 22015
rect 1777 21845 1811 21879
rect 3341 21845 3375 21879
rect 6193 21845 6227 21879
rect 6653 21845 6687 21879
rect 8401 21845 8435 21879
rect 8585 21845 8619 21879
rect 8769 21845 8803 21879
rect 12633 21845 12667 21879
rect 13645 21845 13679 21879
rect 1593 21641 1627 21675
rect 2053 21641 2087 21675
rect 4537 21641 4571 21675
rect 6101 21641 6135 21675
rect 6561 21641 6595 21675
rect 6837 21641 6871 21675
rect 8585 21641 8619 21675
rect 10885 21641 10919 21675
rect 11621 21641 11655 21675
rect 12265 21641 12299 21675
rect 14381 21641 14415 21675
rect 3157 21505 3191 21539
rect 3709 21505 3743 21539
rect 3893 21505 3927 21539
rect 5549 21505 5583 21539
rect 7297 21505 7331 21539
rect 7481 21505 7515 21539
rect 8677 21505 8711 21539
rect 1409 21437 1443 21471
rect 2789 21437 2823 21471
rect 4905 21437 4939 21471
rect 5457 21437 5491 21471
rect 7205 21437 7239 21471
rect 7849 21437 7883 21471
rect 8944 21437 8978 21471
rect 11161 21437 11195 21471
rect 13001 21437 13035 21471
rect 13268 21437 13302 21471
rect 2421 21369 2455 21403
rect 5365 21369 5399 21403
rect 3249 21301 3283 21335
rect 3617 21301 3651 21335
rect 4997 21301 5031 21335
rect 10057 21301 10091 21335
rect 11345 21301 11379 21335
rect 12817 21301 12851 21335
rect 1593 21097 1627 21131
rect 1961 21097 1995 21131
rect 3801 21097 3835 21131
rect 6377 21097 6411 21131
rect 9045 21097 9079 21131
rect 10149 21097 10183 21131
rect 11253 21097 11287 21131
rect 13829 21097 13863 21131
rect 6009 21029 6043 21063
rect 6806 21029 6840 21063
rect 8769 21029 8803 21063
rect 1409 20961 1443 20995
rect 2513 20961 2547 20995
rect 3157 20961 3191 20995
rect 4077 20961 4111 20995
rect 4344 20961 4378 20995
rect 10057 20961 10091 20995
rect 12716 20961 12750 20995
rect 6561 20893 6595 20927
rect 9505 20893 9539 20927
rect 10241 20893 10275 20927
rect 11437 20893 11471 20927
rect 12449 20893 12483 20927
rect 2697 20825 2731 20859
rect 3433 20825 3467 20859
rect 11989 20825 12023 20859
rect 12265 20825 12299 20859
rect 2329 20757 2363 20791
rect 5457 20757 5491 20791
rect 7941 20757 7975 20791
rect 9689 20757 9723 20791
rect 10885 20757 10919 20791
rect 14381 20757 14415 20791
rect 1593 20553 1627 20587
rect 3341 20553 3375 20587
rect 3985 20553 4019 20587
rect 5825 20553 5859 20587
rect 6285 20553 6319 20587
rect 6653 20553 6687 20587
rect 7941 20553 7975 20587
rect 10057 20553 10091 20587
rect 13829 20553 13863 20587
rect 10425 20485 10459 20519
rect 12449 20485 12483 20519
rect 1961 20417 1995 20451
rect 4353 20417 4387 20451
rect 5089 20417 5123 20451
rect 8033 20417 8067 20451
rect 11253 20417 11287 20451
rect 11345 20417 11379 20451
rect 12265 20417 12299 20451
rect 12909 20417 12943 20451
rect 13093 20417 13127 20451
rect 14565 20417 14599 20451
rect 2228 20349 2262 20383
rect 4813 20349 4847 20383
rect 4905 20349 4939 20383
rect 7021 20349 7055 20383
rect 8300 20349 8334 20383
rect 11161 20349 11195 20383
rect 14473 20349 14507 20383
rect 5549 20281 5583 20315
rect 7573 20281 7607 20315
rect 11897 20281 11931 20315
rect 12817 20281 12851 20315
rect 14381 20281 14415 20315
rect 4445 20213 4479 20247
rect 7205 20213 7239 20247
rect 9413 20213 9447 20247
rect 10793 20213 10827 20247
rect 13553 20213 13587 20247
rect 14013 20213 14047 20247
rect 2881 20009 2915 20043
rect 3433 20009 3467 20043
rect 4537 20009 4571 20043
rect 6561 20009 6595 20043
rect 8125 20009 8159 20043
rect 9321 20009 9355 20043
rect 10057 20009 10091 20043
rect 10885 20009 10919 20043
rect 13461 20009 13495 20043
rect 14013 20009 14047 20043
rect 5273 19941 5307 19975
rect 6990 19941 7024 19975
rect 10149 19941 10183 19975
rect 11253 19941 11287 19975
rect 11989 19941 12023 19975
rect 12326 19941 12360 19975
rect 1501 19873 1535 19907
rect 1768 19873 1802 19907
rect 5181 19873 5215 19907
rect 6745 19873 6779 19907
rect 5365 19805 5399 19839
rect 10241 19805 10275 19839
rect 12081 19805 12115 19839
rect 15301 19805 15335 19839
rect 8677 19737 8711 19771
rect 3801 19669 3835 19703
rect 4813 19669 4847 19703
rect 5825 19669 5859 19703
rect 6193 19669 6227 19703
rect 9689 19669 9723 19703
rect 14473 19669 14507 19703
rect 2605 19465 2639 19499
rect 3157 19465 3191 19499
rect 12449 19465 12483 19499
rect 3065 19397 3099 19431
rect 6837 19397 6871 19431
rect 2237 19329 2271 19363
rect 3617 19329 3651 19363
rect 3709 19329 3743 19363
rect 5457 19329 5491 19363
rect 7389 19329 7423 19363
rect 7849 19329 7883 19363
rect 13093 19329 13127 19363
rect 14749 19329 14783 19363
rect 2053 19261 2087 19295
rect 3525 19261 3559 19295
rect 5181 19261 5215 19295
rect 5273 19261 5307 19295
rect 6285 19261 6319 19295
rect 7205 19261 7239 19295
rect 9045 19261 9079 19295
rect 9229 19261 9263 19295
rect 11161 19261 11195 19295
rect 11805 19261 11839 19295
rect 12909 19261 12943 19295
rect 23673 19261 23707 19295
rect 24133 19261 24167 19295
rect 1961 19193 1995 19227
rect 4353 19193 4387 19227
rect 5917 19193 5951 19227
rect 6653 19193 6687 19227
rect 9474 19193 9508 19227
rect 12265 19193 12299 19227
rect 14105 19193 14139 19227
rect 14565 19193 14599 19227
rect 1593 19125 1627 19159
rect 4629 19125 4663 19159
rect 4813 19125 4847 19159
rect 7297 19125 7331 19159
rect 8769 19125 8803 19159
rect 10609 19125 10643 19159
rect 12817 19125 12851 19159
rect 13461 19125 13495 19159
rect 14197 19125 14231 19159
rect 14657 19125 14691 19159
rect 15761 19125 15795 19159
rect 23857 19125 23891 19159
rect 1777 18921 1811 18955
rect 2145 18921 2179 18955
rect 3525 18921 3559 18955
rect 4905 18921 4939 18955
rect 8125 18921 8159 18955
rect 10149 18921 10183 18955
rect 11253 18921 11287 18955
rect 13093 18921 13127 18955
rect 14197 18921 14231 18955
rect 16681 18921 16715 18955
rect 2881 18853 2915 18887
rect 5448 18853 5482 18887
rect 10057 18853 10091 18887
rect 10885 18853 10919 18887
rect 15546 18853 15580 18887
rect 4077 18785 4111 18819
rect 7573 18785 7607 18819
rect 8033 18785 8067 18819
rect 11621 18785 11655 18819
rect 11980 18785 12014 18819
rect 2237 18717 2271 18751
rect 2421 18717 2455 18751
rect 5181 18717 5215 18751
rect 8309 18717 8343 18751
rect 10333 18717 10367 18751
rect 11713 18717 11747 18751
rect 15301 18717 15335 18751
rect 3157 18649 3191 18683
rect 7113 18649 7147 18683
rect 7665 18649 7699 18683
rect 9689 18649 9723 18683
rect 1685 18581 1719 18615
rect 4261 18581 4295 18615
rect 6561 18581 6595 18615
rect 9229 18581 9263 18615
rect 14657 18581 14691 18615
rect 2053 18377 2087 18411
rect 3617 18377 3651 18411
rect 4261 18377 4295 18411
rect 6101 18377 6135 18411
rect 8217 18377 8251 18411
rect 9137 18377 9171 18411
rect 10241 18377 10275 18411
rect 12265 18377 12299 18411
rect 15117 18377 15151 18411
rect 16037 18377 16071 18411
rect 1777 18309 1811 18343
rect 8861 18309 8895 18343
rect 15669 18309 15703 18343
rect 2237 18241 2271 18275
rect 5181 18241 5215 18275
rect 5365 18241 5399 18275
rect 11253 18241 11287 18275
rect 11437 18241 11471 18275
rect 2504 18173 2538 18207
rect 6837 18173 6871 18207
rect 9321 18173 9355 18207
rect 9873 18173 9907 18207
rect 13737 18173 13771 18207
rect 16221 18173 16255 18207
rect 16773 18173 16807 18207
rect 4629 18105 4663 18139
rect 7082 18105 7116 18139
rect 10701 18105 10735 18139
rect 11161 18105 11195 18139
rect 12449 18105 12483 18139
rect 14004 18105 14038 18139
rect 4721 18037 4755 18071
rect 5089 18037 5123 18071
rect 5825 18037 5859 18071
rect 6561 18037 6595 18071
rect 9505 18037 9539 18071
rect 10793 18037 10827 18071
rect 11897 18037 11931 18071
rect 13553 18037 13587 18071
rect 16405 18037 16439 18071
rect 2237 17833 2271 17867
rect 3249 17833 3283 17867
rect 3893 17833 3927 17867
rect 6101 17833 6135 17867
rect 7573 17833 7607 17867
rect 7757 17833 7791 17867
rect 10241 17833 10275 17867
rect 14381 17833 14415 17867
rect 15301 17833 15335 17867
rect 1869 17765 1903 17799
rect 2697 17765 2731 17799
rect 7297 17765 7331 17799
rect 11038 17765 11072 17799
rect 2605 17697 2639 17731
rect 4988 17697 5022 17731
rect 8125 17697 8159 17731
rect 9689 17697 9723 17731
rect 14197 17697 14231 17731
rect 15669 17697 15703 17731
rect 16865 17697 16899 17731
rect 17877 17697 17911 17731
rect 2881 17629 2915 17663
rect 4721 17629 4755 17663
rect 8217 17629 8251 17663
rect 8401 17629 8435 17663
rect 10793 17629 10827 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 13829 17561 13863 17595
rect 4353 17493 4387 17527
rect 6929 17493 6963 17527
rect 8769 17493 8803 17527
rect 9873 17493 9907 17527
rect 12173 17493 12207 17527
rect 15025 17493 15059 17527
rect 17049 17493 17083 17527
rect 1593 17289 1627 17323
rect 2697 17289 2731 17323
rect 3157 17289 3191 17323
rect 3893 17289 3927 17323
rect 4261 17289 4295 17323
rect 7481 17289 7515 17323
rect 7665 17289 7699 17323
rect 10609 17289 10643 17323
rect 13921 17289 13955 17323
rect 14197 17289 14231 17323
rect 16405 17289 16439 17323
rect 16957 17289 16991 17323
rect 2329 17221 2363 17255
rect 5733 17221 5767 17255
rect 8677 17221 8711 17255
rect 9137 17221 9171 17255
rect 12449 17221 12483 17255
rect 14565 17221 14599 17255
rect 18245 17221 18279 17255
rect 4813 17153 4847 17187
rect 4905 17153 4939 17187
rect 7205 17153 7239 17187
rect 8217 17153 8251 17187
rect 9229 17153 9263 17187
rect 13093 17153 13127 17187
rect 1409 17085 1443 17119
rect 2513 17085 2547 17119
rect 3433 17085 3467 17119
rect 4721 17085 4755 17119
rect 6101 17085 6135 17119
rect 8125 17085 8159 17119
rect 9496 17085 9530 17119
rect 12909 17085 12943 17119
rect 14013 17085 14047 17119
rect 15025 17085 15059 17119
rect 18061 17085 18095 17119
rect 18521 17085 18555 17119
rect 6653 17017 6687 17051
rect 8033 17017 8067 17051
rect 12265 17017 12299 17051
rect 12817 17017 12851 17051
rect 13461 17017 13495 17051
rect 15292 17017 15326 17051
rect 4353 16949 4387 16983
rect 5365 16949 5399 16983
rect 11253 16949 11287 16983
rect 11805 16949 11839 16983
rect 14841 16949 14875 16983
rect 1593 16745 1627 16779
rect 2697 16745 2731 16779
rect 3157 16745 3191 16779
rect 3617 16745 3651 16779
rect 4077 16745 4111 16779
rect 5089 16745 5123 16779
rect 6377 16745 6411 16779
rect 8033 16745 8067 16779
rect 9321 16745 9355 16779
rect 9873 16745 9907 16779
rect 10701 16745 10735 16779
rect 12173 16745 12207 16779
rect 12817 16745 12851 16779
rect 13461 16745 13495 16779
rect 15485 16745 15519 16779
rect 15853 16745 15887 16779
rect 17969 16745 18003 16779
rect 6009 16677 6043 16711
rect 6929 16677 6963 16711
rect 7849 16677 7883 16711
rect 8493 16677 8527 16711
rect 11038 16677 11072 16711
rect 15117 16677 15151 16711
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 4445 16609 4479 16643
rect 4537 16609 4571 16643
rect 5641 16609 5675 16643
rect 6837 16609 6871 16643
rect 8401 16609 8435 16643
rect 9689 16609 9723 16643
rect 10241 16609 10275 16643
rect 13829 16609 13863 16643
rect 14565 16609 14599 16643
rect 15301 16609 15335 16643
rect 16856 16609 16890 16643
rect 2329 16541 2363 16575
rect 4629 16541 4663 16575
rect 7021 16541 7055 16575
rect 8677 16541 8711 16575
rect 10793 16541 10827 16575
rect 13921 16541 13955 16575
rect 14105 16541 14139 16575
rect 16589 16541 16623 16575
rect 6469 16405 6503 16439
rect 13369 16405 13403 16439
rect 1593 16201 1627 16235
rect 6561 16201 6595 16235
rect 6929 16201 6963 16235
rect 8033 16201 8067 16235
rect 9045 16201 9079 16235
rect 11253 16201 11287 16235
rect 15577 16201 15611 16235
rect 16589 16201 16623 16235
rect 2973 16133 3007 16167
rect 6837 16133 6871 16167
rect 11621 16133 11655 16167
rect 16221 16133 16255 16167
rect 18245 16133 18279 16167
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 3709 16065 3743 16099
rect 5733 16065 5767 16099
rect 6285 16065 6319 16099
rect 7573 16065 7607 16099
rect 8493 16065 8527 16099
rect 9413 16065 9447 16099
rect 10057 16065 10091 16099
rect 13001 16065 13035 16099
rect 16681 16065 16715 16099
rect 2697 15997 2731 16031
rect 3525 15997 3559 16031
rect 5641 15997 5675 16031
rect 6837 15997 6871 16031
rect 7389 15997 7423 16031
rect 9873 15997 9907 16031
rect 11069 15997 11103 16031
rect 12265 15997 12299 16031
rect 12817 15997 12851 16031
rect 14197 15997 14231 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 19073 15997 19107 16031
rect 19533 15997 19567 16031
rect 1961 15929 1995 15963
rect 3617 15929 3651 15963
rect 5089 15929 5123 15963
rect 9965 15929 9999 15963
rect 14464 15929 14498 15963
rect 3157 15861 3191 15895
rect 4169 15861 4203 15895
rect 4629 15861 4663 15895
rect 5181 15861 5215 15895
rect 5549 15861 5583 15895
rect 7297 15861 7331 15895
rect 9505 15861 9539 15895
rect 10793 15861 10827 15895
rect 12449 15861 12483 15895
rect 12909 15861 12943 15895
rect 13553 15861 13587 15895
rect 14013 15861 14047 15895
rect 17141 15861 17175 15895
rect 19257 15861 19291 15895
rect 2881 15657 2915 15691
rect 3893 15657 3927 15691
rect 6929 15657 6963 15691
rect 7113 15657 7147 15691
rect 8493 15657 8527 15691
rect 9873 15657 9907 15691
rect 12541 15657 12575 15691
rect 12909 15657 12943 15691
rect 13277 15657 13311 15691
rect 15485 15657 15519 15691
rect 17693 15657 17727 15691
rect 21097 15657 21131 15691
rect 7481 15589 7515 15623
rect 10670 15589 10704 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 4896 15521 4930 15555
rect 8217 15521 8251 15555
rect 13737 15521 13771 15555
rect 15301 15521 15335 15555
rect 16580 15521 16614 15555
rect 20913 15521 20947 15555
rect 4629 15453 4663 15487
rect 7573 15453 7607 15487
rect 7757 15453 7791 15487
rect 10425 15453 10459 15487
rect 13829 15453 13863 15487
rect 14013 15453 14047 15487
rect 16313 15453 16347 15487
rect 3525 15385 3559 15419
rect 6653 15385 6687 15419
rect 11805 15385 11839 15419
rect 4353 15317 4387 15351
rect 6009 15317 6043 15351
rect 9137 15317 9171 15351
rect 9505 15317 9539 15351
rect 10333 15317 10367 15351
rect 13369 15317 13403 15351
rect 14381 15317 14415 15351
rect 1593 15113 1627 15147
rect 1961 15113 1995 15147
rect 4261 15113 4295 15147
rect 8217 15113 8251 15147
rect 11161 15113 11195 15147
rect 12817 15113 12851 15147
rect 2697 15045 2731 15079
rect 4813 15045 4847 15079
rect 6653 15045 6687 15079
rect 19625 15045 19659 15079
rect 20913 15045 20947 15079
rect 2881 14977 2915 15011
rect 6837 14977 6871 15011
rect 16957 14977 16991 15011
rect 17417 14977 17451 15011
rect 1409 14909 1443 14943
rect 3148 14909 3182 14943
rect 5365 14909 5399 14943
rect 9781 14909 9815 14943
rect 13921 14909 13955 14943
rect 16221 14909 16255 14943
rect 19441 14909 19475 14943
rect 19901 14909 19935 14943
rect 7104 14841 7138 14875
rect 9321 14841 9355 14875
rect 10026 14841 10060 14875
rect 13369 14841 13403 14875
rect 14188 14841 14222 14875
rect 15945 14841 15979 14875
rect 16773 14841 16807 14875
rect 2329 14773 2363 14807
rect 5273 14773 5307 14807
rect 5549 14773 5583 14807
rect 6193 14773 6227 14807
rect 8861 14773 8895 14807
rect 9689 14773 9723 14807
rect 12909 14773 12943 14807
rect 13737 14773 13771 14807
rect 15301 14773 15335 14807
rect 16405 14773 16439 14807
rect 16865 14773 16899 14807
rect 17785 14773 17819 14807
rect 1961 14569 1995 14603
rect 2421 14569 2455 14603
rect 3525 14569 3559 14603
rect 4077 14569 4111 14603
rect 4537 14569 4571 14603
rect 6009 14569 6043 14603
rect 7481 14569 7515 14603
rect 8401 14569 8435 14603
rect 9045 14569 9079 14603
rect 10793 14569 10827 14603
rect 11069 14569 11103 14603
rect 11621 14569 11655 14603
rect 13645 14569 13679 14603
rect 14105 14569 14139 14603
rect 15485 14569 15519 14603
rect 15945 14569 15979 14603
rect 17509 14569 17543 14603
rect 1409 14501 1443 14535
rect 6368 14501 6402 14535
rect 12081 14501 12115 14535
rect 16405 14501 16439 14535
rect 2789 14433 2823 14467
rect 3893 14433 3927 14467
rect 4445 14433 4479 14467
rect 6101 14433 6135 14467
rect 10057 14433 10091 14467
rect 10149 14433 10183 14467
rect 11989 14433 12023 14467
rect 14013 14433 14047 14467
rect 16313 14433 16347 14467
rect 2881 14365 2915 14399
rect 2973 14365 3007 14399
rect 4629 14365 4663 14399
rect 8033 14365 8067 14399
rect 8585 14365 8619 14399
rect 10333 14365 10367 14399
rect 12265 14365 12299 14399
rect 13369 14365 13403 14399
rect 14197 14365 14231 14399
rect 16589 14365 16623 14399
rect 16957 14365 16991 14399
rect 5549 14297 5583 14331
rect 9505 14297 9539 14331
rect 2237 14229 2271 14263
rect 5273 14229 5307 14263
rect 9689 14229 9723 14263
rect 2605 14025 2639 14059
rect 3157 14025 3191 14059
rect 4169 14025 4203 14059
rect 4629 14025 4663 14059
rect 6193 14025 6227 14059
rect 7113 14025 7147 14059
rect 9045 14025 9079 14059
rect 10517 14025 10551 14059
rect 11989 14025 12023 14059
rect 13185 14025 13219 14059
rect 16405 14025 16439 14059
rect 16681 14025 16715 14059
rect 7573 13957 7607 13991
rect 2053 13889 2087 13923
rect 2237 13889 2271 13923
rect 3709 13889 3743 13923
rect 5089 13889 5123 13923
rect 5733 13889 5767 13923
rect 8125 13889 8159 13923
rect 8677 13889 8711 13923
rect 11161 13889 11195 13923
rect 1961 13821 1995 13855
rect 3065 13821 3099 13855
rect 3617 13821 3651 13855
rect 7389 13821 7423 13855
rect 8033 13821 8067 13855
rect 9137 13821 9171 13855
rect 9404 13821 9438 13855
rect 11621 13821 11655 13855
rect 13737 13821 13771 13855
rect 15945 13821 15979 13855
rect 3525 13753 3559 13787
rect 5641 13753 5675 13787
rect 7941 13753 7975 13787
rect 12449 13753 12483 13787
rect 14004 13753 14038 13787
rect 1593 13685 1627 13719
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 6561 13685 6595 13719
rect 13553 13685 13587 13719
rect 15117 13685 15151 13719
rect 3249 13481 3283 13515
rect 4445 13481 4479 13515
rect 6929 13481 6963 13515
rect 8125 13481 8159 13515
rect 9137 13481 9171 13515
rect 10057 13481 10091 13515
rect 13185 13481 13219 13515
rect 13829 13481 13863 13515
rect 14473 13481 14507 13515
rect 16957 13481 16991 13515
rect 21097 13481 21131 13515
rect 1685 13413 1719 13447
rect 2053 13413 2087 13447
rect 2605 13413 2639 13447
rect 4537 13413 4571 13447
rect 5825 13413 5859 13447
rect 6285 13413 6319 13447
rect 9413 13413 9447 13447
rect 11713 13413 11747 13447
rect 12072 13413 12106 13447
rect 2513 13345 2547 13379
rect 5457 13345 5491 13379
rect 7481 13345 7515 13379
rect 10149 13345 10183 13379
rect 15844 13345 15878 13379
rect 18328 13345 18362 13379
rect 20913 13345 20947 13379
rect 2697 13277 2731 13311
rect 4629 13277 4663 13311
rect 6377 13277 6411 13311
rect 6469 13277 6503 13311
rect 8585 13277 8619 13311
rect 10241 13277 10275 13311
rect 11805 13277 11839 13311
rect 14197 13277 14231 13311
rect 15577 13277 15611 13311
rect 18061 13277 18095 13311
rect 3893 13209 3927 13243
rect 5917 13209 5951 13243
rect 7665 13209 7699 13243
rect 9689 13209 9723 13243
rect 19441 13209 19475 13243
rect 2145 13141 2179 13175
rect 4077 13141 4111 13175
rect 7297 13141 7331 13175
rect 8493 13141 8527 13175
rect 14933 13141 14967 13175
rect 2513 12937 2547 12971
rect 3985 12937 4019 12971
rect 5181 12937 5215 12971
rect 6285 12937 6319 12971
rect 8769 12937 8803 12971
rect 9137 12937 9171 12971
rect 9321 12937 9355 12971
rect 10333 12937 10367 12971
rect 11253 12937 11287 12971
rect 11529 12937 11563 12971
rect 16405 12937 16439 12971
rect 20913 12937 20947 12971
rect 22477 12937 22511 12971
rect 10885 12869 10919 12903
rect 13829 12869 13863 12903
rect 15117 12869 15151 12903
rect 2605 12801 2639 12835
rect 4629 12801 4663 12835
rect 5825 12801 5859 12835
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 9781 12801 9815 12835
rect 9965 12801 9999 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 1409 12733 1443 12767
rect 5549 12733 5583 12767
rect 7093 12733 7127 12767
rect 9689 12733 9723 12767
rect 11337 12733 11371 12767
rect 12449 12733 12483 12767
rect 14933 12733 14967 12767
rect 16313 12733 16347 12767
rect 16773 12733 16807 12767
rect 2145 12665 2179 12699
rect 2850 12665 2884 12699
rect 12694 12665 12728 12699
rect 15577 12665 15611 12699
rect 18061 12733 18095 12767
rect 22293 12733 22327 12767
rect 22753 12733 22787 12767
rect 18521 12665 18555 12699
rect 1593 12597 1627 12631
rect 4997 12597 5031 12631
rect 5641 12597 5675 12631
rect 8217 12597 8251 12631
rect 11897 12597 11931 12631
rect 12265 12597 12299 12631
rect 14841 12597 14875 12631
rect 16865 12597 16899 12631
rect 17325 12597 17359 12631
rect 17509 12597 17543 12631
rect 18981 12597 19015 12631
rect 1685 12393 1719 12427
rect 3893 12393 3927 12427
rect 4261 12393 4295 12427
rect 4721 12393 4755 12427
rect 6837 12393 6871 12427
rect 9413 12393 9447 12427
rect 9689 12393 9723 12427
rect 11253 12393 11287 12427
rect 11621 12393 11655 12427
rect 12541 12393 12575 12427
rect 19165 12393 19199 12427
rect 22017 12393 22051 12427
rect 2789 12325 2823 12359
rect 15546 12325 15580 12359
rect 2145 12257 2179 12291
rect 2237 12257 2271 12291
rect 4077 12257 4111 12291
rect 5724 12257 5758 12291
rect 8309 12257 8343 12291
rect 10057 12257 10091 12291
rect 10149 12257 10183 12291
rect 11713 12257 11747 12291
rect 14013 12257 14047 12291
rect 17785 12257 17819 12291
rect 18052 12257 18086 12291
rect 21833 12257 21867 12291
rect 2329 12189 2363 12223
rect 5457 12189 5491 12223
rect 8401 12189 8435 12223
rect 8585 12189 8619 12223
rect 8953 12189 8987 12223
rect 10333 12189 10367 12223
rect 11805 12189 11839 12223
rect 14105 12189 14139 12223
rect 14289 12189 14323 12223
rect 15301 12189 15335 12223
rect 1777 12121 1811 12155
rect 16681 12121 16715 12155
rect 3157 12053 3191 12087
rect 5181 12053 5215 12087
rect 7481 12053 7515 12087
rect 7941 12053 7975 12087
rect 13093 12053 13127 12087
rect 13461 12053 13495 12087
rect 13645 12053 13679 12087
rect 14749 12053 14783 12087
rect 17233 12053 17267 12087
rect 1685 11849 1719 11883
rect 3525 11849 3559 11883
rect 5181 11849 5215 11883
rect 6285 11849 6319 11883
rect 7941 11849 7975 11883
rect 10793 11849 10827 11883
rect 11253 11849 11287 11883
rect 15301 11849 15335 11883
rect 16037 11849 16071 11883
rect 17785 11849 17819 11883
rect 21373 11849 21407 11883
rect 1961 11781 1995 11815
rect 2145 11713 2179 11747
rect 4721 11713 4755 11747
rect 5825 11713 5859 11747
rect 6561 11713 6595 11747
rect 7389 11713 7423 11747
rect 16497 11713 16531 11747
rect 16681 11713 16715 11747
rect 18521 11713 18555 11747
rect 2412 11645 2446 11679
rect 8125 11645 8159 11679
rect 8401 11645 8435 11679
rect 8668 11645 8702 11679
rect 12173 11645 12207 11679
rect 13185 11645 13219 11679
rect 13369 11645 13403 11679
rect 13625 11645 13659 11679
rect 21189 11645 21223 11679
rect 21649 11645 21683 11679
rect 4077 11577 4111 11611
rect 4997 11577 5031 11611
rect 5641 11577 5675 11611
rect 7297 11577 7331 11611
rect 11345 11577 11379 11611
rect 18061 11577 18095 11611
rect 5549 11509 5583 11543
rect 8125 11509 8159 11543
rect 8217 11509 8251 11543
rect 9781 11509 9815 11543
rect 10333 11509 10367 11543
rect 11805 11509 11839 11543
rect 12909 11509 12943 11543
rect 14749 11509 14783 11543
rect 15853 11509 15887 11543
rect 16405 11509 16439 11543
rect 17141 11509 17175 11543
rect 22017 11509 22051 11543
rect 1961 11305 1995 11339
rect 2881 11305 2915 11339
rect 3801 11305 3835 11339
rect 5273 11305 5307 11339
rect 5641 11305 5675 11339
rect 6101 11305 6135 11339
rect 6929 11305 6963 11339
rect 8493 11305 8527 11339
rect 9873 11305 9907 11339
rect 13277 11305 13311 11339
rect 13737 11305 13771 11339
rect 14473 11305 14507 11339
rect 15301 11305 15335 11339
rect 16405 11305 16439 11339
rect 17785 11305 17819 11339
rect 7380 11237 7414 11271
rect 11152 11237 11186 11271
rect 2329 11169 2363 11203
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 4537 11169 4571 11203
rect 6469 11169 6503 11203
rect 10425 11169 10459 11203
rect 15669 11169 15703 11203
rect 17601 11169 17635 11203
rect 1409 11101 1443 11135
rect 3065 11101 3099 11135
rect 3433 11101 3467 11135
rect 4629 11101 4663 11135
rect 7113 11101 7147 11135
rect 10885 11101 10919 11135
rect 13829 11101 13863 11135
rect 13921 11101 13955 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 4077 11033 4111 11067
rect 13369 11033 13403 11067
rect 15117 11033 15151 11067
rect 2421 10965 2455 10999
rect 12265 10965 12299 10999
rect 12817 10965 12851 10999
rect 3065 10761 3099 10795
rect 3709 10761 3743 10795
rect 6837 10761 6871 10795
rect 8309 10761 8343 10795
rect 11069 10761 11103 10795
rect 13829 10761 13863 10795
rect 15209 10761 15243 10795
rect 16589 10761 16623 10795
rect 16957 10761 16991 10795
rect 18521 10761 18555 10795
rect 6285 10693 6319 10727
rect 1685 10625 1719 10659
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 14657 10625 14691 10659
rect 15853 10625 15887 10659
rect 16221 10625 16255 10659
rect 4077 10557 4111 10591
rect 4169 10557 4203 10591
rect 4425 10557 4459 10591
rect 7849 10557 7883 10591
rect 9505 10557 9539 10591
rect 9689 10557 9723 10591
rect 11621 10557 11655 10591
rect 12173 10557 12207 10591
rect 12449 10557 12483 10591
rect 16773 10557 16807 10591
rect 17233 10557 17267 10591
rect 18337 10557 18371 10591
rect 18889 10557 18923 10591
rect 1952 10489 1986 10523
rect 9229 10489 9263 10523
rect 9956 10489 9990 10523
rect 12694 10489 12728 10523
rect 15669 10489 15703 10523
rect 5549 10421 5583 10455
rect 6561 10421 6595 10455
rect 7205 10421 7239 10455
rect 15025 10421 15059 10455
rect 15577 10421 15611 10455
rect 17601 10421 17635 10455
rect 1869 10217 1903 10251
rect 2789 10217 2823 10251
rect 3801 10217 3835 10251
rect 4537 10217 4571 10251
rect 7205 10217 7239 10251
rect 7665 10217 7699 10251
rect 8125 10217 8159 10251
rect 9689 10217 9723 10251
rect 11253 10217 11287 10251
rect 13553 10217 13587 10251
rect 15117 10217 15151 10251
rect 15577 10217 15611 10251
rect 17141 10217 17175 10251
rect 1777 10149 1811 10183
rect 2513 10149 2547 10183
rect 3525 10149 3559 10183
rect 5426 10149 5460 10183
rect 11713 10149 11747 10183
rect 13461 10149 13495 10183
rect 14013 10149 14047 10183
rect 16028 10149 16062 10183
rect 2973 10081 3007 10115
rect 8033 10081 8067 10115
rect 8677 10081 8711 10115
rect 10057 10081 10091 10115
rect 10977 10081 11011 10115
rect 11621 10081 11655 10115
rect 13921 10081 13955 10115
rect 15761 10081 15795 10115
rect 1961 10013 1995 10047
rect 4077 10013 4111 10047
rect 5181 10013 5215 10047
rect 8217 10013 8251 10047
rect 10149 10013 10183 10047
rect 10333 10013 10367 10047
rect 11897 10013 11931 10047
rect 14105 10013 14139 10047
rect 1409 9945 1443 9979
rect 4905 9945 4939 9979
rect 7573 9945 7607 9979
rect 13093 9945 13127 9979
rect 14565 9945 14599 9979
rect 3157 9877 3191 9911
rect 6561 9877 6595 9911
rect 12541 9877 12575 9911
rect 1961 9673 1995 9707
rect 3525 9673 3559 9707
rect 3893 9673 3927 9707
rect 5365 9673 5399 9707
rect 8217 9673 8251 9707
rect 11069 9673 11103 9707
rect 12081 9673 12115 9707
rect 14013 9673 14047 9707
rect 15853 9673 15887 9707
rect 17141 9673 17175 9707
rect 18245 9673 18279 9707
rect 1593 9605 1627 9639
rect 2329 9605 2363 9639
rect 2697 9605 2731 9639
rect 9689 9605 9723 9639
rect 16405 9605 16439 9639
rect 10333 9537 10367 9571
rect 13001 9537 13035 9571
rect 1409 9469 1443 9503
rect 2505 9469 2539 9503
rect 3985 9469 4019 9503
rect 4241 9469 4275 9503
rect 6009 9469 6043 9503
rect 6653 9469 6687 9503
rect 6837 9469 6871 9503
rect 12817 9469 12851 9503
rect 14473 9469 14507 9503
rect 14729 9469 14763 9503
rect 16957 9469 16991 9503
rect 17417 9469 17451 9503
rect 18061 9469 18095 9503
rect 18521 9469 18555 9503
rect 3065 9401 3099 9435
rect 7082 9401 7116 9435
rect 8861 9401 8895 9435
rect 10057 9401 10091 9435
rect 11253 9401 11287 9435
rect 14381 9401 14415 9435
rect 9137 9333 9171 9367
rect 9505 9333 9539 9367
rect 10149 9333 10183 9367
rect 10701 9333 10735 9367
rect 11713 9333 11747 9367
rect 12449 9333 12483 9367
rect 12909 9333 12943 9367
rect 13553 9333 13587 9367
rect 1869 9129 1903 9163
rect 2329 9129 2363 9163
rect 2605 9129 2639 9163
rect 3341 9129 3375 9163
rect 3893 9129 3927 9163
rect 4077 9129 4111 9163
rect 4445 9129 4479 9163
rect 4537 9129 4571 9163
rect 5273 9129 5307 9163
rect 7757 9129 7791 9163
rect 9505 9129 9539 9163
rect 11989 9129 12023 9163
rect 14657 9129 14691 9163
rect 15393 9129 15427 9163
rect 15945 9129 15979 9163
rect 16589 9129 16623 9163
rect 2973 9061 3007 9095
rect 6377 9061 6411 9095
rect 6469 9061 6503 9095
rect 8493 9061 8527 9095
rect 1409 8993 1443 9027
rect 2421 8993 2455 9027
rect 8401 8993 8435 9027
rect 9956 8993 9990 9027
rect 12725 8993 12759 9027
rect 12981 8993 13015 9027
rect 16405 8993 16439 9027
rect 4629 8925 4663 8959
rect 6561 8925 6595 8959
rect 7021 8925 7055 8959
rect 8677 8925 8711 8959
rect 9689 8925 9723 8959
rect 1593 8857 1627 8891
rect 6009 8857 6043 8891
rect 8033 8857 8067 8891
rect 14105 8857 14139 8891
rect 11069 8789 11103 8823
rect 11621 8789 11655 8823
rect 12541 8789 12575 8823
rect 2053 8585 2087 8619
rect 2421 8585 2455 8619
rect 4445 8585 4479 8619
rect 4813 8585 4847 8619
rect 5733 8585 5767 8619
rect 7481 8585 7515 8619
rect 7757 8585 7791 8619
rect 10793 8585 10827 8619
rect 11897 8585 11931 8619
rect 13829 8585 13863 8619
rect 16405 8585 16439 8619
rect 1685 8517 1719 8551
rect 6101 8517 6135 8551
rect 6469 8517 6503 8551
rect 9321 8517 9355 8551
rect 10333 8517 10367 8551
rect 4169 8449 4203 8483
rect 6929 8449 6963 8483
rect 11253 8449 11287 8483
rect 11437 8449 11471 8483
rect 1501 8381 1535 8415
rect 7941 8381 7975 8415
rect 8208 8381 8242 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 12705 8381 12739 8415
rect 10609 8313 10643 8347
rect 11161 8313 11195 8347
rect 9965 8245 9999 8279
rect 1685 8041 1719 8075
rect 7941 8041 7975 8075
rect 8309 8041 8343 8075
rect 8769 8041 8803 8075
rect 9965 8041 9999 8075
rect 11805 8041 11839 8075
rect 12357 8041 12391 8075
rect 12725 8041 12759 8075
rect 12909 8041 12943 8075
rect 10425 7905 10459 7939
rect 10692 7905 10726 7939
rect 10425 7497 10459 7531
rect 10793 7497 10827 7531
rect 11069 5865 11103 5899
rect 9689 5729 9723 5763
rect 9956 5729 9990 5763
rect 10057 5321 10091 5355
rect 9781 4981 9815 5015
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 3326 25372 3332 25424
rect 3384 25412 3390 25424
rect 7929 25415 7987 25421
rect 7929 25412 7941 25415
rect 3384 25384 7941 25412
rect 3384 25372 3390 25384
rect 7929 25381 7941 25384
rect 7975 25381 7987 25415
rect 7929 25375 7987 25381
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1854 25344 1860 25356
rect 1443 25316 1860 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 2314 25304 2320 25356
rect 2372 25344 2378 25356
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2372 25316 2513 25344
rect 2372 25304 2378 25316
rect 2501 25313 2513 25316
rect 2547 25313 2559 25347
rect 3050 25344 3056 25356
rect 3011 25316 3056 25344
rect 2501 25307 2559 25313
rect 3050 25304 3056 25316
rect 3108 25304 3114 25356
rect 4706 25344 4712 25356
rect 4667 25316 4712 25344
rect 4706 25304 4712 25316
rect 4764 25304 4770 25356
rect 4798 25276 4804 25288
rect 4759 25248 4804 25276
rect 4798 25236 4804 25248
rect 4856 25236 4862 25288
rect 4982 25276 4988 25288
rect 4943 25248 4988 25276
rect 4982 25236 4988 25248
rect 5040 25236 5046 25288
rect 6914 25276 6920 25288
rect 6875 25248 6920 25276
rect 6914 25236 6920 25248
rect 6972 25236 6978 25288
rect 2409 25211 2467 25217
rect 2409 25177 2421 25211
rect 2455 25208 2467 25211
rect 2958 25208 2964 25220
rect 2455 25180 2964 25208
rect 2455 25177 2467 25180
rect 2409 25171 2467 25177
rect 2958 25168 2964 25180
rect 3016 25168 3022 25220
rect 4341 25211 4399 25217
rect 4341 25177 4353 25211
rect 4387 25208 4399 25211
rect 9122 25208 9128 25220
rect 4387 25180 9128 25208
rect 4387 25177 4399 25180
rect 4341 25171 4399 25177
rect 9122 25168 9128 25180
rect 9180 25168 9186 25220
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2866 25140 2872 25152
rect 2731 25112 2872 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 8386 25140 8392 25152
rect 8347 25112 8392 25140
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 12897 25143 12955 25149
rect 12897 25109 12909 25143
rect 12943 25140 12955 25143
rect 13078 25140 13084 25152
rect 12943 25112 13084 25140
rect 12943 25109 12955 25112
rect 12897 25103 12955 25109
rect 13078 25100 13084 25112
rect 13136 25100 13142 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1872 24908 2728 24936
rect 1872 24880 1900 24908
rect 1854 24868 1860 24880
rect 1815 24840 1860 24868
rect 1854 24828 1860 24840
rect 1912 24828 1918 24880
rect 2314 24868 2320 24880
rect 2275 24840 2320 24868
rect 2314 24828 2320 24840
rect 2372 24828 2378 24880
rect 2700 24868 2728 24908
rect 5350 24868 5356 24880
rect 2700 24840 5356 24868
rect 5350 24828 5356 24840
rect 5408 24828 5414 24880
rect 2958 24760 2964 24812
rect 3016 24800 3022 24812
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 3016 24772 3065 24800
rect 3016 24760 3022 24772
rect 3053 24769 3065 24772
rect 3099 24800 3111 24803
rect 4617 24803 4675 24809
rect 4617 24800 4629 24803
rect 3099 24772 4629 24800
rect 3099 24769 3111 24772
rect 3053 24763 3111 24769
rect 4617 24769 4629 24772
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1670 24732 1676 24744
rect 1443 24704 1676 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1670 24692 1676 24704
rect 1728 24692 1734 24744
rect 2774 24692 2780 24744
rect 2832 24732 2838 24744
rect 3234 24732 3240 24744
rect 2832 24704 3240 24732
rect 2832 24692 2838 24704
rect 3234 24692 3240 24704
rect 3292 24692 3298 24744
rect 3418 24692 3424 24744
rect 3476 24732 3482 24744
rect 3513 24735 3571 24741
rect 3513 24732 3525 24735
rect 3476 24704 3525 24732
rect 3476 24692 3482 24704
rect 3513 24701 3525 24704
rect 3559 24732 3571 24735
rect 4341 24735 4399 24741
rect 4341 24732 4353 24735
rect 3559 24704 4353 24732
rect 3559 24701 3571 24704
rect 3513 24695 3571 24701
rect 4341 24701 4353 24704
rect 4387 24732 4399 24735
rect 4632 24732 4660 24763
rect 4706 24760 4712 24812
rect 4764 24800 4770 24812
rect 5077 24803 5135 24809
rect 5077 24800 5089 24803
rect 4764 24772 5089 24800
rect 4764 24760 4770 24772
rect 5077 24769 5089 24772
rect 5123 24800 5135 24803
rect 6825 24803 6883 24809
rect 6825 24800 6837 24803
rect 5123 24772 6837 24800
rect 5123 24769 5135 24772
rect 5077 24763 5135 24769
rect 6825 24769 6837 24772
rect 6871 24769 6883 24803
rect 6825 24763 6883 24769
rect 7745 24803 7803 24809
rect 7745 24769 7757 24803
rect 7791 24800 7803 24803
rect 8202 24800 8208 24812
rect 7791 24772 8208 24800
rect 7791 24769 7803 24772
rect 7745 24763 7803 24769
rect 8202 24760 8208 24772
rect 8260 24800 8266 24812
rect 8297 24803 8355 24809
rect 8297 24800 8309 24803
rect 8260 24772 8309 24800
rect 8260 24760 8266 24772
rect 8297 24769 8309 24772
rect 8343 24769 8355 24803
rect 8297 24763 8355 24769
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 12250 24800 12256 24812
rect 8444 24772 8489 24800
rect 12211 24772 12256 24800
rect 8444 24760 8450 24772
rect 12250 24760 12256 24772
rect 12308 24800 12314 24812
rect 12897 24803 12955 24809
rect 12897 24800 12909 24803
rect 12308 24772 12909 24800
rect 12308 24760 12314 24772
rect 12897 24769 12909 24772
rect 12943 24769 12955 24803
rect 13078 24800 13084 24812
rect 13039 24772 13084 24800
rect 12897 24763 12955 24769
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 5353 24735 5411 24741
rect 5353 24732 5365 24735
rect 4387 24704 4568 24732
rect 4632 24704 5365 24732
rect 4387 24701 4399 24704
rect 4341 24695 4399 24701
rect 2869 24667 2927 24673
rect 2869 24633 2881 24667
rect 2915 24664 2927 24667
rect 3050 24664 3056 24676
rect 2915 24636 3056 24664
rect 2915 24633 2927 24636
rect 2869 24627 2927 24633
rect 3050 24624 3056 24636
rect 3108 24624 3114 24676
rect 3881 24667 3939 24673
rect 3881 24633 3893 24667
rect 3927 24664 3939 24667
rect 4540 24664 4568 24704
rect 5353 24701 5365 24704
rect 5399 24701 5411 24735
rect 5353 24695 5411 24701
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 6178 24732 6184 24744
rect 5583 24704 6184 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 6178 24692 6184 24704
rect 6236 24692 6242 24744
rect 9306 24692 9312 24744
rect 9364 24732 9370 24744
rect 9585 24735 9643 24741
rect 9585 24732 9597 24735
rect 9364 24704 9597 24732
rect 9364 24692 9370 24704
rect 9585 24701 9597 24704
rect 9631 24701 9643 24735
rect 9585 24695 9643 24701
rect 7377 24667 7435 24673
rect 7377 24664 7389 24667
rect 3927 24636 4476 24664
rect 4540 24636 7389 24664
rect 3927 24633 3939 24636
rect 3881 24627 3939 24633
rect 4448 24608 4476 24636
rect 7377 24633 7389 24636
rect 7423 24664 7435 24667
rect 9125 24667 9183 24673
rect 7423 24636 7972 24664
rect 7423 24633 7435 24636
rect 7377 24627 7435 24633
rect 7944 24608 7972 24636
rect 9125 24633 9137 24667
rect 9171 24664 9183 24667
rect 9490 24664 9496 24676
rect 9171 24636 9496 24664
rect 9171 24633 9183 24636
rect 9125 24627 9183 24633
rect 9490 24624 9496 24636
rect 9548 24664 9554 24676
rect 9830 24667 9888 24673
rect 9830 24664 9842 24667
rect 9548 24636 9842 24664
rect 9548 24624 9554 24636
rect 9830 24633 9842 24636
rect 9876 24633 9888 24667
rect 11790 24664 11796 24676
rect 11751 24636 11796 24664
rect 9830 24627 9888 24633
rect 11790 24624 11796 24636
rect 11848 24664 11854 24676
rect 12805 24667 12863 24673
rect 12805 24664 12817 24667
rect 11848 24636 12817 24664
rect 11848 24624 11854 24636
rect 12805 24633 12817 24636
rect 12851 24633 12863 24667
rect 12805 24627 12863 24633
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 1762 24596 1768 24608
rect 1627 24568 1768 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 1762 24556 1768 24568
rect 1820 24556 1826 24608
rect 2406 24596 2412 24608
rect 2367 24568 2412 24596
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 3970 24596 3976 24608
rect 3931 24568 3976 24596
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 4430 24596 4436 24608
rect 4391 24568 4436 24596
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 5534 24556 5540 24608
rect 5592 24596 5598 24608
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5592 24568 5733 24596
rect 5592 24556 5598 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 7834 24596 7840 24608
rect 7795 24568 7840 24596
rect 5721 24559 5779 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 7926 24556 7932 24608
rect 7984 24596 7990 24608
rect 8205 24599 8263 24605
rect 8205 24596 8217 24599
rect 7984 24568 8217 24596
rect 7984 24556 7990 24568
rect 8205 24565 8217 24568
rect 8251 24565 8263 24599
rect 8205 24559 8263 24565
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9401 24599 9459 24605
rect 9401 24596 9413 24599
rect 9364 24568 9413 24596
rect 9364 24556 9370 24568
rect 9401 24565 9413 24568
rect 9447 24565 9459 24599
rect 9401 24559 9459 24565
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 10965 24599 11023 24605
rect 10965 24596 10977 24599
rect 9732 24568 10977 24596
rect 9732 24556 9738 24568
rect 10965 24565 10977 24568
rect 11011 24565 11023 24599
rect 10965 24559 11023 24565
rect 12437 24599 12495 24605
rect 12437 24565 12449 24599
rect 12483 24596 12495 24599
rect 12526 24596 12532 24608
rect 12483 24568 12532 24596
rect 12483 24565 12495 24568
rect 12437 24559 12495 24565
rect 12526 24556 12532 24568
rect 12584 24556 12590 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 2406 24352 2412 24404
rect 2464 24392 2470 24404
rect 2590 24392 2596 24404
rect 2464 24364 2596 24392
rect 2464 24352 2470 24364
rect 2590 24352 2596 24364
rect 2648 24352 2654 24404
rect 3970 24392 3976 24404
rect 2700 24364 3976 24392
rect 2700 24333 2728 24364
rect 3970 24352 3976 24364
rect 4028 24352 4034 24404
rect 8018 24392 8024 24404
rect 7979 24364 8024 24392
rect 8018 24352 8024 24364
rect 8076 24352 8082 24404
rect 9766 24352 9772 24404
rect 9824 24392 9830 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9824 24364 10149 24392
rect 9824 24352 9830 24364
rect 10137 24361 10149 24364
rect 10183 24392 10195 24395
rect 10962 24392 10968 24404
rect 10183 24364 10968 24392
rect 10183 24361 10195 24364
rect 10137 24355 10195 24361
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 15654 24392 15660 24404
rect 15615 24364 15660 24392
rect 15654 24352 15660 24364
rect 15712 24352 15718 24404
rect 17310 24392 17316 24404
rect 17271 24364 17316 24392
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 21818 24392 21824 24404
rect 21779 24364 21824 24392
rect 21818 24352 21824 24364
rect 21876 24352 21882 24404
rect 23477 24395 23535 24401
rect 23477 24361 23489 24395
rect 23523 24392 23535 24395
rect 25314 24392 25320 24404
rect 23523 24364 25320 24392
rect 23523 24361 23535 24364
rect 23477 24355 23535 24361
rect 25314 24352 25320 24364
rect 25372 24352 25378 24404
rect 2133 24327 2191 24333
rect 2133 24293 2145 24327
rect 2179 24324 2191 24327
rect 2685 24327 2743 24333
rect 2685 24324 2697 24327
rect 2179 24296 2697 24324
rect 2179 24293 2191 24296
rect 2133 24287 2191 24293
rect 2685 24293 2697 24296
rect 2731 24293 2743 24327
rect 3234 24324 3240 24336
rect 3195 24296 3240 24324
rect 2685 24287 2743 24293
rect 3234 24284 3240 24296
rect 3292 24284 3298 24336
rect 3881 24327 3939 24333
rect 3881 24293 3893 24327
rect 3927 24324 3939 24327
rect 4798 24324 4804 24336
rect 3927 24296 4804 24324
rect 3927 24293 3939 24296
rect 3881 24287 3939 24293
rect 4798 24284 4804 24296
rect 4856 24284 4862 24336
rect 11606 24284 11612 24336
rect 11664 24333 11670 24336
rect 11664 24327 11728 24333
rect 11664 24293 11682 24327
rect 11716 24293 11728 24327
rect 11664 24287 11728 24293
rect 11664 24284 11670 24287
rect 5074 24265 5080 24268
rect 5068 24256 5080 24265
rect 5035 24228 5080 24256
rect 5068 24219 5080 24228
rect 5074 24216 5080 24219
rect 5132 24216 5138 24268
rect 7006 24216 7012 24268
rect 7064 24256 7070 24268
rect 7929 24259 7987 24265
rect 7929 24256 7941 24259
rect 7064 24228 7941 24256
rect 7064 24216 7070 24228
rect 7929 24225 7941 24228
rect 7975 24225 7987 24259
rect 7929 24219 7987 24225
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9640 24228 10057 24256
rect 9640 24216 9646 24228
rect 10045 24225 10057 24228
rect 10091 24225 10103 24259
rect 10045 24219 10103 24225
rect 15378 24216 15384 24268
rect 15436 24256 15442 24268
rect 15473 24259 15531 24265
rect 15473 24256 15485 24259
rect 15436 24228 15485 24256
rect 15436 24216 15442 24228
rect 15473 24225 15485 24228
rect 15519 24225 15531 24259
rect 17126 24256 17132 24268
rect 17087 24228 17132 24256
rect 15473 24219 15531 24225
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 21634 24256 21640 24268
rect 21595 24228 21640 24256
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 23290 24256 23296 24268
rect 23251 24228 23296 24256
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 2777 24191 2835 24197
rect 2777 24188 2789 24191
rect 2700 24160 2789 24188
rect 2700 24132 2728 24160
rect 2777 24157 2789 24160
rect 2823 24157 2835 24191
rect 2777 24151 2835 24157
rect 4614 24148 4620 24200
rect 4672 24188 4678 24200
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4672 24160 4813 24188
rect 4672 24148 4678 24160
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 8202 24188 8208 24200
rect 8163 24160 8208 24188
rect 4801 24151 4859 24157
rect 8202 24148 8208 24160
rect 8260 24188 8266 24200
rect 8386 24188 8392 24200
rect 8260 24160 8392 24188
rect 8260 24148 8266 24160
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 10318 24188 10324 24200
rect 10231 24160 10324 24188
rect 10318 24148 10324 24160
rect 10376 24188 10382 24200
rect 11422 24188 11428 24200
rect 10376 24160 10824 24188
rect 11383 24160 11428 24188
rect 10376 24148 10382 24160
rect 2682 24080 2688 24132
rect 2740 24080 2746 24132
rect 6917 24123 6975 24129
rect 6917 24089 6929 24123
rect 6963 24120 6975 24123
rect 7558 24120 7564 24132
rect 6963 24092 7564 24120
rect 6963 24089 6975 24092
rect 6917 24083 6975 24089
rect 7558 24080 7564 24092
rect 7616 24080 7622 24132
rect 1670 24052 1676 24064
rect 1631 24024 1676 24052
rect 1670 24012 1676 24024
rect 1728 24012 1734 24064
rect 2222 24052 2228 24064
rect 2183 24024 2228 24052
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 4433 24055 4491 24061
rect 4433 24021 4445 24055
rect 4479 24052 4491 24055
rect 4706 24052 4712 24064
rect 4479 24024 4712 24052
rect 4479 24021 4491 24024
rect 4433 24015 4491 24021
rect 4706 24012 4712 24024
rect 4764 24052 4770 24064
rect 4982 24052 4988 24064
rect 4764 24024 4988 24052
rect 4764 24012 4770 24024
rect 4982 24012 4988 24024
rect 5040 24052 5046 24064
rect 6181 24055 6239 24061
rect 6181 24052 6193 24055
rect 5040 24024 6193 24052
rect 5040 24012 5046 24024
rect 6181 24021 6193 24024
rect 6227 24021 6239 24055
rect 6181 24015 6239 24021
rect 7285 24055 7343 24061
rect 7285 24021 7297 24055
rect 7331 24052 7343 24055
rect 7742 24052 7748 24064
rect 7331 24024 7748 24052
rect 7331 24021 7343 24024
rect 7285 24015 7343 24021
rect 7742 24012 7748 24024
rect 7800 24012 7806 24064
rect 9677 24055 9735 24061
rect 9677 24021 9689 24055
rect 9723 24052 9735 24055
rect 10134 24052 10140 24064
rect 9723 24024 10140 24052
rect 9723 24021 9735 24024
rect 9677 24015 9735 24021
rect 10134 24012 10140 24024
rect 10192 24012 10198 24064
rect 10796 24061 10824 24160
rect 11422 24148 11428 24160
rect 11480 24148 11486 24200
rect 10781 24055 10839 24061
rect 10781 24021 10793 24055
rect 10827 24052 10839 24055
rect 12805 24055 12863 24061
rect 12805 24052 12817 24055
rect 10827 24024 12817 24052
rect 10827 24021 10839 24024
rect 10781 24015 10839 24021
rect 12805 24021 12817 24024
rect 12851 24021 12863 24055
rect 13906 24052 13912 24064
rect 13867 24024 13912 24052
rect 12805 24015 12863 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 4433 23851 4491 23857
rect 4433 23848 4445 23851
rect 4212 23820 4445 23848
rect 4212 23808 4218 23820
rect 4433 23817 4445 23820
rect 4479 23817 4491 23851
rect 4433 23811 4491 23817
rect 2317 23647 2375 23653
rect 2317 23613 2329 23647
rect 2363 23644 2375 23647
rect 2406 23644 2412 23656
rect 2363 23616 2412 23644
rect 2363 23613 2375 23616
rect 2317 23607 2375 23613
rect 2406 23604 2412 23616
rect 2464 23644 2470 23656
rect 4154 23644 4160 23656
rect 2464 23616 4160 23644
rect 2464 23604 2470 23616
rect 4154 23604 4160 23616
rect 4212 23604 4218 23656
rect 2562 23579 2620 23585
rect 2562 23576 2574 23579
rect 1780 23548 2574 23576
rect 1780 23520 1808 23548
rect 2562 23545 2574 23548
rect 2608 23576 2620 23579
rect 2682 23576 2688 23588
rect 2608 23548 2688 23576
rect 2608 23545 2620 23548
rect 2562 23539 2620 23545
rect 2682 23536 2688 23548
rect 2740 23536 2746 23588
rect 4448 23576 4476 23811
rect 4798 23808 4804 23860
rect 4856 23848 4862 23860
rect 4985 23851 5043 23857
rect 4985 23848 4997 23851
rect 4856 23820 4997 23848
rect 4856 23808 4862 23820
rect 4985 23817 4997 23820
rect 5031 23817 5043 23851
rect 6454 23848 6460 23860
rect 6415 23820 6460 23848
rect 4985 23811 5043 23817
rect 6454 23808 6460 23820
rect 6512 23808 6518 23860
rect 7006 23848 7012 23860
rect 6967 23820 7012 23848
rect 7006 23808 7012 23820
rect 7064 23848 7070 23860
rect 9309 23851 9367 23857
rect 9309 23848 9321 23851
rect 7064 23820 9321 23848
rect 7064 23808 7070 23820
rect 9309 23817 9321 23820
rect 9355 23848 9367 23851
rect 9582 23848 9588 23860
rect 9355 23820 9588 23848
rect 9355 23817 9367 23820
rect 9309 23811 9367 23817
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 9766 23848 9772 23860
rect 9727 23820 9772 23848
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 16482 23848 16488 23860
rect 16443 23820 16488 23848
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 18414 23848 18420 23860
rect 18375 23820 18420 23848
rect 18414 23808 18420 23820
rect 18472 23808 18478 23860
rect 19518 23848 19524 23860
rect 19479 23820 19524 23848
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 20622 23848 20628 23860
rect 20583 23820 20628 23848
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 21726 23848 21732 23860
rect 21687 23820 21732 23848
rect 21726 23808 21732 23820
rect 21784 23808 21790 23860
rect 23845 23851 23903 23857
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 24762 23848 24768 23860
rect 23891 23820 24768 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 5074 23672 5080 23724
rect 5132 23712 5138 23724
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5132 23684 5641 23712
rect 5132 23672 5138 23684
rect 5629 23681 5641 23684
rect 5675 23712 5687 23715
rect 6472 23712 6500 23808
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 8205 23783 8263 23789
rect 8205 23780 8217 23783
rect 8076 23752 8217 23780
rect 8076 23740 8082 23752
rect 8205 23749 8217 23752
rect 8251 23749 8263 23783
rect 8205 23743 8263 23749
rect 7742 23712 7748 23724
rect 5675 23684 6500 23712
rect 7703 23684 7748 23712
rect 5675 23681 5687 23684
rect 5629 23675 5687 23681
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 8662 23672 8668 23724
rect 8720 23712 8726 23724
rect 9306 23712 9312 23724
rect 8720 23684 9312 23712
rect 8720 23672 8726 23684
rect 9306 23672 9312 23684
rect 9364 23712 9370 23724
rect 9858 23712 9864 23724
rect 9364 23684 9864 23712
rect 9364 23672 9370 23684
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 15470 23672 15476 23724
rect 15528 23712 15534 23724
rect 16206 23712 16212 23724
rect 15528 23684 16212 23712
rect 15528 23672 15534 23684
rect 16206 23672 16212 23684
rect 16264 23672 16270 23724
rect 4893 23647 4951 23653
rect 4893 23613 4905 23647
rect 4939 23644 4951 23647
rect 5442 23644 5448 23656
rect 4939 23616 5448 23644
rect 4939 23613 4951 23616
rect 4893 23607 4951 23613
rect 5442 23604 5448 23616
rect 5500 23604 5506 23656
rect 7558 23644 7564 23656
rect 7519 23616 7564 23644
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 7653 23647 7711 23653
rect 7653 23613 7665 23647
rect 7699 23644 7711 23647
rect 7834 23644 7840 23656
rect 7699 23616 7840 23644
rect 7699 23613 7711 23616
rect 7653 23607 7711 23613
rect 7834 23604 7840 23616
rect 7892 23604 7898 23656
rect 8202 23604 8208 23656
rect 8260 23644 8266 23656
rect 8573 23647 8631 23653
rect 8573 23644 8585 23647
rect 8260 23616 8585 23644
rect 8260 23604 8266 23616
rect 8573 23613 8585 23616
rect 8619 23613 8631 23647
rect 8573 23607 8631 23613
rect 8849 23647 8907 23653
rect 8849 23613 8861 23647
rect 8895 23644 8907 23647
rect 9674 23644 9680 23656
rect 8895 23616 9680 23644
rect 8895 23613 8907 23616
rect 8849 23607 8907 23613
rect 9674 23604 9680 23616
rect 9732 23604 9738 23656
rect 13817 23647 13875 23653
rect 13817 23644 13829 23647
rect 13648 23616 13829 23644
rect 5258 23576 5264 23588
rect 4448 23548 5264 23576
rect 5258 23536 5264 23548
rect 5316 23576 5322 23588
rect 5353 23579 5411 23585
rect 5353 23576 5365 23579
rect 5316 23548 5365 23576
rect 5316 23536 5322 23548
rect 5353 23545 5365 23548
rect 5399 23545 5411 23579
rect 5353 23539 5411 23545
rect 9582 23536 9588 23588
rect 9640 23576 9646 23588
rect 10128 23579 10186 23585
rect 10128 23576 10140 23579
rect 9640 23548 10140 23576
rect 9640 23536 9646 23548
rect 10128 23545 10140 23548
rect 10174 23576 10186 23579
rect 10318 23576 10324 23588
rect 10174 23548 10324 23576
rect 10174 23545 10186 23548
rect 10128 23539 10186 23545
rect 10318 23536 10324 23548
rect 10376 23536 10382 23588
rect 11054 23536 11060 23588
rect 11112 23576 11118 23588
rect 11606 23576 11612 23588
rect 11112 23548 11612 23576
rect 11112 23536 11118 23548
rect 11606 23536 11612 23548
rect 11664 23576 11670 23588
rect 12161 23579 12219 23585
rect 12161 23576 12173 23579
rect 11664 23548 12173 23576
rect 11664 23536 11670 23548
rect 12161 23545 12173 23548
rect 12207 23576 12219 23579
rect 12342 23576 12348 23588
rect 12207 23548 12348 23576
rect 12207 23545 12219 23548
rect 12161 23539 12219 23545
rect 12342 23536 12348 23548
rect 12400 23536 12406 23588
rect 13648 23520 13676 23616
rect 13817 23613 13829 23616
rect 13863 23613 13875 23647
rect 16301 23647 16359 23653
rect 16301 23644 16313 23647
rect 13817 23607 13875 23613
rect 16132 23616 16313 23644
rect 13906 23536 13912 23588
rect 13964 23576 13970 23588
rect 14062 23579 14120 23585
rect 14062 23576 14074 23579
rect 13964 23548 14074 23576
rect 13964 23536 13970 23548
rect 14062 23545 14074 23548
rect 14108 23545 14120 23579
rect 14062 23539 14120 23545
rect 14826 23536 14832 23588
rect 14884 23576 14890 23588
rect 15378 23576 15384 23588
rect 14884 23548 15384 23576
rect 14884 23536 14890 23548
rect 15378 23536 15384 23548
rect 15436 23576 15442 23588
rect 15749 23579 15807 23585
rect 15749 23576 15761 23579
rect 15436 23548 15761 23576
rect 15436 23536 15442 23548
rect 15749 23545 15761 23548
rect 15795 23545 15807 23579
rect 15749 23539 15807 23545
rect 1762 23508 1768 23520
rect 1723 23480 1768 23508
rect 1762 23468 1768 23480
rect 1820 23468 1826 23520
rect 2225 23511 2283 23517
rect 2225 23477 2237 23511
rect 2271 23508 2283 23511
rect 2406 23508 2412 23520
rect 2271 23480 2412 23508
rect 2271 23477 2283 23480
rect 2225 23471 2283 23477
rect 2406 23468 2412 23480
rect 2464 23468 2470 23520
rect 3697 23511 3755 23517
rect 3697 23477 3709 23511
rect 3743 23508 3755 23511
rect 3878 23508 3884 23520
rect 3743 23480 3884 23508
rect 3743 23477 3755 23480
rect 3697 23471 3755 23477
rect 3878 23468 3884 23480
rect 3936 23468 3942 23520
rect 4614 23468 4620 23520
rect 4672 23508 4678 23520
rect 5997 23511 6055 23517
rect 5997 23508 6009 23511
rect 4672 23480 6009 23508
rect 4672 23468 4678 23480
rect 5997 23477 6009 23480
rect 6043 23508 6055 23511
rect 6822 23508 6828 23520
rect 6043 23480 6828 23508
rect 6043 23477 6055 23480
rect 5997 23471 6055 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 7193 23511 7251 23517
rect 7193 23508 7205 23511
rect 7156 23480 7205 23508
rect 7156 23468 7162 23480
rect 7193 23477 7205 23480
rect 7239 23477 7251 23511
rect 7193 23471 7251 23477
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11241 23511 11299 23517
rect 11241 23508 11253 23511
rect 11020 23480 11253 23508
rect 11020 23468 11026 23480
rect 11241 23477 11253 23480
rect 11287 23477 11299 23511
rect 11241 23471 11299 23477
rect 11422 23468 11428 23520
rect 11480 23508 11486 23520
rect 11793 23511 11851 23517
rect 11793 23508 11805 23511
rect 11480 23480 11805 23508
rect 11480 23468 11486 23480
rect 11793 23477 11805 23480
rect 11839 23477 11851 23511
rect 12802 23508 12808 23520
rect 12763 23480 12808 23508
rect 11793 23471 11851 23477
rect 12802 23468 12808 23480
rect 12860 23468 12866 23520
rect 13630 23508 13636 23520
rect 13591 23480 13636 23508
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 15194 23508 15200 23520
rect 15155 23480 15200 23508
rect 15194 23468 15200 23480
rect 15252 23468 15258 23520
rect 16022 23468 16028 23520
rect 16080 23508 16086 23520
rect 16132 23517 16160 23616
rect 16301 23613 16313 23616
rect 16347 23613 16359 23647
rect 18230 23644 18236 23656
rect 18191 23616 18236 23644
rect 16301 23607 16359 23613
rect 18230 23604 18236 23616
rect 18288 23644 18294 23656
rect 18785 23647 18843 23653
rect 18785 23644 18797 23647
rect 18288 23616 18797 23644
rect 18288 23604 18294 23616
rect 18785 23613 18797 23616
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 19337 23647 19395 23653
rect 19337 23613 19349 23647
rect 19383 23613 19395 23647
rect 19337 23607 19395 23613
rect 19352 23576 19380 23607
rect 19426 23604 19432 23656
rect 19484 23644 19490 23656
rect 20441 23647 20499 23653
rect 20441 23644 20453 23647
rect 19484 23616 20453 23644
rect 19484 23604 19490 23616
rect 20441 23613 20453 23616
rect 20487 23644 20499 23647
rect 20993 23647 21051 23653
rect 20993 23644 21005 23647
rect 20487 23616 21005 23644
rect 20487 23613 20499 23616
rect 20441 23607 20499 23613
rect 20993 23613 21005 23616
rect 21039 23613 21051 23647
rect 20993 23607 21051 23613
rect 21174 23604 21180 23656
rect 21232 23644 21238 23656
rect 21545 23647 21603 23653
rect 21545 23644 21557 23647
rect 21232 23616 21557 23644
rect 21232 23604 21238 23616
rect 21545 23613 21557 23616
rect 21591 23644 21603 23647
rect 22097 23647 22155 23653
rect 22097 23644 22109 23647
rect 21591 23616 22109 23644
rect 21591 23613 21603 23616
rect 21545 23607 21603 23613
rect 22097 23613 22109 23616
rect 22143 23613 22155 23647
rect 22097 23607 22155 23613
rect 23661 23647 23719 23653
rect 23661 23613 23673 23647
rect 23707 23644 23719 23647
rect 24762 23644 24768 23656
rect 23707 23616 24256 23644
rect 24723 23616 24768 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 19889 23579 19947 23585
rect 19889 23576 19901 23579
rect 19352 23548 19901 23576
rect 19352 23520 19380 23548
rect 19889 23545 19901 23548
rect 19935 23545 19947 23579
rect 19889 23539 19947 23545
rect 21634 23536 21640 23588
rect 21692 23576 21698 23588
rect 22465 23579 22523 23585
rect 22465 23576 22477 23579
rect 21692 23548 22477 23576
rect 21692 23536 21698 23548
rect 22465 23545 22477 23548
rect 22511 23545 22523 23579
rect 22465 23539 22523 23545
rect 24228 23520 24256 23616
rect 24762 23604 24768 23616
rect 24820 23644 24826 23656
rect 25317 23647 25375 23653
rect 25317 23644 25329 23647
rect 24820 23616 25329 23644
rect 24820 23604 24826 23616
rect 25317 23613 25329 23616
rect 25363 23613 25375 23647
rect 25317 23607 25375 23613
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 16080 23480 16129 23508
rect 16080 23468 16086 23480
rect 16117 23477 16129 23480
rect 16163 23477 16175 23511
rect 16117 23471 16175 23477
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 17126 23508 17132 23520
rect 16632 23480 17132 23508
rect 16632 23468 16638 23480
rect 17126 23468 17132 23480
rect 17184 23468 17190 23520
rect 19334 23468 19340 23520
rect 19392 23468 19398 23520
rect 22278 23468 22284 23520
rect 22336 23508 22342 23520
rect 23290 23508 23296 23520
rect 22336 23480 23296 23508
rect 22336 23468 22342 23480
rect 23290 23468 23296 23480
rect 23348 23468 23354 23520
rect 24210 23508 24216 23520
rect 24171 23480 24216 23508
rect 24210 23468 24216 23480
rect 24268 23468 24274 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2501 23307 2559 23313
rect 2501 23273 2513 23307
rect 2547 23304 2559 23307
rect 2590 23304 2596 23316
rect 2547 23276 2596 23304
rect 2547 23273 2559 23276
rect 2501 23267 2559 23273
rect 2590 23264 2596 23276
rect 2648 23264 2654 23316
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 3421 23307 3479 23313
rect 3421 23304 3433 23307
rect 2832 23276 3433 23304
rect 2832 23264 2838 23276
rect 3421 23273 3433 23276
rect 3467 23273 3479 23307
rect 3421 23267 3479 23273
rect 4525 23307 4583 23313
rect 4525 23273 4537 23307
rect 4571 23304 4583 23307
rect 4982 23304 4988 23316
rect 4571 23276 4988 23304
rect 4571 23273 4583 23276
rect 4525 23267 4583 23273
rect 4982 23264 4988 23276
rect 5040 23264 5046 23316
rect 7009 23307 7067 23313
rect 7009 23273 7021 23307
rect 7055 23304 7067 23307
rect 7834 23304 7840 23316
rect 7055 23276 7840 23304
rect 7055 23273 7067 23276
rect 7009 23267 7067 23273
rect 7834 23264 7840 23276
rect 7892 23264 7898 23316
rect 8481 23307 8539 23313
rect 8481 23273 8493 23307
rect 8527 23273 8539 23307
rect 8481 23267 8539 23273
rect 9493 23307 9551 23313
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 9582 23304 9588 23316
rect 9539 23276 9588 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 2409 23239 2467 23245
rect 2409 23205 2421 23239
rect 2455 23236 2467 23239
rect 2961 23239 3019 23245
rect 2961 23236 2973 23239
rect 2455 23208 2973 23236
rect 2455 23205 2467 23208
rect 2409 23199 2467 23205
rect 2961 23205 2973 23208
rect 3007 23236 3019 23239
rect 3234 23236 3240 23248
rect 3007 23208 3240 23236
rect 3007 23205 3019 23208
rect 2961 23199 3019 23205
rect 3234 23196 3240 23208
rect 3292 23196 3298 23248
rect 7742 23196 7748 23248
rect 7800 23236 7806 23248
rect 8496 23236 8524 23267
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10045 23307 10103 23313
rect 10045 23304 10057 23307
rect 9732 23276 10057 23304
rect 9732 23264 9738 23276
rect 10045 23273 10057 23276
rect 10091 23273 10103 23307
rect 10045 23267 10103 23273
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 10192 23276 10237 23304
rect 10192 23264 10198 23276
rect 12434 23264 12440 23316
rect 12492 23304 12498 23316
rect 13357 23307 13415 23313
rect 13357 23304 13369 23307
rect 12492 23276 13369 23304
rect 12492 23264 12498 23276
rect 13357 23273 13369 23276
rect 13403 23273 13415 23307
rect 13357 23267 13415 23273
rect 15473 23307 15531 23313
rect 15473 23273 15485 23307
rect 15519 23304 15531 23307
rect 16482 23304 16488 23316
rect 15519 23276 16488 23304
rect 15519 23273 15531 23276
rect 15473 23267 15531 23273
rect 16482 23264 16488 23276
rect 16540 23264 16546 23316
rect 16758 23304 16764 23316
rect 16719 23276 16764 23304
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 19061 23307 19119 23313
rect 19061 23273 19073 23307
rect 19107 23304 19119 23307
rect 19242 23304 19248 23316
rect 19107 23276 19248 23304
rect 19107 23273 19119 23276
rect 19061 23267 19119 23273
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 21085 23307 21143 23313
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 21634 23304 21640 23316
rect 21131 23276 21640 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 22370 23304 22376 23316
rect 22331 23276 22376 23304
rect 22370 23264 22376 23276
rect 22428 23264 22434 23316
rect 24026 23304 24032 23316
rect 23987 23276 24032 23304
rect 24026 23264 24032 23276
rect 24084 23264 24090 23316
rect 7800 23208 8524 23236
rect 7800 23196 7806 23208
rect 9858 23196 9864 23248
rect 9916 23236 9922 23248
rect 10689 23239 10747 23245
rect 10689 23236 10701 23239
rect 9916 23208 10701 23236
rect 9916 23196 9922 23208
rect 10689 23205 10701 23208
rect 10735 23236 10747 23239
rect 11422 23236 11428 23248
rect 10735 23208 11428 23236
rect 10735 23205 10747 23208
rect 10689 23199 10747 23205
rect 11422 23196 11428 23208
rect 11480 23236 11486 23248
rect 12250 23245 12256 23248
rect 12244 23236 12256 23245
rect 11480 23208 12020 23236
rect 12211 23208 12256 23236
rect 11480 23196 11486 23208
rect 11992 23180 12020 23208
rect 12244 23199 12256 23208
rect 12250 23196 12256 23199
rect 12308 23196 12314 23248
rect 1949 23171 2007 23177
rect 1949 23137 1961 23171
rect 1995 23168 2007 23171
rect 2314 23168 2320 23180
rect 1995 23140 2320 23168
rect 1995 23137 2007 23140
rect 1949 23131 2007 23137
rect 2314 23128 2320 23140
rect 2372 23168 2378 23180
rect 3050 23168 3056 23180
rect 2372 23140 3056 23168
rect 2372 23128 2378 23140
rect 3050 23128 3056 23140
rect 3108 23168 3114 23180
rect 3418 23168 3424 23180
rect 3108 23140 3424 23168
rect 3108 23128 3114 23140
rect 3418 23128 3424 23140
rect 3476 23128 3482 23180
rect 4154 23128 4160 23180
rect 4212 23168 4218 23180
rect 4614 23168 4620 23180
rect 4212 23140 4620 23168
rect 4212 23128 4218 23140
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 4706 23128 4712 23180
rect 4764 23168 4770 23180
rect 4873 23171 4931 23177
rect 4873 23168 4885 23171
rect 4764 23140 4885 23168
rect 4764 23128 4770 23140
rect 4873 23137 4885 23140
rect 4919 23137 4931 23171
rect 4873 23131 4931 23137
rect 7190 23128 7196 23180
rect 7248 23168 7254 23180
rect 7357 23171 7415 23177
rect 7357 23168 7369 23171
rect 7248 23140 7369 23168
rect 7248 23128 7254 23140
rect 7357 23137 7369 23140
rect 7403 23137 7415 23171
rect 11974 23168 11980 23180
rect 11887 23140 11980 23168
rect 7357 23131 7415 23137
rect 11974 23128 11980 23140
rect 12032 23128 12038 23180
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 16577 23171 16635 23177
rect 16577 23137 16589 23171
rect 16623 23168 16635 23171
rect 17310 23168 17316 23180
rect 16623 23140 17316 23168
rect 16623 23137 16635 23140
rect 16577 23131 16635 23137
rect 17310 23128 17316 23140
rect 17368 23128 17374 23180
rect 17862 23168 17868 23180
rect 17823 23140 17868 23168
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 18874 23168 18880 23180
rect 18835 23140 18880 23168
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 20806 23128 20812 23180
rect 20864 23168 20870 23180
rect 20901 23171 20959 23177
rect 20901 23168 20913 23171
rect 20864 23140 20913 23168
rect 20864 23128 20870 23140
rect 20901 23137 20913 23140
rect 20947 23137 20959 23171
rect 22186 23168 22192 23180
rect 22147 23140 22192 23168
rect 20901 23131 20959 23137
rect 22186 23128 22192 23140
rect 22244 23128 22250 23180
rect 23842 23168 23848 23180
rect 23803 23140 23848 23168
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 1762 23060 1768 23112
rect 1820 23100 1826 23112
rect 2593 23103 2651 23109
rect 2593 23100 2605 23103
rect 1820 23072 2605 23100
rect 1820 23060 1826 23072
rect 2593 23069 2605 23072
rect 2639 23100 2651 23103
rect 2639 23072 3188 23100
rect 2639 23069 2651 23072
rect 2593 23063 2651 23069
rect 2961 23035 3019 23041
rect 2961 23001 2973 23035
rect 3007 23032 3019 23035
rect 3050 23032 3056 23044
rect 3007 23004 3056 23032
rect 3007 23001 3019 23004
rect 2961 22995 3019 23001
rect 3050 22992 3056 23004
rect 3108 22992 3114 23044
rect 3160 23041 3188 23072
rect 6822 23060 6828 23112
rect 6880 23100 6886 23112
rect 7006 23100 7012 23112
rect 6880 23072 7012 23100
rect 6880 23060 6886 23072
rect 7006 23060 7012 23072
rect 7064 23100 7070 23112
rect 7101 23103 7159 23109
rect 7101 23100 7113 23103
rect 7064 23072 7113 23100
rect 7064 23060 7070 23072
rect 7101 23069 7113 23072
rect 7147 23069 7159 23103
rect 7101 23063 7159 23069
rect 9490 23060 9496 23112
rect 9548 23100 9554 23112
rect 10229 23103 10287 23109
rect 10229 23100 10241 23103
rect 9548 23072 10241 23100
rect 9548 23060 9554 23072
rect 10229 23069 10241 23072
rect 10275 23100 10287 23103
rect 10962 23100 10968 23112
rect 10275 23072 10968 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 10962 23060 10968 23072
rect 11020 23060 11026 23112
rect 3145 23035 3203 23041
rect 3145 23001 3157 23035
rect 3191 23032 3203 23035
rect 18049 23035 18107 23041
rect 3191 23004 3280 23032
rect 3191 23001 3203 23004
rect 3145 22995 3203 23001
rect 3252 22976 3280 23004
rect 18049 23001 18061 23035
rect 18095 23032 18107 23035
rect 19334 23032 19340 23044
rect 18095 23004 19340 23032
rect 18095 23001 18107 23004
rect 18049 22995 18107 23001
rect 19334 22992 19340 23004
rect 19392 22992 19398 23044
rect 2038 22964 2044 22976
rect 1999 22936 2044 22964
rect 2038 22924 2044 22936
rect 2096 22924 2102 22976
rect 3234 22924 3240 22976
rect 3292 22924 3298 22976
rect 5997 22967 6055 22973
rect 5997 22933 6009 22967
rect 6043 22964 6055 22967
rect 6270 22964 6276 22976
rect 6043 22936 6276 22964
rect 6043 22933 6055 22936
rect 5997 22927 6055 22933
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 6638 22964 6644 22976
rect 6599 22936 6644 22964
rect 6638 22924 6644 22936
rect 6696 22924 6702 22976
rect 9677 22967 9735 22973
rect 9677 22933 9689 22967
rect 9723 22964 9735 22967
rect 10042 22964 10048 22976
rect 9723 22936 10048 22964
rect 9723 22933 9735 22936
rect 9677 22927 9735 22933
rect 10042 22924 10048 22936
rect 10100 22924 10106 22976
rect 10962 22924 10968 22976
rect 11020 22964 11026 22976
rect 11057 22967 11115 22973
rect 11057 22964 11069 22967
rect 11020 22936 11069 22964
rect 11020 22924 11026 22936
rect 11057 22933 11069 22936
rect 11103 22933 11115 22967
rect 11057 22927 11115 22933
rect 11146 22924 11152 22976
rect 11204 22964 11210 22976
rect 11425 22967 11483 22973
rect 11425 22964 11437 22967
rect 11204 22936 11437 22964
rect 11204 22924 11210 22936
rect 11425 22933 11437 22936
rect 11471 22933 11483 22967
rect 11425 22927 11483 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2406 22760 2412 22772
rect 2148 22732 2412 22760
rect 2148 22565 2176 22732
rect 2406 22720 2412 22732
rect 2464 22720 2470 22772
rect 3234 22720 3240 22772
rect 3292 22760 3298 22772
rect 3513 22763 3571 22769
rect 3513 22760 3525 22763
rect 3292 22732 3525 22760
rect 3292 22720 3298 22732
rect 3513 22729 3525 22732
rect 3559 22729 3571 22763
rect 3513 22723 3571 22729
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 4249 22763 4307 22769
rect 4249 22760 4261 22763
rect 4212 22732 4261 22760
rect 4212 22720 4218 22732
rect 4249 22729 4261 22732
rect 4295 22729 4307 22763
rect 4614 22760 4620 22772
rect 4575 22732 4620 22760
rect 4249 22723 4307 22729
rect 4614 22720 4620 22732
rect 4672 22720 4678 22772
rect 6641 22763 6699 22769
rect 6641 22729 6653 22763
rect 6687 22760 6699 22763
rect 7190 22760 7196 22772
rect 6687 22732 7196 22760
rect 6687 22729 6699 22732
rect 6641 22723 6699 22729
rect 7190 22720 7196 22732
rect 7248 22760 7254 22772
rect 8110 22760 8116 22772
rect 7248 22732 8116 22760
rect 7248 22720 7254 22732
rect 8110 22720 8116 22732
rect 8168 22720 8174 22772
rect 9674 22760 9680 22772
rect 9635 22732 9680 22760
rect 9674 22720 9680 22732
rect 9732 22720 9738 22772
rect 11330 22720 11336 22772
rect 11388 22760 11394 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 11388 22732 11713 22760
rect 11388 22720 11394 22732
rect 11701 22729 11713 22732
rect 11747 22760 11759 22763
rect 12250 22760 12256 22772
rect 11747 22732 12256 22760
rect 11747 22729 11759 22732
rect 11701 22723 11759 22729
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 16485 22763 16543 22769
rect 16485 22760 16497 22763
rect 16448 22732 16497 22760
rect 16448 22720 16454 22732
rect 16485 22729 16497 22732
rect 16531 22729 16543 22763
rect 16485 22723 16543 22729
rect 7006 22652 7012 22704
rect 7064 22692 7070 22704
rect 7101 22695 7159 22701
rect 7101 22692 7113 22695
rect 7064 22664 7113 22692
rect 7064 22652 7070 22664
rect 7101 22661 7113 22664
rect 7147 22692 7159 22695
rect 7561 22695 7619 22701
rect 7561 22692 7573 22695
rect 7147 22664 7573 22692
rect 7147 22661 7159 22664
rect 7101 22655 7159 22661
rect 7561 22661 7573 22664
rect 7607 22661 7619 22695
rect 11974 22692 11980 22704
rect 11935 22664 11980 22692
rect 7561 22655 7619 22661
rect 5077 22627 5135 22633
rect 5077 22593 5089 22627
rect 5123 22624 5135 22627
rect 5626 22624 5632 22636
rect 5123 22596 5632 22624
rect 5123 22593 5135 22596
rect 5077 22587 5135 22593
rect 5626 22584 5632 22596
rect 5684 22584 5690 22636
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 6270 22624 6276 22636
rect 5859 22596 6276 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 6270 22584 6276 22596
rect 6328 22584 6334 22636
rect 7576 22624 7604 22655
rect 11974 22652 11980 22664
rect 12032 22692 12038 22704
rect 12342 22692 12348 22704
rect 12032 22664 12348 22692
rect 12032 22652 12038 22664
rect 12342 22652 12348 22664
rect 12400 22652 12406 22704
rect 22741 22695 22799 22701
rect 22741 22661 22753 22695
rect 22787 22692 22799 22695
rect 23842 22692 23848 22704
rect 22787 22664 23848 22692
rect 22787 22661 22799 22664
rect 22741 22655 22799 22661
rect 23842 22652 23848 22664
rect 23900 22652 23906 22704
rect 7745 22627 7803 22633
rect 7745 22624 7757 22627
rect 7576 22596 7757 22624
rect 7745 22593 7757 22596
rect 7791 22593 7803 22627
rect 11054 22624 11060 22636
rect 11015 22596 11060 22624
rect 7745 22587 7803 22593
rect 2133 22559 2191 22565
rect 2133 22556 2145 22559
rect 1688 22528 2145 22556
rect 1688 22432 1716 22528
rect 2133 22525 2145 22528
rect 2179 22525 2191 22559
rect 2133 22519 2191 22525
rect 4614 22516 4620 22568
rect 4672 22556 4678 22568
rect 5537 22559 5595 22565
rect 5537 22556 5549 22559
rect 4672 22528 5549 22556
rect 4672 22516 4678 22528
rect 5537 22525 5549 22528
rect 5583 22556 5595 22559
rect 6546 22556 6552 22568
rect 5583 22528 6552 22556
rect 5583 22525 5595 22528
rect 5537 22519 5595 22525
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 7760 22556 7788 22587
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 10962 22556 10968 22568
rect 7760 22528 8156 22556
rect 10923 22528 10968 22556
rect 8128 22500 8156 22528
rect 10962 22516 10968 22528
rect 11020 22516 11026 22568
rect 13265 22559 13323 22565
rect 13265 22525 13277 22559
rect 13311 22556 13323 22559
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 13311 22528 13553 22556
rect 13311 22525 13323 22528
rect 13265 22519 13323 22525
rect 13541 22525 13553 22528
rect 13587 22556 13599 22559
rect 13630 22556 13636 22568
rect 13587 22528 13636 22556
rect 13587 22525 13599 22528
rect 13541 22519 13599 22525
rect 13630 22516 13636 22528
rect 13688 22516 13694 22568
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 16301 22559 16359 22565
rect 16301 22556 16313 22559
rect 15620 22528 16313 22556
rect 15620 22516 15626 22528
rect 16301 22525 16313 22528
rect 16347 22556 16359 22559
rect 16761 22559 16819 22565
rect 16761 22556 16773 22559
rect 16347 22528 16773 22556
rect 16347 22525 16359 22528
rect 16301 22519 16359 22525
rect 16761 22525 16773 22528
rect 16807 22525 16819 22559
rect 22554 22556 22560 22568
rect 22515 22528 22560 22556
rect 16761 22519 16819 22525
rect 22554 22516 22560 22528
rect 22612 22556 22618 22568
rect 23017 22559 23075 22565
rect 23017 22556 23029 22559
rect 22612 22528 23029 22556
rect 22612 22516 22618 22528
rect 23017 22525 23029 22528
rect 23063 22525 23075 22559
rect 23017 22519 23075 22525
rect 2314 22448 2320 22500
rect 2372 22497 2378 22500
rect 2372 22491 2436 22497
rect 2372 22457 2390 22491
rect 2424 22457 2436 22491
rect 2372 22451 2436 22457
rect 2372 22448 2378 22451
rect 7834 22448 7840 22500
rect 7892 22488 7898 22500
rect 7990 22491 8048 22497
rect 7990 22488 8002 22491
rect 7892 22460 8002 22488
rect 7892 22448 7898 22460
rect 7990 22457 8002 22460
rect 8036 22457 8048 22491
rect 7990 22451 8048 22457
rect 8110 22448 8116 22500
rect 8168 22448 8174 22500
rect 9766 22448 9772 22500
rect 9824 22488 9830 22500
rect 10413 22491 10471 22497
rect 10413 22488 10425 22491
rect 9824 22460 10425 22488
rect 9824 22448 9830 22460
rect 10413 22457 10425 22460
rect 10459 22488 10471 22491
rect 10873 22491 10931 22497
rect 10873 22488 10885 22491
rect 10459 22460 10885 22488
rect 10459 22457 10471 22460
rect 10413 22451 10471 22457
rect 10873 22457 10885 22460
rect 10919 22457 10931 22491
rect 12434 22488 12440 22500
rect 12395 22460 12440 22488
rect 10873 22451 10931 22457
rect 12434 22448 12440 22460
rect 12492 22448 12498 22500
rect 13078 22488 13084 22500
rect 12991 22460 13084 22488
rect 13078 22448 13084 22460
rect 13136 22488 13142 22500
rect 13808 22491 13866 22497
rect 13808 22488 13820 22491
rect 13136 22460 13820 22488
rect 13136 22448 13142 22460
rect 13808 22457 13820 22460
rect 13854 22488 13866 22491
rect 14366 22488 14372 22500
rect 13854 22460 14372 22488
rect 13854 22457 13866 22460
rect 13808 22451 13866 22457
rect 14366 22448 14372 22460
rect 14424 22448 14430 22500
rect 16206 22448 16212 22500
rect 16264 22488 16270 22500
rect 17862 22488 17868 22500
rect 16264 22460 17868 22488
rect 16264 22448 16270 22460
rect 17862 22448 17868 22460
rect 17920 22488 17926 22500
rect 18233 22491 18291 22497
rect 18233 22488 18245 22491
rect 17920 22460 18245 22488
rect 17920 22448 17926 22460
rect 18233 22457 18245 22460
rect 18279 22457 18291 22491
rect 18233 22451 18291 22457
rect 1670 22420 1676 22432
rect 1631 22392 1676 22420
rect 1670 22380 1676 22392
rect 1728 22380 1734 22432
rect 2041 22423 2099 22429
rect 2041 22389 2053 22423
rect 2087 22420 2099 22423
rect 2590 22420 2596 22432
rect 2087 22392 2596 22420
rect 2087 22389 2099 22392
rect 2041 22383 2099 22389
rect 2590 22380 2596 22392
rect 2648 22380 2654 22432
rect 5169 22423 5227 22429
rect 5169 22389 5181 22423
rect 5215 22420 5227 22423
rect 5442 22420 5448 22432
rect 5215 22392 5448 22420
rect 5215 22389 5227 22392
rect 5169 22383 5227 22389
rect 5442 22380 5448 22392
rect 5500 22380 5506 22432
rect 6270 22420 6276 22432
rect 6231 22392 6276 22420
rect 6270 22380 6276 22392
rect 6328 22380 6334 22432
rect 8938 22380 8944 22432
rect 8996 22420 9002 22432
rect 9125 22423 9183 22429
rect 9125 22420 9137 22423
rect 8996 22392 9137 22420
rect 8996 22380 9002 22392
rect 9125 22389 9137 22392
rect 9171 22389 9183 22423
rect 9125 22383 9183 22389
rect 10505 22423 10563 22429
rect 10505 22389 10517 22423
rect 10551 22420 10563 22423
rect 10686 22420 10692 22432
rect 10551 22392 10692 22420
rect 10551 22389 10563 22392
rect 10505 22383 10563 22389
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 13265 22423 13323 22429
rect 13265 22420 13277 22423
rect 12400 22392 13277 22420
rect 12400 22380 12406 22392
rect 13265 22389 13277 22392
rect 13311 22420 13323 22423
rect 13357 22423 13415 22429
rect 13357 22420 13369 22423
rect 13311 22392 13369 22420
rect 13311 22389 13323 22392
rect 13265 22383 13323 22389
rect 13357 22389 13369 22392
rect 13403 22389 13415 22423
rect 13357 22383 13415 22389
rect 13906 22380 13912 22432
rect 13964 22420 13970 22432
rect 14921 22423 14979 22429
rect 14921 22420 14933 22423
rect 13964 22392 14933 22420
rect 13964 22380 13970 22392
rect 14921 22389 14933 22392
rect 14967 22389 14979 22423
rect 14921 22383 14979 22389
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 15565 22423 15623 22429
rect 15565 22420 15577 22423
rect 15344 22392 15577 22420
rect 15344 22380 15350 22392
rect 15565 22389 15577 22392
rect 15611 22420 15623 22423
rect 15930 22420 15936 22432
rect 15611 22392 15936 22420
rect 15611 22389 15623 22392
rect 15565 22383 15623 22389
rect 15930 22380 15936 22392
rect 15988 22380 15994 22432
rect 17221 22423 17279 22429
rect 17221 22389 17233 22423
rect 17267 22420 17279 22423
rect 17310 22420 17316 22432
rect 17267 22392 17316 22420
rect 17267 22389 17279 22392
rect 17221 22383 17279 22389
rect 17310 22380 17316 22392
rect 17368 22380 17374 22432
rect 18874 22420 18880 22432
rect 18835 22392 18880 22420
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 20806 22380 20812 22432
rect 20864 22420 20870 22432
rect 20901 22423 20959 22429
rect 20901 22420 20913 22423
rect 20864 22392 20913 22420
rect 20864 22380 20870 22392
rect 20901 22389 20913 22392
rect 20947 22389 20959 22423
rect 22186 22420 22192 22432
rect 22147 22392 22192 22420
rect 20901 22383 20959 22389
rect 22186 22380 22192 22392
rect 22244 22380 22250 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1673 22219 1731 22225
rect 1673 22185 1685 22219
rect 1719 22216 1731 22219
rect 1762 22216 1768 22228
rect 1719 22188 1768 22216
rect 1719 22185 1731 22188
rect 1673 22179 1731 22185
rect 1762 22176 1768 22188
rect 1820 22176 1826 22228
rect 2038 22176 2044 22228
rect 2096 22216 2102 22228
rect 2133 22219 2191 22225
rect 2133 22216 2145 22219
rect 2096 22188 2145 22216
rect 2096 22176 2102 22188
rect 2133 22185 2145 22188
rect 2179 22185 2191 22219
rect 2133 22179 2191 22185
rect 2148 22148 2176 22179
rect 2222 22176 2228 22228
rect 2280 22216 2286 22228
rect 2280 22188 2325 22216
rect 2280 22176 2286 22188
rect 2498 22176 2504 22228
rect 2556 22216 2562 22228
rect 4065 22219 4123 22225
rect 4065 22216 4077 22219
rect 2556 22188 4077 22216
rect 2556 22176 2562 22188
rect 4065 22185 4077 22188
rect 4111 22185 4123 22219
rect 4706 22216 4712 22228
rect 4667 22188 4712 22216
rect 4065 22179 4123 22185
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 5074 22216 5080 22228
rect 5035 22188 5080 22216
rect 5074 22176 5080 22188
rect 5132 22176 5138 22228
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 7009 22219 7067 22225
rect 7009 22216 7021 22219
rect 6696 22188 7021 22216
rect 6696 22176 6702 22188
rect 7009 22185 7021 22188
rect 7055 22185 7067 22219
rect 7742 22216 7748 22228
rect 7703 22188 7748 22216
rect 7009 22179 7067 22185
rect 7742 22176 7748 22188
rect 7800 22216 7806 22228
rect 8021 22219 8079 22225
rect 8021 22216 8033 22219
rect 7800 22188 8033 22216
rect 7800 22176 7806 22188
rect 8021 22185 8033 22188
rect 8067 22185 8079 22219
rect 9766 22216 9772 22228
rect 9727 22188 9772 22216
rect 8021 22179 8079 22185
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 10781 22219 10839 22225
rect 10781 22185 10793 22219
rect 10827 22216 10839 22219
rect 10962 22216 10968 22228
rect 10827 22188 10968 22216
rect 10827 22185 10839 22188
rect 10781 22179 10839 22185
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 12342 22176 12348 22228
rect 12400 22216 12406 22228
rect 12802 22216 12808 22228
rect 12400 22188 12808 22216
rect 12400 22176 12406 22188
rect 12802 22176 12808 22188
rect 12860 22216 12866 22228
rect 12989 22219 13047 22225
rect 12989 22216 13001 22219
rect 12860 22188 13001 22216
rect 12860 22176 12866 22188
rect 12989 22185 13001 22188
rect 13035 22185 13047 22219
rect 12989 22179 13047 22185
rect 2682 22148 2688 22160
rect 2148 22120 2688 22148
rect 2682 22108 2688 22120
rect 2740 22108 2746 22160
rect 5445 22151 5503 22157
rect 5445 22117 5457 22151
rect 5491 22148 5503 22151
rect 6362 22148 6368 22160
rect 5491 22120 6368 22148
rect 5491 22117 5503 22120
rect 5445 22111 5503 22117
rect 6362 22108 6368 22120
rect 6420 22108 6426 22160
rect 7926 22108 7932 22160
rect 7984 22148 7990 22160
rect 8110 22148 8116 22160
rect 7984 22120 8116 22148
rect 7984 22108 7990 22120
rect 8110 22108 8116 22120
rect 8168 22108 8174 22160
rect 10134 22148 10140 22160
rect 9600 22120 10140 22148
rect 2869 22083 2927 22089
rect 2869 22049 2881 22083
rect 2915 22080 2927 22083
rect 3050 22080 3056 22092
rect 2915 22052 3056 22080
rect 2915 22049 2927 22052
rect 2869 22043 2927 22049
rect 3050 22040 3056 22052
rect 3108 22040 3114 22092
rect 8205 22083 8263 22089
rect 8205 22049 8217 22083
rect 8251 22080 8263 22083
rect 8573 22083 8631 22089
rect 8573 22080 8585 22083
rect 8251 22052 8585 22080
rect 8251 22049 8263 22052
rect 8205 22043 8263 22049
rect 8573 22049 8585 22052
rect 8619 22049 8631 22083
rect 9490 22080 9496 22092
rect 9451 22052 9496 22080
rect 8573 22043 8631 22049
rect 9490 22040 9496 22052
rect 9548 22040 9554 22092
rect 2406 22012 2412 22024
rect 2367 21984 2412 22012
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 5534 22012 5540 22024
rect 5495 21984 5540 22012
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 5721 22015 5779 22021
rect 5721 21981 5733 22015
rect 5767 22012 5779 22015
rect 5994 22012 6000 22024
rect 5767 21984 6000 22012
rect 5767 21981 5779 21984
rect 5721 21975 5779 21981
rect 5994 21972 6000 21984
rect 6052 21972 6058 22024
rect 7098 22012 7104 22024
rect 7059 21984 7104 22012
rect 7098 21972 7104 21984
rect 7156 21972 7162 22024
rect 7193 22015 7251 22021
rect 7193 21981 7205 22015
rect 7239 22012 7251 22015
rect 8938 22012 8944 22024
rect 7239 21984 8944 22012
rect 7239 21981 7251 21984
rect 7193 21975 7251 21981
rect 2222 21904 2228 21956
rect 2280 21944 2286 21956
rect 3697 21947 3755 21953
rect 3697 21944 3709 21947
rect 2280 21916 3709 21944
rect 2280 21904 2286 21916
rect 3697 21913 3709 21916
rect 3743 21913 3755 21947
rect 3697 21907 3755 21913
rect 6549 21947 6607 21953
rect 6549 21913 6561 21947
rect 6595 21944 6607 21947
rect 7208 21944 7236 21975
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9600 22012 9628 22120
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 10597 22151 10655 22157
rect 10597 22117 10609 22151
rect 10643 22148 10655 22151
rect 11054 22148 11060 22160
rect 10643 22120 11060 22148
rect 10643 22117 10655 22120
rect 10597 22111 10655 22117
rect 11054 22108 11060 22120
rect 11112 22108 11118 22160
rect 11149 22151 11207 22157
rect 11149 22117 11161 22151
rect 11195 22148 11207 22151
rect 11606 22148 11612 22160
rect 11195 22120 11612 22148
rect 11195 22117 11207 22120
rect 11149 22111 11207 22117
rect 11606 22108 11612 22120
rect 11664 22108 11670 22160
rect 10870 22040 10876 22092
rect 10928 22080 10934 22092
rect 11241 22083 11299 22089
rect 11241 22080 11253 22083
rect 10928 22052 11253 22080
rect 10928 22040 10934 22052
rect 11241 22049 11253 22052
rect 11287 22080 11299 22083
rect 11698 22080 11704 22092
rect 11287 22052 11704 22080
rect 11287 22049 11299 22052
rect 11241 22043 11299 22049
rect 11698 22040 11704 22052
rect 11756 22040 11762 22092
rect 12161 22083 12219 22089
rect 12161 22049 12173 22083
rect 12207 22080 12219 22083
rect 12526 22080 12532 22092
rect 12207 22052 12532 22080
rect 12207 22049 12219 22052
rect 12161 22043 12219 22049
rect 12526 22040 12532 22052
rect 12584 22080 12590 22092
rect 13081 22083 13139 22089
rect 13081 22080 13093 22083
rect 12584 22052 13093 22080
rect 12584 22040 12590 22052
rect 13081 22049 13093 22052
rect 13127 22049 13139 22083
rect 13081 22043 13139 22049
rect 11330 22012 11336 22024
rect 9171 21984 9628 22012
rect 11291 21984 11336 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 11330 21972 11336 21984
rect 11388 21972 11394 22024
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 22012 12495 22015
rect 13265 22015 13323 22021
rect 13265 22012 13277 22015
rect 12483 21984 13277 22012
rect 12483 21981 12495 21984
rect 12437 21975 12495 21981
rect 13265 21981 13277 21984
rect 13311 22012 13323 22015
rect 13906 22012 13912 22024
rect 13311 21984 13912 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 6595 21916 7236 21944
rect 6595 21913 6607 21916
rect 6549 21907 6607 21913
rect 8018 21904 8024 21956
rect 8076 21944 8082 21956
rect 8662 21944 8668 21956
rect 8076 21916 8668 21944
rect 8076 21904 8082 21916
rect 8662 21904 8668 21916
rect 8720 21904 8726 21956
rect 1765 21879 1823 21885
rect 1765 21845 1777 21879
rect 1811 21876 1823 21879
rect 2038 21876 2044 21888
rect 1811 21848 2044 21876
rect 1811 21845 1823 21848
rect 1765 21839 1823 21845
rect 2038 21836 2044 21848
rect 2096 21836 2102 21888
rect 3326 21876 3332 21888
rect 3239 21848 3332 21876
rect 3326 21836 3332 21848
rect 3384 21876 3390 21888
rect 3602 21876 3608 21888
rect 3384 21848 3608 21876
rect 3384 21836 3390 21848
rect 3602 21836 3608 21848
rect 3660 21836 3666 21888
rect 6178 21876 6184 21888
rect 6139 21848 6184 21876
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 6638 21876 6644 21888
rect 6599 21848 6644 21876
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 8389 21879 8447 21885
rect 8389 21845 8401 21879
rect 8435 21876 8447 21879
rect 8478 21876 8484 21888
rect 8435 21848 8484 21876
rect 8435 21845 8447 21848
rect 8389 21839 8447 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 8573 21879 8631 21885
rect 8573 21845 8585 21879
rect 8619 21876 8631 21879
rect 8757 21879 8815 21885
rect 8757 21876 8769 21879
rect 8619 21848 8769 21876
rect 8619 21845 8631 21848
rect 8573 21839 8631 21845
rect 8757 21845 8769 21848
rect 8803 21876 8815 21879
rect 9582 21876 9588 21888
rect 8803 21848 9588 21876
rect 8803 21845 8815 21848
rect 8757 21839 8815 21845
rect 9582 21836 9588 21848
rect 9640 21836 9646 21888
rect 12621 21879 12679 21885
rect 12621 21845 12633 21879
rect 12667 21876 12679 21879
rect 12710 21876 12716 21888
rect 12667 21848 12716 21876
rect 12667 21845 12679 21848
rect 12621 21839 12679 21845
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 13630 21876 13636 21888
rect 13591 21848 13636 21876
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 2041 21675 2099 21681
rect 2041 21641 2053 21675
rect 2087 21672 2099 21675
rect 2130 21672 2136 21684
rect 2087 21644 2136 21672
rect 2087 21641 2099 21644
rect 2041 21635 2099 21641
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21468 1455 21471
rect 2056 21468 2084 21635
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 4522 21672 4528 21684
rect 4483 21644 4528 21672
rect 4522 21632 4528 21644
rect 4580 21632 4586 21684
rect 6089 21675 6147 21681
rect 6089 21641 6101 21675
rect 6135 21672 6147 21675
rect 6362 21672 6368 21684
rect 6135 21644 6368 21672
rect 6135 21641 6147 21644
rect 6089 21635 6147 21641
rect 6362 21632 6368 21644
rect 6420 21632 6426 21684
rect 6546 21672 6552 21684
rect 6507 21644 6552 21672
rect 6546 21632 6552 21644
rect 6604 21632 6610 21684
rect 6730 21632 6736 21684
rect 6788 21672 6794 21684
rect 6825 21675 6883 21681
rect 6825 21672 6837 21675
rect 6788 21644 6837 21672
rect 6788 21632 6794 21644
rect 6825 21641 6837 21644
rect 6871 21641 6883 21675
rect 6825 21635 6883 21641
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21672 8631 21675
rect 8662 21672 8668 21684
rect 8619 21644 8668 21672
rect 8619 21641 8631 21644
rect 8573 21635 8631 21641
rect 8662 21632 8668 21644
rect 8720 21632 8726 21684
rect 10870 21672 10876 21684
rect 10831 21644 10876 21672
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 11606 21672 11612 21684
rect 11567 21644 11612 21672
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 12253 21675 12311 21681
rect 12253 21641 12265 21675
rect 12299 21672 12311 21675
rect 12342 21672 12348 21684
rect 12299 21644 12348 21672
rect 12299 21641 12311 21644
rect 12253 21635 12311 21641
rect 12342 21632 12348 21644
rect 12400 21632 12406 21684
rect 14366 21672 14372 21684
rect 14327 21644 14372 21672
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 3145 21539 3203 21545
rect 3145 21505 3157 21539
rect 3191 21536 3203 21539
rect 3694 21536 3700 21548
rect 3191 21508 3700 21536
rect 3191 21505 3203 21508
rect 3145 21499 3203 21505
rect 3694 21496 3700 21508
rect 3752 21496 3758 21548
rect 3881 21539 3939 21545
rect 3881 21505 3893 21539
rect 3927 21536 3939 21539
rect 3970 21536 3976 21548
rect 3927 21508 3976 21536
rect 3927 21505 3939 21508
rect 3881 21499 3939 21505
rect 1443 21440 2084 21468
rect 2777 21471 2835 21477
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 2777 21437 2789 21471
rect 2823 21468 2835 21471
rect 3896 21468 3924 21499
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 5074 21496 5080 21548
rect 5132 21536 5138 21548
rect 5537 21539 5595 21545
rect 5537 21536 5549 21539
rect 5132 21508 5549 21536
rect 5132 21496 5138 21508
rect 5537 21505 5549 21508
rect 5583 21536 5595 21539
rect 6178 21536 6184 21548
rect 5583 21508 6184 21536
rect 5583 21505 5595 21508
rect 5537 21499 5595 21505
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 6564 21536 6592 21632
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 6564 21508 7297 21536
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 7742 21536 7748 21548
rect 7515 21508 7748 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 8680 21545 8708 21632
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 2823 21440 3924 21468
rect 2823 21437 2835 21440
rect 2777 21431 2835 21437
rect 4062 21428 4068 21480
rect 4120 21468 4126 21480
rect 4890 21468 4896 21480
rect 4120 21440 4896 21468
rect 4120 21428 4126 21440
rect 4890 21428 4896 21440
rect 4948 21468 4954 21480
rect 5445 21471 5503 21477
rect 5445 21468 5457 21471
rect 4948 21440 5457 21468
rect 4948 21428 4954 21440
rect 5445 21437 5457 21440
rect 5491 21437 5503 21471
rect 5445 21431 5503 21437
rect 6914 21428 6920 21480
rect 6972 21468 6978 21480
rect 8938 21477 8944 21480
rect 7193 21471 7251 21477
rect 7193 21468 7205 21471
rect 6972 21440 7205 21468
rect 6972 21428 6978 21440
rect 7193 21437 7205 21440
rect 7239 21468 7251 21471
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7239 21440 7849 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 8932 21468 8944 21477
rect 8899 21440 8944 21468
rect 7837 21431 7895 21437
rect 8932 21431 8944 21440
rect 8938 21428 8944 21431
rect 8996 21428 9002 21480
rect 11146 21468 11152 21480
rect 11107 21440 11152 21468
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 12989 21471 13047 21477
rect 12989 21468 13001 21471
rect 12820 21440 13001 21468
rect 2406 21400 2412 21412
rect 2319 21372 2412 21400
rect 2406 21360 2412 21372
rect 2464 21400 2470 21412
rect 3878 21400 3884 21412
rect 2464 21372 3884 21400
rect 2464 21360 2470 21372
rect 3878 21360 3884 21372
rect 3936 21400 3942 21412
rect 4338 21400 4344 21412
rect 3936 21372 4344 21400
rect 3936 21360 3942 21372
rect 4338 21360 4344 21372
rect 4396 21360 4402 21412
rect 4522 21360 4528 21412
rect 4580 21400 4586 21412
rect 5350 21400 5356 21412
rect 4580 21372 5356 21400
rect 4580 21360 4586 21372
rect 5350 21360 5356 21372
rect 5408 21360 5414 21412
rect 3234 21332 3240 21344
rect 3195 21304 3240 21332
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 3602 21332 3608 21344
rect 3563 21304 3608 21332
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 4982 21332 4988 21344
rect 4943 21304 4988 21332
rect 4982 21292 4988 21304
rect 5040 21292 5046 21344
rect 9950 21292 9956 21344
rect 10008 21332 10014 21344
rect 10045 21335 10103 21341
rect 10045 21332 10057 21335
rect 10008 21304 10057 21332
rect 10008 21292 10014 21304
rect 10045 21301 10057 21304
rect 10091 21301 10103 21335
rect 10045 21295 10103 21301
rect 11238 21292 11244 21344
rect 11296 21332 11302 21344
rect 11333 21335 11391 21341
rect 11333 21332 11345 21335
rect 11296 21304 11345 21332
rect 11296 21292 11302 21304
rect 11333 21301 11345 21304
rect 11379 21301 11391 21335
rect 11333 21295 11391 21301
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12820 21341 12848 21440
rect 12989 21437 13001 21440
rect 13035 21437 13047 21471
rect 12989 21431 13047 21437
rect 13256 21471 13314 21477
rect 13256 21437 13268 21471
rect 13302 21468 13314 21471
rect 13630 21468 13636 21480
rect 13302 21440 13636 21468
rect 13302 21437 13314 21440
rect 13256 21431 13314 21437
rect 13630 21428 13636 21440
rect 13688 21428 13694 21480
rect 26234 21360 26240 21412
rect 26292 21400 26298 21412
rect 27614 21400 27620 21412
rect 26292 21372 27620 21400
rect 26292 21360 26298 21372
rect 27614 21360 27620 21372
rect 27672 21360 27678 21412
rect 12805 21335 12863 21341
rect 12805 21332 12817 21335
rect 12492 21304 12817 21332
rect 12492 21292 12498 21304
rect 12805 21301 12817 21304
rect 12851 21301 12863 21335
rect 12805 21295 12863 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 1762 21088 1768 21140
rect 1820 21128 1826 21140
rect 1949 21131 2007 21137
rect 1949 21128 1961 21131
rect 1820 21100 1961 21128
rect 1820 21088 1826 21100
rect 1949 21097 1961 21100
rect 1995 21097 2007 21131
rect 1949 21091 2007 21097
rect 2774 21088 2780 21140
rect 2832 21128 2838 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 2832 21100 3801 21128
rect 2832 21088 2838 21100
rect 3789 21097 3801 21100
rect 3835 21097 3847 21131
rect 3789 21091 3847 21097
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 6365 21131 6423 21137
rect 6365 21128 6377 21131
rect 5592 21100 6377 21128
rect 5592 21088 5598 21100
rect 6365 21097 6377 21100
rect 6411 21097 6423 21131
rect 6365 21091 6423 21097
rect 7098 21088 7104 21140
rect 7156 21128 7162 21140
rect 9033 21131 9091 21137
rect 9033 21128 9045 21131
rect 7156 21100 9045 21128
rect 7156 21088 7162 21100
rect 9033 21097 9045 21100
rect 9079 21097 9091 21131
rect 10134 21128 10140 21140
rect 10095 21100 10140 21128
rect 9033 21091 9091 21097
rect 10134 21088 10140 21100
rect 10192 21088 10198 21140
rect 11241 21131 11299 21137
rect 11241 21097 11253 21131
rect 11287 21128 11299 21131
rect 11330 21128 11336 21140
rect 11287 21100 11336 21128
rect 11287 21097 11299 21100
rect 11241 21091 11299 21097
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 13630 21088 13636 21140
rect 13688 21128 13694 21140
rect 13817 21131 13875 21137
rect 13817 21128 13829 21131
rect 13688 21100 13829 21128
rect 13688 21088 13694 21100
rect 13817 21097 13829 21100
rect 13863 21097 13875 21131
rect 13817 21091 13875 21097
rect 5994 21060 6000 21072
rect 5955 21032 6000 21060
rect 5994 21020 6000 21032
rect 6052 21020 6058 21072
rect 6270 21020 6276 21072
rect 6328 21060 6334 21072
rect 6794 21063 6852 21069
rect 6794 21060 6806 21063
rect 6328 21032 6806 21060
rect 6328 21020 6334 21032
rect 6794 21029 6806 21032
rect 6840 21029 6852 21063
rect 6794 21023 6852 21029
rect 8757 21063 8815 21069
rect 8757 21029 8769 21063
rect 8803 21060 8815 21063
rect 8938 21060 8944 21072
rect 8803 21032 8944 21060
rect 8803 21029 8815 21032
rect 8757 21023 8815 21029
rect 8938 21020 8944 21032
rect 8996 21020 9002 21072
rect 1394 20992 1400 21004
rect 1355 20964 1400 20992
rect 1394 20952 1400 20964
rect 1452 20952 1458 21004
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 3142 20992 3148 21004
rect 2547 20964 3148 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 3142 20952 3148 20964
rect 3200 20952 3206 21004
rect 4062 20992 4068 21004
rect 4023 20964 4068 20992
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 4338 21001 4344 21004
rect 4332 20992 4344 21001
rect 4299 20964 4344 20992
rect 4332 20955 4344 20964
rect 4338 20952 4344 20955
rect 4396 20952 4402 21004
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 10410 20992 10416 21004
rect 10091 20964 10416 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 12704 20995 12762 21001
rect 12704 20992 12716 20995
rect 12268 20964 12716 20992
rect 6546 20924 6552 20936
rect 6507 20896 6552 20924
rect 6546 20884 6552 20896
rect 6604 20884 6610 20936
rect 9490 20924 9496 20936
rect 9403 20896 9496 20924
rect 9490 20884 9496 20896
rect 9548 20924 9554 20936
rect 9950 20924 9956 20936
rect 9548 20896 9956 20924
rect 9548 20884 9554 20896
rect 9950 20884 9956 20896
rect 10008 20924 10014 20936
rect 10229 20927 10287 20933
rect 10229 20924 10241 20927
rect 10008 20896 10241 20924
rect 10008 20884 10014 20896
rect 10229 20893 10241 20896
rect 10275 20893 10287 20927
rect 11422 20924 11428 20936
rect 11383 20896 11428 20924
rect 10229 20887 10287 20893
rect 11422 20884 11428 20896
rect 11480 20884 11486 20936
rect 2682 20856 2688 20868
rect 2643 20828 2688 20856
rect 2682 20816 2688 20828
rect 2740 20816 2746 20868
rect 2774 20816 2780 20868
rect 2832 20856 2838 20868
rect 12268 20865 12296 20964
rect 12704 20961 12716 20964
rect 12750 20992 12762 20995
rect 13446 20992 13452 21004
rect 12750 20964 13452 20992
rect 12750 20961 12762 20964
rect 12704 20955 12762 20961
rect 13446 20952 13452 20964
rect 13504 20952 13510 21004
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 12492 20896 12537 20924
rect 12492 20884 12498 20896
rect 3421 20859 3479 20865
rect 3421 20856 3433 20859
rect 2832 20828 3433 20856
rect 2832 20816 2838 20828
rect 3421 20825 3433 20828
rect 3467 20825 3479 20859
rect 3421 20819 3479 20825
rect 11977 20859 12035 20865
rect 11977 20825 11989 20859
rect 12023 20856 12035 20859
rect 12253 20859 12311 20865
rect 12253 20856 12265 20859
rect 12023 20828 12265 20856
rect 12023 20825 12035 20828
rect 11977 20819 12035 20825
rect 12253 20825 12265 20828
rect 12299 20825 12311 20859
rect 12253 20819 12311 20825
rect 2222 20748 2228 20800
rect 2280 20788 2286 20800
rect 2317 20791 2375 20797
rect 2317 20788 2329 20791
rect 2280 20760 2329 20788
rect 2280 20748 2286 20760
rect 2317 20757 2329 20760
rect 2363 20757 2375 20791
rect 2317 20751 2375 20757
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 5445 20791 5503 20797
rect 5445 20788 5457 20791
rect 5132 20760 5457 20788
rect 5132 20748 5138 20760
rect 5445 20757 5457 20760
rect 5491 20757 5503 20791
rect 5445 20751 5503 20757
rect 5994 20748 6000 20800
rect 6052 20788 6058 20800
rect 7929 20791 7987 20797
rect 7929 20788 7941 20791
rect 6052 20760 7941 20788
rect 6052 20748 6058 20760
rect 7929 20757 7941 20760
rect 7975 20757 7987 20791
rect 9674 20788 9680 20800
rect 9635 20760 9680 20788
rect 7929 20751 7987 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 10873 20791 10931 20797
rect 10873 20757 10885 20791
rect 10919 20788 10931 20791
rect 11330 20788 11336 20800
rect 10919 20760 11336 20788
rect 10919 20757 10931 20760
rect 10873 20751 10931 20757
rect 11330 20748 11336 20760
rect 11388 20788 11394 20800
rect 13630 20788 13636 20800
rect 11388 20760 13636 20788
rect 11388 20748 11394 20760
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 14366 20788 14372 20800
rect 14327 20760 14372 20788
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1394 20544 1400 20596
rect 1452 20584 1458 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1452 20556 1593 20584
rect 1452 20544 1458 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 3329 20587 3387 20593
rect 3329 20553 3341 20587
rect 3375 20584 3387 20587
rect 3418 20584 3424 20596
rect 3375 20556 3424 20584
rect 3375 20553 3387 20556
rect 3329 20547 3387 20553
rect 3418 20544 3424 20556
rect 3476 20544 3482 20596
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 4062 20584 4068 20596
rect 4019 20556 4068 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 4062 20544 4068 20556
rect 4120 20544 4126 20596
rect 4338 20544 4344 20596
rect 4396 20584 4402 20596
rect 5813 20587 5871 20593
rect 5813 20584 5825 20587
rect 4396 20556 5825 20584
rect 4396 20544 4402 20556
rect 5813 20553 5825 20556
rect 5859 20553 5871 20587
rect 6270 20584 6276 20596
rect 6231 20556 6276 20584
rect 5813 20547 5871 20553
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 6546 20544 6552 20596
rect 6604 20584 6610 20596
rect 6641 20587 6699 20593
rect 6641 20584 6653 20587
rect 6604 20556 6653 20584
rect 6604 20544 6610 20556
rect 6641 20553 6653 20556
rect 6687 20584 6699 20587
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 6687 20556 7941 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 7929 20553 7941 20556
rect 7975 20584 7987 20587
rect 8018 20584 8024 20596
rect 7975 20556 8024 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 8018 20544 8024 20556
rect 8076 20544 8082 20596
rect 10045 20587 10103 20593
rect 10045 20553 10057 20587
rect 10091 20584 10103 20587
rect 10134 20584 10140 20596
rect 10091 20556 10140 20584
rect 10091 20553 10103 20556
rect 10045 20547 10103 20553
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 13814 20584 13820 20596
rect 13775 20556 13820 20584
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 1762 20408 1768 20460
rect 1820 20448 1826 20460
rect 8036 20457 8064 20544
rect 10410 20516 10416 20528
rect 10371 20488 10416 20516
rect 10410 20476 10416 20488
rect 10468 20476 10474 20528
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 11256 20488 12449 20516
rect 11256 20460 11284 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12437 20479 12495 20485
rect 1949 20451 2007 20457
rect 1949 20448 1961 20451
rect 1820 20420 1961 20448
rect 1820 20408 1826 20420
rect 1949 20417 1961 20420
rect 1995 20417 2007 20451
rect 1949 20411 2007 20417
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 5077 20451 5135 20457
rect 4387 20420 4936 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 4908 20392 4936 20420
rect 5077 20417 5089 20451
rect 5123 20448 5135 20451
rect 8021 20451 8079 20457
rect 5123 20420 5580 20448
rect 5123 20417 5135 20420
rect 5077 20411 5135 20417
rect 2222 20389 2228 20392
rect 2216 20380 2228 20389
rect 2183 20352 2228 20380
rect 2216 20343 2228 20352
rect 2222 20340 2228 20343
rect 2280 20340 2286 20392
rect 4522 20340 4528 20392
rect 4580 20380 4586 20392
rect 4801 20383 4859 20389
rect 4801 20380 4813 20383
rect 4580 20352 4813 20380
rect 4580 20340 4586 20352
rect 4801 20349 4813 20352
rect 4847 20349 4859 20383
rect 4801 20343 4859 20349
rect 4890 20340 4896 20392
rect 4948 20380 4954 20392
rect 4948 20352 4993 20380
rect 4948 20340 4954 20352
rect 3970 20272 3976 20324
rect 4028 20312 4034 20324
rect 5092 20312 5120 20411
rect 5552 20321 5580 20420
rect 8021 20417 8033 20451
rect 8067 20417 8079 20451
rect 11238 20448 11244 20460
rect 11151 20420 11244 20448
rect 8021 20411 8079 20417
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 11330 20408 11336 20460
rect 11388 20448 11394 20460
rect 12253 20451 12311 20457
rect 11388 20420 11433 20448
rect 11388 20408 11394 20420
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12894 20448 12900 20460
rect 12299 20420 12900 20448
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13081 20451 13139 20457
rect 13081 20417 13093 20451
rect 13127 20448 13139 20451
rect 13446 20448 13452 20460
rect 13127 20420 13452 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 14366 20408 14372 20460
rect 14424 20448 14430 20460
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 14424 20420 14565 20448
rect 14424 20408 14430 20420
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 7009 20383 7067 20389
rect 7009 20349 7021 20383
rect 7055 20380 7067 20383
rect 7926 20380 7932 20392
rect 7055 20352 7932 20380
rect 7055 20349 7067 20352
rect 7009 20343 7067 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8294 20389 8300 20392
rect 8288 20380 8300 20389
rect 8220 20352 8300 20380
rect 4028 20284 5120 20312
rect 5537 20315 5595 20321
rect 4028 20272 4034 20284
rect 5537 20281 5549 20315
rect 5583 20312 5595 20315
rect 7561 20315 7619 20321
rect 5583 20284 7328 20312
rect 5583 20281 5595 20284
rect 5537 20275 5595 20281
rect 1670 20204 1676 20256
rect 1728 20244 1734 20256
rect 2314 20244 2320 20256
rect 1728 20216 2320 20244
rect 1728 20204 1734 20216
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 4430 20244 4436 20256
rect 4391 20216 4436 20244
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 7193 20247 7251 20253
rect 7193 20244 7205 20247
rect 7064 20216 7205 20244
rect 7064 20204 7070 20216
rect 7193 20213 7205 20216
rect 7239 20213 7251 20247
rect 7300 20244 7328 20284
rect 7561 20281 7573 20315
rect 7607 20312 7619 20315
rect 8220 20312 8248 20352
rect 8288 20343 8300 20352
rect 8294 20340 8300 20343
rect 8352 20340 8358 20392
rect 11149 20383 11207 20389
rect 11149 20349 11161 20383
rect 11195 20380 11207 20383
rect 11422 20380 11428 20392
rect 11195 20352 11428 20380
rect 11195 20349 11207 20352
rect 11149 20343 11207 20349
rect 11422 20340 11428 20352
rect 11480 20340 11486 20392
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 13872 20352 14473 20380
rect 13872 20340 13878 20352
rect 14461 20349 14473 20352
rect 14507 20349 14519 20383
rect 14461 20343 14519 20349
rect 9582 20312 9588 20324
rect 7607 20284 8248 20312
rect 8303 20284 9588 20312
rect 7607 20281 7619 20284
rect 7561 20275 7619 20281
rect 8303 20244 8331 20284
rect 9582 20272 9588 20284
rect 9640 20272 9646 20324
rect 11882 20312 11888 20324
rect 11795 20284 11888 20312
rect 11882 20272 11888 20284
rect 11940 20312 11946 20324
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 11940 20284 12817 20312
rect 11940 20272 11946 20284
rect 12805 20281 12817 20284
rect 12851 20281 12863 20315
rect 12805 20275 12863 20281
rect 13906 20272 13912 20324
rect 13964 20312 13970 20324
rect 14369 20315 14427 20321
rect 14369 20312 14381 20315
rect 13964 20284 14381 20312
rect 13964 20272 13970 20284
rect 14369 20281 14381 20284
rect 14415 20281 14427 20315
rect 14369 20275 14427 20281
rect 9398 20244 9404 20256
rect 7300 20216 8331 20244
rect 9359 20216 9404 20244
rect 7193 20207 7251 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 10781 20247 10839 20253
rect 10781 20213 10793 20247
rect 10827 20244 10839 20247
rect 10962 20244 10968 20256
rect 10827 20216 10968 20244
rect 10827 20213 10839 20216
rect 10781 20207 10839 20213
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 13541 20247 13599 20253
rect 13541 20213 13553 20247
rect 13587 20244 13599 20247
rect 13722 20244 13728 20256
rect 13587 20216 13728 20244
rect 13587 20213 13599 20216
rect 13541 20207 13599 20213
rect 13722 20204 13728 20216
rect 13780 20204 13786 20256
rect 13998 20244 14004 20256
rect 13959 20216 14004 20244
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1762 20040 1768 20052
rect 1504 20012 1768 20040
rect 1504 19913 1532 20012
rect 1762 20000 1768 20012
rect 1820 20000 1826 20052
rect 2222 20000 2228 20052
rect 2280 20040 2286 20052
rect 2590 20040 2596 20052
rect 2280 20012 2596 20040
rect 2280 20000 2286 20012
rect 2590 20000 2596 20012
rect 2648 20040 2654 20052
rect 2869 20043 2927 20049
rect 2869 20040 2881 20043
rect 2648 20012 2881 20040
rect 2648 20000 2654 20012
rect 2869 20009 2881 20012
rect 2915 20009 2927 20043
rect 2869 20003 2927 20009
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 3421 20043 3479 20049
rect 3421 20040 3433 20043
rect 3292 20012 3433 20040
rect 3292 20000 3298 20012
rect 3421 20009 3433 20012
rect 3467 20009 3479 20043
rect 4522 20040 4528 20052
rect 4483 20012 4528 20040
rect 3421 20003 3479 20009
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 6549 20043 6607 20049
rect 6549 20040 6561 20043
rect 5040 20012 6561 20040
rect 5040 20000 5046 20012
rect 6549 20009 6561 20012
rect 6595 20009 6607 20043
rect 6549 20003 6607 20009
rect 8113 20043 8171 20049
rect 8113 20009 8125 20043
rect 8159 20040 8171 20043
rect 8294 20040 8300 20052
rect 8159 20012 8300 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 9309 20043 9367 20049
rect 9309 20009 9321 20043
rect 9355 20040 9367 20043
rect 9398 20040 9404 20052
rect 9355 20012 9404 20040
rect 9355 20009 9367 20012
rect 9309 20003 9367 20009
rect 9398 20000 9404 20012
rect 9456 20000 9462 20052
rect 10042 20040 10048 20052
rect 10003 20012 10048 20040
rect 10042 20000 10048 20012
rect 10100 20040 10106 20052
rect 10778 20040 10784 20052
rect 10100 20012 10784 20040
rect 10100 20000 10106 20012
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 10873 20043 10931 20049
rect 10873 20009 10885 20043
rect 10919 20040 10931 20043
rect 11422 20040 11428 20052
rect 10919 20012 11428 20040
rect 10919 20009 10931 20012
rect 10873 20003 10931 20009
rect 11422 20000 11428 20012
rect 11480 20000 11486 20052
rect 13446 20040 13452 20052
rect 13407 20012 13452 20040
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 13906 20000 13912 20052
rect 13964 20040 13970 20052
rect 14001 20043 14059 20049
rect 14001 20040 14013 20043
rect 13964 20012 14013 20040
rect 13964 20000 13970 20012
rect 14001 20009 14013 20012
rect 14047 20009 14059 20043
rect 14001 20003 14059 20009
rect 5258 19972 5264 19984
rect 5219 19944 5264 19972
rect 5258 19932 5264 19944
rect 5316 19932 5322 19984
rect 5994 19932 6000 19984
rect 6052 19972 6058 19984
rect 6978 19975 7036 19981
rect 6978 19972 6990 19975
rect 6052 19944 6990 19972
rect 6052 19932 6058 19944
rect 6978 19941 6990 19944
rect 7024 19941 7036 19975
rect 6978 19935 7036 19941
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 10137 19975 10195 19981
rect 10137 19972 10149 19975
rect 8904 19944 10149 19972
rect 8904 19932 8910 19944
rect 10137 19941 10149 19944
rect 10183 19941 10195 19975
rect 11238 19972 11244 19984
rect 11199 19944 11244 19972
rect 10137 19935 10195 19941
rect 11238 19932 11244 19944
rect 11296 19932 11302 19984
rect 12342 19981 12348 19984
rect 11977 19975 12035 19981
rect 11977 19941 11989 19975
rect 12023 19972 12035 19975
rect 12314 19975 12348 19981
rect 12314 19972 12326 19975
rect 12023 19944 12326 19972
rect 12023 19941 12035 19944
rect 11977 19935 12035 19941
rect 12314 19941 12326 19944
rect 12314 19935 12348 19941
rect 12342 19932 12348 19935
rect 12400 19932 12406 19984
rect 1489 19907 1547 19913
rect 1489 19873 1501 19907
rect 1535 19873 1547 19907
rect 1489 19867 1547 19873
rect 1756 19907 1814 19913
rect 1756 19873 1768 19907
rect 1802 19904 1814 19907
rect 2314 19904 2320 19916
rect 1802 19876 2320 19904
rect 1802 19873 1814 19876
rect 1756 19867 1814 19873
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4580 19876 5181 19904
rect 4580 19864 4586 19876
rect 5169 19873 5181 19876
rect 5215 19873 5227 19907
rect 5169 19867 5227 19873
rect 6546 19864 6552 19916
rect 6604 19904 6610 19916
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 6604 19876 6745 19904
rect 6604 19864 6610 19876
rect 6733 19873 6745 19876
rect 6779 19873 6791 19907
rect 6733 19867 6791 19873
rect 5074 19796 5080 19848
rect 5132 19836 5138 19848
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 5132 19808 5365 19836
rect 5132 19796 5138 19808
rect 5353 19805 5365 19808
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 10192 19808 10241 19836
rect 10192 19796 10198 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 15378 19836 15384 19848
rect 15335 19808 15384 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 8018 19728 8024 19780
rect 8076 19768 8082 19780
rect 8665 19771 8723 19777
rect 8665 19768 8677 19771
rect 8076 19740 8677 19768
rect 8076 19728 8082 19740
rect 8665 19737 8677 19740
rect 8711 19737 8723 19771
rect 8665 19731 8723 19737
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3200 19672 3801 19700
rect 3200 19660 3206 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 3789 19663 3847 19669
rect 4801 19703 4859 19709
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 5166 19700 5172 19712
rect 4847 19672 5172 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 5813 19703 5871 19709
rect 5813 19700 5825 19703
rect 5500 19672 5825 19700
rect 5500 19660 5506 19672
rect 5813 19669 5825 19672
rect 5859 19669 5871 19703
rect 6178 19700 6184 19712
rect 6139 19672 6184 19700
rect 5813 19663 5871 19669
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 9674 19700 9680 19712
rect 9635 19672 9680 19700
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 12084 19700 12112 19799
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 12434 19700 12440 19712
rect 12084 19672 12440 19700
rect 12434 19660 12440 19672
rect 12492 19700 12498 19712
rect 13722 19700 13728 19712
rect 12492 19672 13728 19700
rect 12492 19660 12498 19672
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 14458 19700 14464 19712
rect 14419 19672 14464 19700
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2590 19496 2596 19508
rect 2551 19468 2596 19496
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 3142 19496 3148 19508
rect 3103 19468 3148 19496
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 12066 19456 12072 19508
rect 12124 19496 12130 19508
rect 12437 19499 12495 19505
rect 12437 19496 12449 19499
rect 12124 19468 12449 19496
rect 12124 19456 12130 19468
rect 12437 19465 12449 19468
rect 12483 19465 12495 19499
rect 12437 19459 12495 19465
rect 1946 19388 1952 19440
rect 2004 19428 2010 19440
rect 2406 19428 2412 19440
rect 2004 19400 2412 19428
rect 2004 19388 2010 19400
rect 2406 19388 2412 19400
rect 2464 19388 2470 19440
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 2608 19360 2636 19456
rect 3053 19431 3111 19437
rect 3053 19397 3065 19431
rect 3099 19428 3111 19431
rect 3326 19428 3332 19440
rect 3099 19400 3332 19428
rect 3099 19397 3111 19400
rect 3053 19391 3111 19397
rect 3326 19388 3332 19400
rect 3384 19428 3390 19440
rect 3384 19400 3740 19428
rect 3384 19388 3390 19400
rect 2271 19332 2636 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 3234 19320 3240 19372
rect 3292 19360 3298 19372
rect 3712 19369 3740 19400
rect 6178 19388 6184 19440
rect 6236 19428 6242 19440
rect 6825 19431 6883 19437
rect 6825 19428 6837 19431
rect 6236 19400 6837 19428
rect 6236 19388 6242 19400
rect 6825 19397 6837 19400
rect 6871 19397 6883 19431
rect 6825 19391 6883 19397
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 12676 19400 13124 19428
rect 12676 19388 12682 19400
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 3292 19332 3617 19360
rect 3292 19320 3298 19332
rect 3605 19329 3617 19332
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 4430 19360 4436 19372
rect 3697 19323 3755 19329
rect 4080 19332 4436 19360
rect 2041 19295 2099 19301
rect 2041 19261 2053 19295
rect 2087 19292 2099 19295
rect 3142 19292 3148 19304
rect 2087 19264 3148 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 3142 19252 3148 19264
rect 3200 19252 3206 19304
rect 3510 19292 3516 19304
rect 3423 19264 3516 19292
rect 3510 19252 3516 19264
rect 3568 19292 3574 19304
rect 4080 19292 4108 19332
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 5442 19360 5448 19372
rect 5403 19332 5448 19360
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 7374 19360 7380 19372
rect 7335 19332 7380 19360
rect 7374 19320 7380 19332
rect 7432 19360 7438 19372
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7432 19332 7849 19360
rect 7432 19320 7438 19332
rect 7837 19329 7849 19332
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 13096 19369 13124 19400
rect 13081 19363 13139 19369
rect 10836 19332 11008 19360
rect 10836 19320 10842 19332
rect 3568 19264 4108 19292
rect 3568 19252 3574 19264
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 5169 19295 5227 19301
rect 5169 19292 5181 19295
rect 5040 19264 5181 19292
rect 5040 19252 5046 19264
rect 5169 19261 5181 19264
rect 5215 19261 5227 19295
rect 5169 19255 5227 19261
rect 5261 19295 5319 19301
rect 5261 19261 5273 19295
rect 5307 19292 5319 19295
rect 6178 19292 6184 19304
rect 5307 19264 6184 19292
rect 5307 19261 5319 19264
rect 5261 19255 5319 19261
rect 6178 19252 6184 19264
rect 6236 19252 6242 19304
rect 6273 19295 6331 19301
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 7190 19292 7196 19304
rect 6319 19264 7196 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 8904 19264 9045 19292
rect 8904 19252 8910 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9214 19292 9220 19304
rect 9175 19264 9220 19292
rect 9033 19255 9091 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 10980 19292 11008 19332
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 14458 19320 14464 19372
rect 14516 19360 14522 19372
rect 14737 19363 14795 19369
rect 14737 19360 14749 19363
rect 14516 19332 14749 19360
rect 14516 19320 14522 19332
rect 14737 19329 14749 19332
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 10980 19264 11161 19292
rect 11149 19261 11161 19264
rect 11195 19292 11207 19295
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11195 19264 11805 19292
rect 11195 19261 11207 19264
rect 11149 19255 11207 19261
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 11793 19255 11851 19261
rect 12897 19295 12955 19301
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 13354 19292 13360 19304
rect 12943 19264 13360 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 1762 19184 1768 19236
rect 1820 19224 1826 19236
rect 1949 19227 2007 19233
rect 1949 19224 1961 19227
rect 1820 19196 1961 19224
rect 1820 19184 1826 19196
rect 1949 19193 1961 19196
rect 1995 19224 2007 19227
rect 2682 19224 2688 19236
rect 1995 19196 2688 19224
rect 1995 19193 2007 19196
rect 1949 19187 2007 19193
rect 2682 19184 2688 19196
rect 2740 19184 2746 19236
rect 4341 19227 4399 19233
rect 4341 19193 4353 19227
rect 4387 19224 4399 19227
rect 5905 19227 5963 19233
rect 4387 19196 5028 19224
rect 4387 19193 4399 19196
rect 4341 19187 4399 19193
rect 5000 19168 5028 19196
rect 5905 19193 5917 19227
rect 5951 19224 5963 19227
rect 5994 19224 6000 19236
rect 5951 19196 6000 19224
rect 5951 19193 5963 19196
rect 5905 19187 5963 19193
rect 5994 19184 6000 19196
rect 6052 19184 6058 19236
rect 6641 19227 6699 19233
rect 6641 19193 6653 19227
rect 6687 19224 6699 19227
rect 6687 19196 7328 19224
rect 6687 19193 6699 19196
rect 6641 19187 6699 19193
rect 7300 19168 7328 19196
rect 9398 19184 9404 19236
rect 9456 19233 9462 19236
rect 9456 19227 9520 19233
rect 9456 19193 9474 19227
rect 9508 19193 9520 19227
rect 9456 19187 9520 19193
rect 9456 19184 9462 19187
rect 1581 19159 1639 19165
rect 1581 19125 1593 19159
rect 1627 19156 1639 19159
rect 2130 19156 2136 19168
rect 1627 19128 2136 19156
rect 1627 19125 1639 19128
rect 1581 19119 1639 19125
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 4522 19116 4528 19168
rect 4580 19156 4586 19168
rect 4617 19159 4675 19165
rect 4617 19156 4629 19159
rect 4580 19128 4629 19156
rect 4580 19116 4586 19128
rect 4617 19125 4629 19128
rect 4663 19125 4675 19159
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4617 19119 4675 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 4982 19116 4988 19168
rect 5040 19116 5046 19168
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 8757 19159 8815 19165
rect 7340 19128 7385 19156
rect 7340 19116 7346 19128
rect 8757 19125 8769 19159
rect 8803 19156 8815 19159
rect 10134 19156 10140 19168
rect 8803 19128 10140 19156
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 10134 19116 10140 19128
rect 10192 19156 10198 19168
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 10192 19128 10609 19156
rect 10192 19116 10198 19128
rect 10597 19125 10609 19128
rect 10643 19156 10655 19159
rect 10870 19156 10876 19168
rect 10643 19128 10876 19156
rect 10643 19125 10655 19128
rect 10597 19119 10655 19125
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11808 19156 11836 19255
rect 12253 19227 12311 19233
rect 12253 19193 12265 19227
rect 12299 19224 12311 19227
rect 12912 19224 12940 19255
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 23658 19292 23664 19304
rect 23619 19264 23664 19292
rect 23658 19252 23664 19264
rect 23716 19292 23722 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23716 19264 24133 19292
rect 23716 19252 23722 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24121 19255 24179 19261
rect 14090 19224 14096 19236
rect 12299 19196 12940 19224
rect 14003 19196 14096 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 14090 19184 14096 19196
rect 14148 19224 14154 19236
rect 14553 19227 14611 19233
rect 14553 19224 14565 19227
rect 14148 19196 14565 19224
rect 14148 19184 14154 19196
rect 14553 19193 14565 19196
rect 14599 19193 14611 19227
rect 14553 19187 14611 19193
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 11808 19128 12817 19156
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 13446 19156 13452 19168
rect 13407 19128 13452 19156
rect 12805 19119 12863 19125
rect 13446 19116 13452 19128
rect 13504 19156 13510 19168
rect 13722 19156 13728 19168
rect 13504 19128 13728 19156
rect 13504 19116 13510 19128
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 14182 19156 14188 19168
rect 14143 19128 14188 19156
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 14642 19156 14648 19168
rect 14603 19128 14648 19156
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 15746 19156 15752 19168
rect 15707 19128 15752 19156
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 23845 19159 23903 19165
rect 23845 19125 23857 19159
rect 23891 19156 23903 19159
rect 24762 19156 24768 19168
rect 23891 19128 24768 19156
rect 23891 19125 23903 19128
rect 23845 19119 23903 19125
rect 24762 19116 24768 19128
rect 24820 19116 24826 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 1854 18912 1860 18964
rect 1912 18952 1918 18964
rect 2133 18955 2191 18961
rect 2133 18952 2145 18955
rect 1912 18924 2145 18952
rect 1912 18912 1918 18924
rect 2133 18921 2145 18924
rect 2179 18952 2191 18955
rect 2498 18952 2504 18964
rect 2179 18924 2504 18952
rect 2179 18921 2191 18924
rect 2133 18915 2191 18921
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 3510 18952 3516 18964
rect 3471 18924 3516 18952
rect 3510 18912 3516 18924
rect 3568 18912 3574 18964
rect 4154 18912 4160 18964
rect 4212 18952 4218 18964
rect 4893 18955 4951 18961
rect 4893 18952 4905 18955
rect 4212 18924 4905 18952
rect 4212 18912 4218 18924
rect 4893 18921 4905 18924
rect 4939 18952 4951 18955
rect 5258 18952 5264 18964
rect 4939 18924 5264 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 7558 18912 7564 18964
rect 7616 18952 7622 18964
rect 8110 18952 8116 18964
rect 7616 18924 8116 18952
rect 7616 18912 7622 18924
rect 8110 18912 8116 18924
rect 8168 18912 8174 18964
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 10134 18952 10140 18964
rect 9732 18924 10140 18952
rect 9732 18912 9738 18924
rect 10134 18912 10140 18924
rect 10192 18912 10198 18964
rect 11238 18952 11244 18964
rect 11151 18924 11244 18952
rect 11238 18912 11244 18924
rect 11296 18952 11302 18964
rect 12434 18952 12440 18964
rect 11296 18924 12440 18952
rect 11296 18912 11302 18924
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 13081 18955 13139 18961
rect 13081 18921 13093 18955
rect 13127 18921 13139 18955
rect 13081 18915 13139 18921
rect 2866 18884 2872 18896
rect 2779 18856 2872 18884
rect 2866 18844 2872 18856
rect 2924 18884 2930 18896
rect 3970 18884 3976 18896
rect 2924 18856 3976 18884
rect 2924 18844 2930 18856
rect 3970 18844 3976 18856
rect 4028 18844 4034 18896
rect 5442 18893 5448 18896
rect 5436 18884 5448 18893
rect 5403 18856 5448 18884
rect 5436 18847 5448 18856
rect 5442 18844 5448 18847
rect 5500 18844 5506 18896
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18884 10103 18887
rect 10226 18884 10232 18896
rect 10091 18856 10232 18884
rect 10091 18853 10103 18856
rect 10045 18847 10103 18853
rect 10226 18844 10232 18856
rect 10284 18884 10290 18896
rect 10686 18884 10692 18896
rect 10284 18856 10692 18884
rect 10284 18844 10290 18856
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 10873 18887 10931 18893
rect 10873 18853 10885 18887
rect 10919 18884 10931 18887
rect 11422 18884 11428 18896
rect 10919 18856 11428 18884
rect 10919 18853 10931 18856
rect 10873 18847 10931 18853
rect 11422 18844 11428 18856
rect 11480 18884 11486 18896
rect 12342 18884 12348 18896
rect 11480 18856 12348 18884
rect 11480 18844 11486 18856
rect 12342 18844 12348 18856
rect 12400 18884 12406 18896
rect 13096 18884 13124 18915
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14185 18955 14243 18961
rect 14185 18952 14197 18955
rect 14148 18924 14197 18952
rect 14148 18912 14154 18924
rect 14185 18921 14197 18924
rect 14231 18921 14243 18955
rect 14185 18915 14243 18921
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16669 18955 16727 18961
rect 16669 18952 16681 18955
rect 16632 18924 16681 18952
rect 16632 18912 16638 18924
rect 16669 18921 16681 18924
rect 16715 18921 16727 18955
rect 16669 18915 16727 18921
rect 12400 18856 13124 18884
rect 12400 18844 12406 18856
rect 14458 18844 14464 18896
rect 14516 18884 14522 18896
rect 15286 18884 15292 18896
rect 14516 18856 15292 18884
rect 14516 18844 14522 18856
rect 15286 18844 15292 18856
rect 15344 18884 15350 18896
rect 15534 18887 15592 18893
rect 15534 18884 15546 18887
rect 15344 18856 15546 18884
rect 15344 18844 15350 18856
rect 15534 18853 15546 18856
rect 15580 18853 15592 18887
rect 15534 18847 15592 18853
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4338 18816 4344 18828
rect 4111 18788 4344 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4338 18776 4344 18788
rect 4396 18776 4402 18828
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 7742 18816 7748 18828
rect 7607 18788 7748 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 7742 18776 7748 18788
rect 7800 18816 7806 18828
rect 8021 18819 8079 18825
rect 8021 18816 8033 18819
rect 7800 18788 8033 18816
rect 7800 18776 7806 18788
rect 8021 18785 8033 18788
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 11609 18819 11667 18825
rect 11609 18785 11621 18819
rect 11655 18816 11667 18819
rect 11968 18819 12026 18825
rect 11968 18816 11980 18819
rect 11655 18788 11980 18816
rect 11655 18785 11667 18788
rect 11609 18779 11667 18785
rect 11968 18785 11980 18788
rect 12014 18816 12026 18819
rect 12526 18816 12532 18828
rect 12014 18788 12532 18816
rect 12014 18785 12026 18788
rect 11968 18779 12026 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 2222 18748 2228 18760
rect 2183 18720 2228 18748
rect 2222 18708 2228 18720
rect 2280 18708 2286 18760
rect 2406 18708 2412 18760
rect 2464 18748 2470 18760
rect 2464 18720 2509 18748
rect 2464 18708 2470 18720
rect 4614 18708 4620 18760
rect 4672 18748 4678 18760
rect 5169 18751 5227 18757
rect 5169 18748 5181 18751
rect 4672 18720 5181 18748
rect 4672 18708 4678 18720
rect 5169 18717 5181 18720
rect 5215 18717 5227 18751
rect 5169 18711 5227 18717
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 9398 18748 9404 18760
rect 8343 18720 9404 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 11701 18751 11759 18757
rect 11701 18717 11713 18751
rect 11747 18717 11759 18751
rect 11701 18711 11759 18717
rect 2424 18680 2452 18708
rect 3145 18683 3203 18689
rect 3145 18680 3157 18683
rect 2424 18652 3157 18680
rect 3145 18649 3157 18652
rect 3191 18680 3203 18683
rect 3326 18680 3332 18692
rect 3191 18652 3332 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3326 18640 3332 18652
rect 3384 18640 3390 18692
rect 6822 18640 6828 18692
rect 6880 18680 6886 18692
rect 7101 18683 7159 18689
rect 7101 18680 7113 18683
rect 6880 18652 7113 18680
rect 6880 18640 6886 18652
rect 7101 18649 7113 18652
rect 7147 18649 7159 18683
rect 7650 18680 7656 18692
rect 7611 18652 7656 18680
rect 7101 18643 7159 18649
rect 1670 18612 1676 18624
rect 1631 18584 1676 18612
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 3970 18572 3976 18624
rect 4028 18612 4034 18624
rect 4249 18615 4307 18621
rect 4249 18612 4261 18615
rect 4028 18584 4261 18612
rect 4028 18572 4034 18584
rect 4249 18581 4261 18584
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 6914 18612 6920 18624
rect 6595 18584 6920 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7116 18612 7144 18643
rect 7650 18640 7656 18652
rect 7708 18640 7714 18692
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 9766 18680 9772 18692
rect 9723 18652 9772 18680
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 9214 18612 9220 18624
rect 7116 18584 9220 18612
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 11716 18612 11744 18711
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 13504 18720 15301 18748
rect 13504 18708 13510 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 11882 18612 11888 18624
rect 11716 18584 11888 18612
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 14642 18612 14648 18624
rect 13872 18584 14648 18612
rect 13872 18572 13878 18584
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 15304 18612 15332 18711
rect 15654 18612 15660 18624
rect 15304 18584 15660 18612
rect 15654 18572 15660 18584
rect 15712 18572 15718 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2041 18411 2099 18417
rect 2041 18408 2053 18411
rect 1728 18380 2053 18408
rect 1728 18368 1734 18380
rect 2041 18377 2053 18380
rect 2087 18377 2099 18411
rect 2041 18371 2099 18377
rect 1765 18343 1823 18349
rect 1765 18309 1777 18343
rect 1811 18340 1823 18343
rect 1854 18340 1860 18352
rect 1811 18312 1860 18340
rect 1811 18309 1823 18312
rect 1765 18303 1823 18309
rect 1854 18300 1860 18312
rect 1912 18300 1918 18352
rect 2056 18272 2084 18371
rect 3326 18368 3332 18420
rect 3384 18408 3390 18420
rect 3605 18411 3663 18417
rect 3605 18408 3617 18411
rect 3384 18380 3617 18408
rect 3384 18368 3390 18380
rect 3605 18377 3617 18380
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 4249 18411 4307 18417
rect 4249 18377 4261 18411
rect 4295 18408 4307 18411
rect 5442 18408 5448 18420
rect 4295 18380 5448 18408
rect 4295 18377 4307 18380
rect 4249 18371 4307 18377
rect 5442 18368 5448 18380
rect 5500 18408 5506 18420
rect 6086 18408 6092 18420
rect 5500 18380 6092 18408
rect 5500 18368 5506 18380
rect 6086 18368 6092 18380
rect 6144 18368 6150 18420
rect 8202 18408 8208 18420
rect 8163 18380 8208 18408
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 9122 18408 9128 18420
rect 9083 18380 9128 18408
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 10226 18408 10232 18420
rect 10187 18380 10232 18408
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 12253 18411 12311 18417
rect 12253 18377 12265 18411
rect 12299 18408 12311 18411
rect 12526 18408 12532 18420
rect 12299 18380 12532 18408
rect 12299 18377 12311 18380
rect 12253 18371 12311 18377
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 15105 18411 15163 18417
rect 15105 18377 15117 18411
rect 15151 18408 15163 18411
rect 15286 18408 15292 18420
rect 15151 18380 15292 18408
rect 15151 18377 15163 18380
rect 15105 18371 15163 18377
rect 15286 18368 15292 18380
rect 15344 18408 15350 18420
rect 16025 18411 16083 18417
rect 16025 18408 16037 18411
rect 15344 18380 16037 18408
rect 15344 18368 15350 18380
rect 16025 18377 16037 18380
rect 16071 18377 16083 18411
rect 16025 18371 16083 18377
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 2056 18244 2237 18272
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 5166 18272 5172 18284
rect 4120 18244 5172 18272
rect 4120 18232 4126 18244
rect 5166 18232 5172 18244
rect 5224 18232 5230 18284
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 5460 18272 5488 18368
rect 8849 18343 8907 18349
rect 8849 18309 8861 18343
rect 8895 18340 8907 18343
rect 9398 18340 9404 18352
rect 8895 18312 9404 18340
rect 8895 18309 8907 18312
rect 8849 18303 8907 18309
rect 9398 18300 9404 18312
rect 9456 18300 9462 18352
rect 15654 18340 15660 18352
rect 15615 18312 15660 18340
rect 15654 18300 15660 18312
rect 15712 18300 15718 18352
rect 11238 18272 11244 18284
rect 5399 18244 5488 18272
rect 11199 18244 11244 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 11422 18272 11428 18284
rect 11383 18244 11428 18272
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 2492 18207 2550 18213
rect 2492 18173 2504 18207
rect 2538 18204 2550 18207
rect 2866 18204 2872 18216
rect 2538 18176 2872 18204
rect 2538 18173 2550 18176
rect 2492 18167 2550 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 6822 18204 6828 18216
rect 6564 18176 6828 18204
rect 4617 18139 4675 18145
rect 4617 18105 4629 18139
rect 4663 18136 4675 18139
rect 4663 18108 5120 18136
rect 4663 18105 4675 18108
rect 4617 18099 4675 18105
rect 5092 18080 5120 18108
rect 4706 18068 4712 18080
rect 4667 18040 4712 18068
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 6564 18077 6592 18176
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 9180 18176 9321 18204
rect 9180 18164 9186 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9861 18207 9919 18213
rect 9861 18173 9873 18207
rect 9907 18204 9919 18207
rect 10318 18204 10324 18216
rect 9907 18176 10324 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10318 18164 10324 18176
rect 10376 18204 10382 18216
rect 11054 18204 11060 18216
rect 10376 18176 11060 18204
rect 10376 18164 10382 18176
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 13446 18164 13452 18216
rect 13504 18204 13510 18216
rect 13725 18207 13783 18213
rect 13725 18204 13737 18207
rect 13504 18176 13737 18204
rect 13504 18164 13510 18176
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 7070 18139 7128 18145
rect 7070 18136 7082 18139
rect 6972 18108 7082 18136
rect 6972 18096 6978 18108
rect 7070 18105 7082 18108
rect 7116 18105 7128 18139
rect 7070 18099 7128 18105
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 11149 18139 11207 18145
rect 11149 18136 11161 18139
rect 10735 18108 11161 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 11149 18105 11161 18108
rect 11195 18136 11207 18139
rect 12437 18139 12495 18145
rect 12437 18136 12449 18139
rect 11195 18108 12449 18136
rect 11195 18105 11207 18108
rect 11149 18099 11207 18105
rect 12437 18105 12449 18108
rect 12483 18105 12495 18139
rect 12437 18099 12495 18105
rect 5813 18071 5871 18077
rect 5813 18037 5825 18071
rect 5859 18068 5871 18071
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 5859 18040 6561 18068
rect 5859 18037 5871 18040
rect 5813 18031 5871 18037
rect 6549 18037 6561 18040
rect 6595 18037 6607 18071
rect 6549 18031 6607 18037
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 9493 18071 9551 18077
rect 9493 18068 9505 18071
rect 8352 18040 9505 18068
rect 8352 18028 8358 18040
rect 9493 18037 9505 18040
rect 9539 18037 9551 18071
rect 10778 18068 10784 18080
rect 10739 18040 10784 18068
rect 9493 18031 9551 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11882 18068 11888 18080
rect 11843 18040 11888 18068
rect 11882 18028 11888 18040
rect 11940 18068 11946 18080
rect 13556 18077 13584 18176
rect 13725 18173 13737 18176
rect 13771 18173 13783 18207
rect 13725 18167 13783 18173
rect 15194 18164 15200 18216
rect 15252 18204 15258 18216
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 15252 18176 16221 18204
rect 15252 18164 15258 18176
rect 16209 18173 16221 18176
rect 16255 18204 16267 18207
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16255 18176 16773 18204
rect 16255 18173 16267 18176
rect 16209 18167 16267 18173
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 13998 18145 14004 18148
rect 13992 18136 14004 18145
rect 13959 18108 14004 18136
rect 13992 18099 14004 18108
rect 13998 18096 14004 18099
rect 14056 18096 14062 18148
rect 13541 18071 13599 18077
rect 13541 18068 13553 18071
rect 11940 18040 13553 18068
rect 11940 18028 11946 18040
rect 13541 18037 13553 18040
rect 13587 18037 13599 18071
rect 16390 18068 16396 18080
rect 16351 18040 16396 18068
rect 13541 18031 13599 18037
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2222 17864 2228 17876
rect 2183 17836 2228 17864
rect 2222 17824 2228 17836
rect 2280 17864 2286 17876
rect 3237 17867 3295 17873
rect 3237 17864 3249 17867
rect 2280 17836 3249 17864
rect 2280 17824 2286 17836
rect 3237 17833 3249 17836
rect 3283 17833 3295 17867
rect 3237 17827 3295 17833
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 4062 17864 4068 17876
rect 3927 17836 4068 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 6086 17864 6092 17876
rect 6047 17836 6092 17864
rect 6086 17824 6092 17836
rect 6144 17824 6150 17876
rect 7558 17864 7564 17876
rect 7519 17836 7564 17864
rect 7558 17824 7564 17836
rect 7616 17824 7622 17876
rect 7742 17864 7748 17876
rect 7703 17836 7748 17864
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 10229 17867 10287 17873
rect 10229 17864 10241 17867
rect 10192 17836 10241 17864
rect 10192 17824 10198 17836
rect 10229 17833 10241 17836
rect 10275 17833 10287 17867
rect 10229 17827 10287 17833
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 15102 17864 15108 17876
rect 14415 17836 15108 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 15289 17867 15347 17873
rect 15289 17833 15301 17867
rect 15335 17833 15347 17867
rect 15289 17827 15347 17833
rect 1857 17799 1915 17805
rect 1857 17765 1869 17799
rect 1903 17796 1915 17799
rect 2406 17796 2412 17808
rect 1903 17768 2412 17796
rect 1903 17765 1915 17768
rect 1857 17759 1915 17765
rect 2406 17756 2412 17768
rect 2464 17756 2470 17808
rect 2685 17799 2743 17805
rect 2685 17765 2697 17799
rect 2731 17796 2743 17799
rect 3142 17796 3148 17808
rect 2731 17768 3148 17796
rect 2731 17765 2743 17768
rect 2685 17759 2743 17765
rect 3142 17756 3148 17768
rect 3200 17796 3206 17808
rect 4154 17796 4160 17808
rect 3200 17768 4160 17796
rect 3200 17756 3206 17768
rect 4154 17756 4160 17768
rect 4212 17756 4218 17808
rect 7285 17799 7343 17805
rect 7285 17765 7297 17799
rect 7331 17796 7343 17799
rect 7926 17796 7932 17808
rect 7331 17768 7932 17796
rect 7331 17765 7343 17768
rect 7285 17759 7343 17765
rect 7926 17756 7932 17768
rect 7984 17756 7990 17808
rect 10870 17756 10876 17808
rect 10928 17796 10934 17808
rect 11026 17799 11084 17805
rect 11026 17796 11038 17799
rect 10928 17768 11038 17796
rect 10928 17756 10934 17768
rect 11026 17765 11038 17768
rect 11072 17765 11084 17799
rect 11026 17759 11084 17765
rect 2590 17728 2596 17740
rect 2551 17700 2596 17728
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 4982 17737 4988 17740
rect 4976 17728 4988 17737
rect 4943 17700 4988 17728
rect 4976 17691 4988 17700
rect 4982 17688 4988 17691
rect 5040 17688 5046 17740
rect 8110 17728 8116 17740
rect 8071 17700 8116 17728
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 9858 17728 9864 17740
rect 9723 17700 9864 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 9858 17688 9864 17700
rect 9916 17688 9922 17740
rect 11882 17728 11888 17740
rect 10796 17700 11888 17728
rect 2866 17660 2872 17672
rect 2827 17632 2872 17660
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 4614 17620 4620 17672
rect 4672 17660 4678 17672
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 4672 17632 4721 17660
rect 4672 17620 4678 17632
rect 4709 17629 4721 17632
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7524 17632 8217 17660
rect 7524 17620 7530 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8386 17660 8392 17672
rect 8347 17632 8392 17660
rect 8205 17623 8263 17629
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 10686 17660 10692 17672
rect 9272 17632 10692 17660
rect 9272 17620 9278 17632
rect 10686 17620 10692 17632
rect 10744 17660 10750 17672
rect 10796 17669 10824 17700
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14185 17731 14243 17737
rect 14185 17728 14197 17731
rect 13964 17700 14197 17728
rect 13964 17688 13970 17700
rect 14185 17697 14197 17700
rect 14231 17728 14243 17731
rect 15304 17728 15332 17827
rect 14231 17700 15332 17728
rect 15657 17731 15715 17737
rect 14231 17697 14243 17700
rect 14185 17691 14243 17697
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 16482 17728 16488 17740
rect 15703 17700 16488 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 10781 17663 10839 17669
rect 10781 17660 10793 17663
rect 10744 17632 10793 17660
rect 10744 17620 10750 17632
rect 10781 17629 10793 17632
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15672 17660 15700 17691
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 16850 17728 16856 17740
rect 16811 17700 16856 17728
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 17862 17728 17868 17740
rect 17823 17700 17868 17728
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 14608 17632 15700 17660
rect 15749 17663 15807 17669
rect 14608 17620 14614 17632
rect 15749 17629 15761 17663
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 1394 17552 1400 17604
rect 1452 17592 1458 17604
rect 3050 17592 3056 17604
rect 1452 17564 3056 17592
rect 1452 17552 1458 17564
rect 3050 17552 3056 17564
rect 3108 17552 3114 17604
rect 13817 17595 13875 17601
rect 13817 17561 13829 17595
rect 13863 17592 13875 17595
rect 13998 17592 14004 17604
rect 13863 17564 14004 17592
rect 13863 17561 13875 17564
rect 13817 17555 13875 17561
rect 13998 17552 14004 17564
rect 14056 17592 14062 17604
rect 15286 17592 15292 17604
rect 14056 17564 15292 17592
rect 14056 17552 14062 17564
rect 15286 17552 15292 17564
rect 15344 17552 15350 17604
rect 4338 17524 4344 17536
rect 4299 17496 4344 17524
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 4890 17484 4896 17536
rect 4948 17524 4954 17536
rect 6914 17524 6920 17536
rect 4948 17496 6920 17524
rect 4948 17484 4954 17496
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 8754 17524 8760 17536
rect 8715 17496 8760 17524
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 9824 17496 9873 17524
rect 9824 17484 9830 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 9861 17487 9919 17493
rect 11054 17484 11060 17536
rect 11112 17524 11118 17536
rect 12066 17524 12072 17536
rect 11112 17496 12072 17524
rect 11112 17484 11118 17496
rect 12066 17484 12072 17496
rect 12124 17524 12130 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 12124 17496 12173 17524
rect 12124 17484 12130 17496
rect 12161 17493 12173 17496
rect 12207 17493 12219 17527
rect 12161 17487 12219 17493
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 15013 17527 15071 17533
rect 15013 17524 15025 17527
rect 14792 17496 15025 17524
rect 14792 17484 14798 17496
rect 15013 17493 15025 17496
rect 15059 17524 15071 17527
rect 15764 17524 15792 17623
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 15896 17632 15941 17660
rect 15896 17620 15902 17632
rect 17034 17524 17040 17536
rect 15059 17496 15792 17524
rect 16995 17496 17040 17524
rect 15059 17493 15071 17496
rect 15013 17487 15071 17493
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2682 17320 2688 17332
rect 2643 17292 2688 17320
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 3142 17320 3148 17332
rect 3103 17292 3148 17320
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 3878 17320 3884 17332
rect 3839 17292 3884 17320
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 4249 17323 4307 17329
rect 4249 17289 4261 17323
rect 4295 17320 4307 17323
rect 4890 17320 4896 17332
rect 4295 17292 4896 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 4890 17280 4896 17292
rect 4948 17280 4954 17332
rect 7466 17320 7472 17332
rect 7427 17292 7472 17320
rect 7466 17280 7472 17292
rect 7524 17280 7530 17332
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 8018 17320 8024 17332
rect 7699 17292 8024 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 8220 17292 10609 17320
rect 2317 17255 2375 17261
rect 2317 17221 2329 17255
rect 2363 17252 2375 17255
rect 2590 17252 2596 17264
rect 2363 17224 2596 17252
rect 2363 17221 2375 17224
rect 2317 17215 2375 17221
rect 2590 17212 2596 17224
rect 2648 17212 2654 17264
rect 3896 17184 3924 17280
rect 5721 17255 5779 17261
rect 5721 17252 5733 17255
rect 4816 17224 5733 17252
rect 4816 17196 4844 17224
rect 5721 17221 5733 17224
rect 5767 17221 5779 17255
rect 5721 17215 5779 17221
rect 4798 17184 4804 17196
rect 1412 17156 3924 17184
rect 4759 17156 4804 17184
rect 1412 17125 1440 17156
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 4890 17144 4896 17196
rect 4948 17184 4954 17196
rect 8220 17193 8248 17292
rect 10597 17289 10609 17292
rect 10643 17320 10655 17323
rect 10962 17320 10968 17332
rect 10643 17292 10968 17320
rect 10643 17289 10655 17292
rect 10597 17283 10655 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 13906 17320 13912 17332
rect 13867 17292 13912 17320
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 14826 17320 14832 17332
rect 14231 17292 14832 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 14826 17280 14832 17292
rect 14884 17280 14890 17332
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 16393 17323 16451 17329
rect 16393 17320 16405 17323
rect 15344 17292 16405 17320
rect 15344 17280 15350 17292
rect 16393 17289 16405 17292
rect 16439 17289 16451 17323
rect 16393 17283 16451 17289
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 16945 17323 17003 17329
rect 16945 17320 16957 17323
rect 16908 17292 16957 17320
rect 16908 17280 16914 17292
rect 16945 17289 16957 17292
rect 16991 17289 17003 17323
rect 16945 17283 17003 17289
rect 8386 17212 8392 17264
rect 8444 17252 8450 17264
rect 8665 17255 8723 17261
rect 8665 17252 8677 17255
rect 8444 17224 8677 17252
rect 8444 17212 8450 17224
rect 8665 17221 8677 17224
rect 8711 17221 8723 17255
rect 9122 17252 9128 17264
rect 9083 17224 9128 17252
rect 8665 17215 8723 17221
rect 9122 17212 9128 17224
rect 9180 17252 9186 17264
rect 12437 17255 12495 17261
rect 9180 17224 9260 17252
rect 9180 17212 9186 17224
rect 9232 17193 9260 17224
rect 12437 17221 12449 17255
rect 12483 17252 12495 17255
rect 13814 17252 13820 17264
rect 12483 17224 13820 17252
rect 12483 17221 12495 17224
rect 12437 17215 12495 17221
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 13998 17212 14004 17264
rect 14056 17212 14062 17264
rect 14550 17252 14556 17264
rect 14511 17224 14556 17252
rect 14550 17212 14556 17224
rect 14608 17212 14614 17264
rect 18230 17252 18236 17264
rect 18191 17224 18236 17252
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 19334 17212 19340 17264
rect 19392 17252 19398 17264
rect 20254 17252 20260 17264
rect 19392 17224 20260 17252
rect 19392 17212 19398 17224
rect 20254 17212 20260 17224
rect 20312 17212 20318 17264
rect 7193 17187 7251 17193
rect 4948 17156 4993 17184
rect 4948 17144 4954 17156
rect 7193 17153 7205 17187
rect 7239 17184 7251 17187
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 7239 17156 8217 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12860 17156 13093 17184
rect 12860 17144 12866 17156
rect 13081 17153 13093 17156
rect 13127 17184 13139 17187
rect 14016 17184 14044 17212
rect 13127 17156 14044 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 1397 17079 1455 17085
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2501 17119 2559 17125
rect 2501 17116 2513 17119
rect 2004 17088 2513 17116
rect 2004 17076 2010 17088
rect 2501 17085 2513 17088
rect 2547 17116 2559 17119
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 2547 17088 3433 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 3421 17085 3433 17088
rect 3467 17085 3479 17119
rect 4706 17116 4712 17128
rect 4667 17088 4712 17116
rect 3421 17079 3479 17085
rect 4706 17076 4712 17088
rect 4764 17116 4770 17128
rect 6089 17119 6147 17125
rect 6089 17116 6101 17119
rect 4764 17088 6101 17116
rect 4764 17076 4770 17088
rect 6089 17085 6101 17088
rect 6135 17085 6147 17119
rect 6089 17079 6147 17085
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 9490 17125 9496 17128
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 7984 17088 8125 17116
rect 7984 17076 7990 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 9484 17116 9496 17125
rect 9451 17088 9496 17116
rect 8113 17079 8171 17085
rect 9484 17079 9496 17088
rect 9490 17076 9496 17079
rect 9548 17076 9554 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 11808 17088 12909 17116
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17048 6699 17051
rect 8018 17048 8024 17060
rect 6687 17020 8024 17048
rect 6687 17017 6699 17020
rect 6641 17011 6699 17017
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 4338 16980 4344 16992
rect 4299 16952 4344 16980
rect 4338 16940 4344 16952
rect 4396 16940 4402 16992
rect 4614 16940 4620 16992
rect 4672 16980 4678 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 4672 16952 5365 16980
rect 4672 16940 4678 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 5353 16943 5411 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 10744 16952 11253 16980
rect 10744 16940 10750 16952
rect 11241 16949 11253 16952
rect 11287 16949 11299 16983
rect 11241 16943 11299 16949
rect 11698 16940 11704 16992
rect 11756 16980 11762 16992
rect 11808 16989 11836 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 14001 17079 14059 17085
rect 14844 17088 15025 17116
rect 12158 17008 12164 17060
rect 12216 17048 12222 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 12216 17020 12265 17048
rect 12216 17008 12222 17020
rect 12253 17017 12265 17020
rect 12299 17048 12311 17051
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 12299 17020 12817 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 13446 17048 13452 17060
rect 13407 17020 13452 17048
rect 12805 17011 12863 17017
rect 13446 17008 13452 17020
rect 13504 17048 13510 17060
rect 14016 17048 14044 17079
rect 13504 17020 14044 17048
rect 13504 17008 13510 17020
rect 14844 16992 14872 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 18046 17116 18052 17128
rect 18007 17088 18052 17116
rect 15013 17079 15071 17085
rect 18046 17076 18052 17088
rect 18104 17116 18110 17128
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18104 17088 18521 17116
rect 18104 17076 18110 17088
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 15280 17051 15338 17057
rect 15280 17017 15292 17051
rect 15326 17048 15338 17051
rect 15838 17048 15844 17060
rect 15326 17020 15844 17048
rect 15326 17017 15338 17020
rect 15280 17011 15338 17017
rect 15838 17008 15844 17020
rect 15896 17008 15902 17060
rect 11793 16983 11851 16989
rect 11793 16980 11805 16983
rect 11756 16952 11805 16980
rect 11756 16940 11762 16952
rect 11793 16949 11805 16952
rect 11839 16949 11851 16983
rect 14826 16980 14832 16992
rect 14787 16952 14832 16980
rect 11793 16943 11851 16949
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1486 16736 1492 16788
rect 1544 16776 1550 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1544 16748 1593 16776
rect 1544 16736 1550 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 1581 16739 1639 16745
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 2556 16748 2697 16776
rect 2556 16736 2562 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 2685 16739 2743 16745
rect 3050 16736 3056 16788
rect 3108 16776 3114 16788
rect 3145 16779 3203 16785
rect 3145 16776 3157 16779
rect 3108 16748 3157 16776
rect 3108 16736 3114 16748
rect 3145 16745 3157 16748
rect 3191 16745 3203 16779
rect 3602 16776 3608 16788
rect 3563 16748 3608 16776
rect 3145 16739 3203 16745
rect 3602 16736 3608 16748
rect 3660 16736 3666 16788
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3936 16748 4077 16776
rect 3936 16736 3942 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4065 16739 4123 16745
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5077 16779 5135 16785
rect 5077 16776 5089 16779
rect 5040 16748 5089 16776
rect 5040 16736 5046 16748
rect 5077 16745 5089 16748
rect 5123 16745 5135 16779
rect 5077 16739 5135 16745
rect 6365 16779 6423 16785
rect 6365 16745 6377 16779
rect 6411 16776 6423 16779
rect 6546 16776 6552 16788
rect 6411 16748 6552 16776
rect 6411 16745 6423 16748
rect 6365 16739 6423 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16776 9367 16779
rect 9490 16776 9496 16788
rect 9355 16748 9496 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 9861 16779 9919 16785
rect 9861 16745 9873 16779
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16776 10747 16779
rect 10870 16776 10876 16788
rect 10735 16748 10876 16776
rect 10735 16745 10747 16748
rect 10689 16739 10747 16745
rect 3620 16708 3648 16736
rect 2516 16680 3648 16708
rect 5997 16711 6055 16717
rect 2516 16649 2544 16680
rect 5997 16677 6009 16711
rect 6043 16708 6055 16711
rect 6917 16711 6975 16717
rect 6917 16708 6929 16711
rect 6043 16680 6929 16708
rect 6043 16677 6055 16680
rect 5997 16671 6055 16677
rect 6917 16677 6929 16680
rect 6963 16708 6975 16711
rect 7098 16708 7104 16720
rect 6963 16680 7104 16708
rect 6963 16677 6975 16680
rect 6917 16671 6975 16677
rect 7098 16668 7104 16680
rect 7156 16668 7162 16720
rect 7837 16711 7895 16717
rect 7837 16677 7849 16711
rect 7883 16708 7895 16711
rect 8110 16708 8116 16720
rect 7883 16680 8116 16708
rect 7883 16677 7895 16680
rect 7837 16671 7895 16677
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 8481 16711 8539 16717
rect 8481 16708 8493 16711
rect 8220 16680 8493 16708
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 2501 16643 2559 16649
rect 1443 16612 1716 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1688 16436 1716 16612
rect 2501 16609 2513 16643
rect 2547 16609 2559 16643
rect 4430 16640 4436 16652
rect 4391 16612 4436 16640
rect 2501 16603 2559 16609
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 4706 16640 4712 16652
rect 4571 16612 4712 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 6822 16640 6828 16652
rect 5675 16612 6828 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 8220 16640 8248 16680
rect 8481 16677 8493 16680
rect 8527 16677 8539 16711
rect 8481 16671 8539 16677
rect 9766 16668 9772 16720
rect 9824 16708 9830 16720
rect 9876 16708 9904 16739
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12161 16779 12219 16785
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 12526 16776 12532 16788
rect 12207 16748 12532 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 13449 16779 13507 16785
rect 13449 16745 13461 16779
rect 13495 16776 13507 16779
rect 14734 16776 14740 16788
rect 13495 16748 14740 16776
rect 13495 16745 13507 16748
rect 13449 16739 13507 16745
rect 14734 16736 14740 16748
rect 14792 16736 14798 16788
rect 15470 16776 15476 16788
rect 15431 16748 15476 16776
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 15838 16776 15844 16788
rect 15799 16748 15844 16776
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 17954 16776 17960 16788
rect 17915 16748 17960 16776
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 9824 16680 9904 16708
rect 9824 16668 9830 16680
rect 10962 16668 10968 16720
rect 11020 16717 11026 16720
rect 11020 16711 11084 16717
rect 11020 16677 11038 16711
rect 11072 16677 11084 16711
rect 11020 16671 11084 16677
rect 15105 16711 15163 16717
rect 15105 16677 15117 16711
rect 15151 16708 15163 16711
rect 15856 16708 15884 16736
rect 15151 16680 15884 16708
rect 15151 16677 15163 16680
rect 15105 16671 15163 16677
rect 11020 16668 11026 16671
rect 8386 16640 8392 16652
rect 7524 16612 8248 16640
rect 8347 16612 8392 16640
rect 7524 16600 7530 16612
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 9858 16600 9864 16652
rect 9916 16640 9922 16652
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 9916 16612 10241 16640
rect 9916 16600 9922 16612
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 13817 16643 13875 16649
rect 13817 16640 13829 16643
rect 10229 16603 10287 16609
rect 13740 16612 13829 16640
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16572 2375 16575
rect 2866 16572 2872 16584
rect 2363 16544 2872 16572
rect 2363 16541 2375 16544
rect 2317 16535 2375 16541
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3602 16532 3608 16584
rect 3660 16572 3666 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 3660 16544 4629 16572
rect 3660 16532 3666 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 7009 16575 7067 16581
rect 7009 16572 7021 16575
rect 6604 16544 7021 16572
rect 6604 16532 6610 16544
rect 7009 16541 7021 16544
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 8665 16575 8723 16581
rect 8665 16541 8677 16575
rect 8711 16572 8723 16575
rect 9490 16572 9496 16584
rect 8711 16544 9496 16572
rect 8711 16541 8723 16544
rect 8665 16535 8723 16541
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 10686 16532 10692 16584
rect 10744 16572 10750 16584
rect 10781 16575 10839 16581
rect 10781 16572 10793 16575
rect 10744 16544 10793 16572
rect 10744 16532 10750 16544
rect 10781 16541 10793 16544
rect 10827 16541 10839 16575
rect 10781 16535 10839 16541
rect 13538 16532 13544 16584
rect 13596 16572 13602 16584
rect 13740 16572 13768 16612
rect 13817 16609 13829 16612
rect 13863 16609 13875 16643
rect 14550 16640 14556 16652
rect 13817 16603 13875 16609
rect 14108 16612 14556 16640
rect 14108 16581 14136 16612
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 16850 16649 16856 16652
rect 16844 16603 16856 16649
rect 16908 16640 16914 16652
rect 16908 16612 16944 16640
rect 16850 16600 16856 16603
rect 16908 16600 16914 16612
rect 13596 16544 13768 16572
rect 13909 16575 13967 16581
rect 13596 16532 13602 16544
rect 13909 16541 13921 16575
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 13924 16504 13952 16535
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 16577 16575 16635 16581
rect 16577 16572 16589 16575
rect 16356 16544 16589 16572
rect 16356 16532 16362 16544
rect 16577 16541 16589 16544
rect 16623 16541 16635 16575
rect 16577 16535 16635 16541
rect 13464 16476 13952 16504
rect 13464 16448 13492 16476
rect 4154 16436 4160 16448
rect 1688 16408 4160 16436
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 13446 16436 13452 16448
rect 13403 16408 13452 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 3234 16192 3240 16244
rect 3292 16232 3298 16244
rect 4798 16232 4804 16244
rect 3292 16204 4804 16232
rect 3292 16192 3298 16204
rect 4798 16192 4804 16204
rect 4856 16232 4862 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 4856 16204 6561 16232
rect 4856 16192 4862 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 6914 16232 6920 16244
rect 6875 16204 6920 16232
rect 6549 16195 6607 16201
rect 14 16124 20 16176
rect 72 16164 78 16176
rect 2961 16167 3019 16173
rect 2961 16164 2973 16167
rect 72 16136 2973 16164
rect 72 16124 78 16136
rect 2961 16133 2973 16136
rect 3007 16133 3019 16167
rect 6564 16164 6592 16195
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 7466 16192 7472 16244
rect 7524 16232 7530 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7524 16204 8033 16232
rect 7524 16192 7530 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9490 16232 9496 16244
rect 9079 16204 9496 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 11238 16232 11244 16244
rect 11199 16204 11244 16232
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 15565 16235 15623 16241
rect 15565 16201 15577 16235
rect 15611 16232 15623 16235
rect 15838 16232 15844 16244
rect 15611 16204 15844 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16577 16235 16635 16241
rect 16577 16201 16589 16235
rect 16623 16232 16635 16235
rect 16850 16232 16856 16244
rect 16623 16204 16856 16232
rect 16623 16201 16635 16204
rect 16577 16195 16635 16201
rect 16850 16192 16856 16204
rect 16908 16192 16914 16244
rect 6825 16167 6883 16173
rect 6825 16164 6837 16167
rect 6564 16136 6837 16164
rect 2961 16127 3019 16133
rect 6825 16133 6837 16136
rect 6871 16133 6883 16167
rect 6825 16127 6883 16133
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16065 2283 16099
rect 2225 16059 2283 16065
rect 2240 16028 2268 16059
rect 2685 16031 2743 16037
rect 2685 16028 2697 16031
rect 2240 16000 2697 16028
rect 2685 15997 2697 16000
rect 2731 15997 2743 16031
rect 2685 15991 2743 15997
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2590 15960 2596 15972
rect 1995 15932 2596 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2590 15920 2596 15932
rect 2648 15920 2654 15972
rect 2700 15892 2728 15991
rect 2976 15960 3004 16127
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11609 16167 11667 16173
rect 11609 16164 11621 16167
rect 11112 16136 11621 16164
rect 11112 16124 11118 16136
rect 11609 16133 11621 16136
rect 11655 16133 11667 16167
rect 11609 16127 11667 16133
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 16209 16167 16267 16173
rect 16209 16164 16221 16167
rect 15344 16136 16221 16164
rect 15344 16124 15350 16136
rect 16209 16133 16221 16136
rect 16255 16164 16267 16167
rect 18233 16167 18291 16173
rect 18233 16164 18245 16167
rect 16255 16136 18245 16164
rect 16255 16133 16267 16136
rect 16209 16127 16267 16133
rect 18233 16133 18245 16136
rect 18279 16133 18291 16167
rect 18233 16127 18291 16133
rect 3602 16056 3608 16108
rect 3660 16096 3666 16108
rect 3697 16099 3755 16105
rect 3697 16096 3709 16099
rect 3660 16068 3709 16096
rect 3660 16056 3666 16068
rect 3697 16065 3709 16068
rect 3743 16065 3755 16099
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 3697 16059 3755 16065
rect 5276 16068 5733 16096
rect 3050 15988 3056 16040
rect 3108 16028 3114 16040
rect 3510 16028 3516 16040
rect 3108 16000 3516 16028
rect 3108 15988 3114 16000
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 5276 15972 5304 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 6273 16099 6331 16105
rect 6273 16065 6285 16099
rect 6319 16096 6331 16099
rect 7561 16099 7619 16105
rect 7561 16096 7573 16099
rect 6319 16068 7573 16096
rect 6319 16065 6331 16068
rect 6273 16059 6331 16065
rect 7561 16065 7573 16068
rect 7607 16096 7619 16099
rect 7742 16096 7748 16108
rect 7607 16068 7748 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 8444 16068 8493 16096
rect 8444 16056 8450 16068
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 10042 16096 10048 16108
rect 9447 16068 10048 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 12526 16056 12532 16108
rect 12584 16096 12590 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12584 16068 13001 16096
rect 12584 16056 12590 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 6454 16028 6460 16040
rect 5675 16000 6460 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 6871 16000 7389 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7377 15997 7389 16000
rect 7423 16028 7435 16031
rect 8754 16028 8760 16040
rect 7423 16000 8760 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 8754 15988 8760 16000
rect 8812 15988 8818 16040
rect 9306 15988 9312 16040
rect 9364 16028 9370 16040
rect 9861 16031 9919 16037
rect 9861 16028 9873 16031
rect 9364 16000 9873 16028
rect 9364 15988 9370 16000
rect 9861 15997 9873 16000
rect 9907 15997 9919 16031
rect 9861 15991 9919 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11514 16028 11520 16040
rect 11103 16000 11520 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 12802 16028 12808 16040
rect 12299 16000 12808 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 12802 15988 12808 16000
rect 12860 15988 12866 16040
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 14016 16000 14197 16028
rect 3234 15960 3240 15972
rect 2976 15932 3240 15960
rect 3234 15920 3240 15932
rect 3292 15960 3298 15972
rect 3605 15963 3663 15969
rect 3605 15960 3617 15963
rect 3292 15932 3617 15960
rect 3292 15920 3298 15932
rect 3605 15929 3617 15932
rect 3651 15929 3663 15963
rect 3605 15923 3663 15929
rect 5077 15963 5135 15969
rect 5077 15929 5089 15963
rect 5123 15960 5135 15963
rect 5258 15960 5264 15972
rect 5123 15932 5264 15960
rect 5123 15929 5135 15932
rect 5077 15923 5135 15929
rect 5258 15920 5264 15932
rect 5316 15920 5322 15972
rect 9766 15920 9772 15972
rect 9824 15960 9830 15972
rect 9953 15963 10011 15969
rect 9953 15960 9965 15963
rect 9824 15932 9965 15960
rect 9824 15920 9830 15932
rect 9953 15929 9965 15932
rect 9999 15929 10011 15963
rect 9953 15923 10011 15929
rect 2866 15892 2872 15904
rect 2700 15864 2872 15892
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 3142 15892 3148 15904
rect 3103 15864 3148 15892
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3694 15852 3700 15904
rect 3752 15892 3758 15904
rect 4157 15895 4215 15901
rect 4157 15892 4169 15895
rect 3752 15864 4169 15892
rect 3752 15852 3758 15864
rect 4157 15861 4169 15864
rect 4203 15892 4215 15895
rect 4430 15892 4436 15904
rect 4203 15864 4436 15892
rect 4203 15861 4215 15864
rect 4157 15855 4215 15861
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15892 4675 15895
rect 4706 15892 4712 15904
rect 4663 15864 4712 15892
rect 4663 15861 4675 15864
rect 4617 15855 4675 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 5537 15895 5595 15901
rect 5537 15861 5549 15895
rect 5583 15892 5595 15895
rect 5994 15892 6000 15904
rect 5583 15864 6000 15892
rect 5583 15861 5595 15864
rect 5537 15855 5595 15861
rect 5994 15852 6000 15864
rect 6052 15852 6058 15904
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7282 15892 7288 15904
rect 6972 15864 7288 15892
rect 6972 15852 6978 15864
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 9490 15892 9496 15904
rect 9451 15864 9496 15892
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 12894 15892 12900 15904
rect 12492 15864 12537 15892
rect 12855 15864 12900 15892
rect 12492 15852 12498 15864
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 13538 15892 13544 15904
rect 13499 15864 13544 15892
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14016 15901 14044 16000
rect 14185 15997 14197 16000
rect 14231 16028 14243 16031
rect 14826 16028 14832 16040
rect 14231 16000 14832 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 16028 18110 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18104 16000 18521 16028
rect 18104 15988 18110 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 19058 16028 19064 16040
rect 19019 16000 19064 16028
rect 18509 15991 18567 15997
rect 19058 15988 19064 16000
rect 19116 16028 19122 16040
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19116 16000 19533 16028
rect 19116 15988 19122 16000
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 19521 15991 19579 15997
rect 14452 15963 14510 15969
rect 14452 15929 14464 15963
rect 14498 15960 14510 15963
rect 14550 15960 14556 15972
rect 14498 15932 14556 15960
rect 14498 15929 14510 15932
rect 14452 15923 14510 15929
rect 14550 15920 14556 15932
rect 14608 15920 14614 15972
rect 14001 15895 14059 15901
rect 14001 15892 14013 15895
rect 13780 15864 14013 15892
rect 13780 15852 13786 15864
rect 14001 15861 14013 15864
rect 14047 15861 14059 15895
rect 14001 15855 14059 15861
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 17129 15895 17187 15901
rect 17129 15892 17141 15895
rect 16356 15864 17141 15892
rect 16356 15852 16362 15864
rect 17129 15861 17141 15864
rect 17175 15861 17187 15895
rect 19242 15892 19248 15904
rect 19203 15864 19248 15892
rect 17129 15855 17187 15861
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2866 15688 2872 15700
rect 2827 15660 2872 15688
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4154 15688 4160 15700
rect 3927 15660 4160 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 6914 15688 6920 15700
rect 6875 15660 6920 15688
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 7098 15688 7104 15700
rect 7059 15660 7104 15688
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 8478 15688 8484 15700
rect 8439 15660 8484 15688
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9732 15660 9873 15688
rect 9732 15648 9738 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 12526 15688 12532 15700
rect 12487 15660 12532 15688
rect 9861 15651 9919 15657
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 12894 15688 12900 15700
rect 12855 15660 12900 15688
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 13265 15691 13323 15697
rect 13265 15657 13277 15691
rect 13311 15688 13323 15691
rect 14550 15688 14556 15700
rect 13311 15660 14556 15688
rect 13311 15657 13323 15660
rect 13265 15651 13323 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 15473 15691 15531 15697
rect 15473 15657 15485 15691
rect 15519 15688 15531 15691
rect 15930 15688 15936 15700
rect 15519 15660 15936 15688
rect 15519 15657 15531 15660
rect 15473 15651 15531 15657
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 16850 15648 16856 15700
rect 16908 15688 16914 15700
rect 17681 15691 17739 15697
rect 17681 15688 17693 15691
rect 16908 15660 17693 15688
rect 16908 15648 16914 15660
rect 17681 15657 17693 15660
rect 17727 15657 17739 15691
rect 21082 15688 21088 15700
rect 21043 15660 21088 15688
rect 17681 15651 17739 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 1670 15620 1676 15632
rect 1504 15592 1676 15620
rect 1504 15561 1532 15592
rect 1670 15580 1676 15592
rect 1728 15580 1734 15632
rect 1946 15580 1952 15632
rect 2004 15620 2010 15632
rect 2774 15620 2780 15632
rect 2004 15592 2780 15620
rect 2004 15580 2010 15592
rect 2774 15580 2780 15592
rect 2832 15620 2838 15632
rect 7469 15623 7527 15629
rect 7469 15620 7481 15623
rect 2832 15592 7481 15620
rect 2832 15580 2838 15592
rect 7469 15589 7481 15592
rect 7515 15620 7527 15623
rect 8846 15620 8852 15632
rect 7515 15592 8852 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 10042 15580 10048 15632
rect 10100 15620 10106 15632
rect 10658 15623 10716 15629
rect 10658 15620 10670 15623
rect 10100 15592 10670 15620
rect 10100 15580 10106 15592
rect 10658 15589 10670 15592
rect 10704 15620 10716 15623
rect 11054 15620 11060 15632
rect 10704 15592 11060 15620
rect 10704 15589 10716 15592
rect 10658 15583 10716 15589
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 17034 15620 17040 15632
rect 12032 15592 17040 15620
rect 12032 15580 12038 15592
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15521 1547 15555
rect 1489 15515 1547 15521
rect 1756 15555 1814 15561
rect 1756 15521 1768 15555
rect 1802 15552 1814 15555
rect 2498 15552 2504 15564
rect 1802 15524 2504 15552
rect 1802 15521 1814 15524
rect 1756 15515 1814 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 4884 15555 4942 15561
rect 4884 15521 4896 15555
rect 4930 15552 4942 15555
rect 5258 15552 5264 15564
rect 4930 15524 5264 15552
rect 4930 15521 4942 15524
rect 4884 15515 4942 15521
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 8205 15555 8263 15561
rect 8205 15521 8217 15555
rect 8251 15552 8263 15555
rect 8386 15552 8392 15564
rect 8251 15524 8392 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 13725 15555 13783 15561
rect 13725 15552 13737 15555
rect 13412 15524 13737 15552
rect 13412 15512 13418 15524
rect 13725 15521 13737 15524
rect 13771 15521 13783 15555
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 13725 15515 13783 15521
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16574 15561 16580 15564
rect 16568 15515 16580 15561
rect 16632 15552 16638 15564
rect 20898 15552 20904 15564
rect 16632 15524 16668 15552
rect 20859 15524 20904 15552
rect 16574 15512 16580 15515
rect 16632 15512 16638 15524
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 2866 15444 2872 15496
rect 2924 15484 2930 15496
rect 4614 15484 4620 15496
rect 2924 15456 4620 15484
rect 2924 15444 2930 15456
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 6914 15444 6920 15496
rect 6972 15484 6978 15496
rect 7098 15484 7104 15496
rect 6972 15456 7104 15484
rect 6972 15444 6978 15456
rect 7098 15444 7104 15456
rect 7156 15484 7162 15496
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7156 15456 7573 15484
rect 7156 15444 7162 15456
rect 7561 15453 7573 15456
rect 7607 15453 7619 15487
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7561 15447 7619 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 10410 15484 10416 15496
rect 10371 15456 10416 15484
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 13446 15444 13452 15496
rect 13504 15484 13510 15496
rect 13817 15487 13875 15493
rect 13817 15484 13829 15487
rect 13504 15456 13829 15484
rect 13504 15444 13510 15456
rect 13817 15453 13829 15456
rect 13863 15453 13875 15487
rect 13817 15447 13875 15453
rect 14001 15487 14059 15493
rect 14001 15453 14013 15487
rect 14047 15484 14059 15487
rect 14090 15484 14096 15496
rect 14047 15456 14096 15484
rect 14047 15453 14059 15456
rect 14001 15447 14059 15453
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 16298 15484 16304 15496
rect 16259 15456 16304 15484
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 3513 15419 3571 15425
rect 3513 15385 3525 15419
rect 3559 15416 3571 15419
rect 3602 15416 3608 15428
rect 3559 15388 3608 15416
rect 3559 15385 3571 15388
rect 3513 15379 3571 15385
rect 3602 15376 3608 15388
rect 3660 15416 3666 15428
rect 6641 15419 6699 15425
rect 3660 15388 4384 15416
rect 3660 15376 3666 15388
rect 4356 15357 4384 15388
rect 6641 15385 6653 15419
rect 6687 15416 6699 15419
rect 7760 15416 7788 15444
rect 11790 15416 11796 15428
rect 6687 15388 7788 15416
rect 11751 15388 11796 15416
rect 6687 15385 6699 15388
rect 6641 15379 6699 15385
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 12894 15416 12900 15428
rect 12400 15388 12900 15416
rect 12400 15376 12406 15388
rect 12894 15376 12900 15388
rect 12952 15376 12958 15428
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 5997 15351 6055 15357
rect 5997 15348 6009 15351
rect 4387 15320 6009 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 5997 15317 6009 15320
rect 6043 15317 6055 15351
rect 5997 15311 6055 15317
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9306 15348 9312 15360
rect 9171 15320 9312 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 9766 15348 9772 15360
rect 9539 15320 9772 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 9766 15308 9772 15320
rect 9824 15308 9830 15360
rect 10321 15351 10379 15357
rect 10321 15317 10333 15351
rect 10367 15348 10379 15351
rect 11514 15348 11520 15360
rect 10367 15320 11520 15348
rect 10367 15317 10379 15320
rect 10321 15311 10379 15317
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 13357 15351 13415 15357
rect 13357 15317 13369 15351
rect 13403 15348 13415 15351
rect 13814 15348 13820 15360
rect 13403 15320 13820 15348
rect 13403 15317 13415 15320
rect 13357 15311 13415 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14182 15308 14188 15360
rect 14240 15348 14246 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 14240 15320 14381 15348
rect 14240 15308 14246 15320
rect 14369 15317 14381 15320
rect 14415 15317 14427 15351
rect 14369 15311 14427 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 1581 15147 1639 15153
rect 1581 15144 1593 15147
rect 1452 15116 1593 15144
rect 1452 15104 1458 15116
rect 1581 15113 1593 15116
rect 1627 15113 1639 15147
rect 1581 15107 1639 15113
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1949 15147 2007 15153
rect 1949 15144 1961 15147
rect 1728 15116 1961 15144
rect 1728 15104 1734 15116
rect 1949 15113 1961 15116
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 1964 15076 1992 15107
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 2556 15116 4261 15144
rect 2556 15104 2562 15116
rect 4249 15113 4261 15116
rect 4295 15144 4307 15147
rect 4614 15144 4620 15156
rect 4295 15116 4620 15144
rect 4295 15113 4307 15116
rect 4249 15107 4307 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 6546 15104 6552 15156
rect 6604 15144 6610 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 6604 15116 8217 15144
rect 6604 15104 6610 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 11112 15116 11161 15144
rect 11112 15104 11118 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 11149 15107 11207 15113
rect 12805 15147 12863 15153
rect 12805 15113 12817 15147
rect 12851 15144 12863 15147
rect 14090 15144 14096 15156
rect 12851 15116 14096 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 2590 15076 2596 15088
rect 1964 15048 2596 15076
rect 2590 15036 2596 15048
rect 2648 15076 2654 15088
rect 2685 15079 2743 15085
rect 2685 15076 2697 15079
rect 2648 15048 2697 15076
rect 2648 15036 2654 15048
rect 2685 15045 2697 15048
rect 2731 15045 2743 15079
rect 2685 15039 2743 15045
rect 2700 15008 2728 15039
rect 4522 15036 4528 15088
rect 4580 15076 4586 15088
rect 4801 15079 4859 15085
rect 4801 15076 4813 15079
rect 4580 15048 4813 15076
rect 4580 15036 4586 15048
rect 4801 15045 4813 15048
rect 4847 15076 4859 15079
rect 6178 15076 6184 15088
rect 4847 15048 6184 15076
rect 4847 15045 4859 15048
rect 4801 15039 4859 15045
rect 6178 15036 6184 15048
rect 6236 15076 6242 15088
rect 6641 15079 6699 15085
rect 6641 15076 6653 15079
rect 6236 15048 6653 15076
rect 6236 15036 6242 15048
rect 6641 15045 6653 15048
rect 6687 15076 6699 15079
rect 19613 15079 19671 15085
rect 6687 15048 6868 15076
rect 6687 15045 6699 15048
rect 6641 15039 6699 15045
rect 2866 15008 2872 15020
rect 2700 14980 2872 15008
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 6840 15017 6868 15048
rect 19613 15045 19625 15079
rect 19659 15076 19671 15079
rect 20898 15076 20904 15088
rect 19659 15048 20904 15076
rect 19659 15045 19671 15048
rect 19613 15039 19671 15045
rect 20898 15036 20904 15048
rect 20956 15036 20962 15088
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 9122 14968 9128 15020
rect 9180 15008 9186 15020
rect 9180 14980 9812 15008
rect 9180 14968 9186 14980
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 1412 14872 1440 14903
rect 2314 14900 2320 14952
rect 2372 14940 2378 14952
rect 3136 14943 3194 14949
rect 3136 14940 3148 14943
rect 2372 14912 3148 14940
rect 2372 14900 2378 14912
rect 3136 14909 3148 14912
rect 3182 14940 3194 14943
rect 3602 14940 3608 14952
rect 3182 14912 3608 14940
rect 3182 14909 3194 14912
rect 3136 14903 3194 14909
rect 3602 14900 3608 14912
rect 3660 14900 3666 14952
rect 5350 14940 5356 14952
rect 5311 14912 5356 14940
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 6730 14940 6736 14952
rect 5920 14912 6736 14940
rect 3510 14872 3516 14884
rect 1412 14844 3516 14872
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 5074 14832 5080 14884
rect 5132 14872 5138 14884
rect 5920 14872 5948 14912
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 9784 14949 9812 14980
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16908 14980 16957 15008
rect 16908 14968 16914 14980
rect 16945 14977 16957 14980
rect 16991 15008 17003 15011
rect 17405 15011 17463 15017
rect 17405 15008 17417 15011
rect 16991 14980 17417 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 17405 14977 17417 14980
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10410 14940 10416 14952
rect 9815 14912 10416 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 5132 14844 5948 14872
rect 5132 14832 5138 14844
rect 2314 14804 2320 14816
rect 2275 14776 2320 14804
rect 2314 14764 2320 14776
rect 2372 14764 2378 14816
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 5920 14804 5948 14844
rect 6086 14832 6092 14884
rect 6144 14872 6150 14884
rect 7092 14875 7150 14881
rect 7092 14872 7104 14875
rect 6144 14844 7104 14872
rect 6144 14832 6150 14844
rect 7092 14841 7104 14844
rect 7138 14872 7150 14875
rect 7742 14872 7748 14884
rect 7138 14844 7748 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 9309 14875 9367 14881
rect 9309 14841 9321 14875
rect 9355 14872 9367 14875
rect 10014 14875 10072 14881
rect 10014 14872 10026 14875
rect 9355 14844 10026 14872
rect 9355 14841 9367 14844
rect 9309 14835 9367 14841
rect 10014 14841 10026 14844
rect 10060 14872 10072 14875
rect 10134 14872 10140 14884
rect 10060 14844 10140 14872
rect 10060 14841 10072 14844
rect 10014 14835 10072 14841
rect 10134 14832 10140 14844
rect 10192 14832 10198 14884
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5920 14776 6193 14804
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 8846 14804 8852 14816
rect 8807 14776 8852 14804
rect 6181 14767 6239 14773
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 9677 14807 9735 14813
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 10244 14804 10272 14912
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13740 14912 13921 14940
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 13354 14872 13360 14884
rect 12676 14844 13360 14872
rect 12676 14832 12682 14844
rect 13354 14832 13360 14844
rect 13412 14832 13418 14884
rect 13740 14816 13768 14912
rect 13909 14909 13921 14912
rect 13955 14940 13967 14943
rect 16209 14943 16267 14949
rect 16209 14940 16221 14943
rect 13955 14912 16221 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 16209 14909 16221 14912
rect 16255 14940 16267 14943
rect 16298 14940 16304 14952
rect 16255 14912 16304 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16298 14900 16304 14912
rect 16356 14900 16362 14952
rect 19426 14940 19432 14952
rect 19387 14912 19432 14940
rect 19426 14900 19432 14912
rect 19484 14940 19490 14952
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19484 14912 19901 14940
rect 19484 14900 19490 14912
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 19889 14903 19947 14909
rect 14182 14881 14188 14884
rect 14176 14872 14188 14881
rect 14143 14844 14188 14872
rect 14176 14835 14188 14844
rect 14182 14832 14188 14835
rect 14240 14832 14246 14884
rect 15933 14875 15991 14881
rect 15933 14841 15945 14875
rect 15979 14872 15991 14875
rect 16761 14875 16819 14881
rect 16761 14872 16773 14875
rect 15979 14844 16773 14872
rect 15979 14841 15991 14844
rect 15933 14835 15991 14841
rect 16761 14841 16773 14844
rect 16807 14872 16819 14875
rect 17494 14872 17500 14884
rect 16807 14844 17500 14872
rect 16807 14841 16819 14844
rect 16761 14835 16819 14841
rect 17494 14832 17500 14844
rect 17552 14832 17558 14884
rect 10778 14804 10784 14816
rect 9723 14776 10784 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 10778 14764 10784 14776
rect 10836 14804 10842 14816
rect 11790 14804 11796 14816
rect 10836 14776 11796 14804
rect 10836 14764 10842 14776
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13170 14804 13176 14816
rect 12943 14776 13176 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13722 14804 13728 14816
rect 13683 14776 13728 14804
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 15286 14804 15292 14816
rect 15247 14776 15292 14804
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 16390 14804 16396 14816
rect 16351 14776 16396 14804
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16850 14804 16856 14816
rect 16763 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14804 16914 14816
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 16908 14776 17785 14804
rect 16908 14764 16914 14776
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 17773 14767 17831 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2130 14560 2136 14612
rect 2188 14600 2194 14612
rect 2409 14603 2467 14609
rect 2409 14600 2421 14603
rect 2188 14572 2421 14600
rect 2188 14560 2194 14572
rect 2409 14569 2421 14572
rect 2455 14569 2467 14603
rect 2409 14563 2467 14569
rect 2498 14560 2504 14612
rect 2556 14600 2562 14612
rect 3510 14600 3516 14612
rect 2556 14572 3004 14600
rect 3471 14572 3516 14600
rect 2556 14560 2562 14572
rect 1397 14535 1455 14541
rect 1397 14501 1409 14535
rect 1443 14532 1455 14535
rect 2866 14532 2872 14544
rect 1443 14504 2872 14532
rect 1443 14501 1455 14504
rect 1397 14495 1455 14501
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 2832 14436 2877 14464
rect 2832 14424 2838 14436
rect 2976 14405 3004 14572
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4062 14600 4068 14612
rect 4023 14572 4068 14600
rect 4062 14560 4068 14572
rect 4120 14560 4126 14612
rect 4522 14600 4528 14612
rect 4483 14572 4528 14600
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 5997 14603 6055 14609
rect 5997 14569 6009 14603
rect 6043 14600 6055 14603
rect 6086 14600 6092 14612
rect 6043 14572 6092 14600
rect 6043 14569 6055 14572
rect 5997 14563 6055 14569
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 7466 14600 7472 14612
rect 7427 14572 7472 14600
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 8386 14600 8392 14612
rect 8347 14572 8392 14600
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 9030 14600 9036 14612
rect 8991 14572 9036 14600
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 10778 14600 10784 14612
rect 10739 14572 10784 14600
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11609 14603 11667 14609
rect 11609 14569 11621 14603
rect 11655 14600 11667 14603
rect 12342 14600 12348 14612
rect 11655 14572 12348 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 13630 14600 13636 14612
rect 13591 14572 13636 14600
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13872 14572 14105 14600
rect 13872 14560 13878 14572
rect 14093 14569 14105 14572
rect 14139 14600 14151 14603
rect 14458 14600 14464 14612
rect 14139 14572 14464 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 15378 14560 15384 14612
rect 15436 14600 15442 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 15436 14572 15485 14600
rect 15436 14560 15442 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 15473 14563 15531 14569
rect 15933 14603 15991 14609
rect 15933 14569 15945 14603
rect 15979 14600 15991 14603
rect 16850 14600 16856 14612
rect 15979 14572 16856 14600
rect 15979 14569 15991 14572
rect 15933 14563 15991 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17494 14600 17500 14612
rect 17455 14572 17500 14600
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 6356 14535 6414 14541
rect 6356 14501 6368 14535
rect 6402 14532 6414 14535
rect 6546 14532 6552 14544
rect 6402 14504 6552 14532
rect 6402 14501 6414 14504
rect 6356 14495 6414 14501
rect 6546 14492 6552 14504
rect 6604 14492 6610 14544
rect 11698 14492 11704 14544
rect 11756 14532 11762 14544
rect 12069 14535 12127 14541
rect 12069 14532 12081 14535
rect 11756 14504 12081 14532
rect 11756 14492 11762 14504
rect 12069 14501 12081 14504
rect 12115 14501 12127 14535
rect 12069 14495 12127 14501
rect 14734 14492 14740 14544
rect 14792 14532 14798 14544
rect 16390 14532 16396 14544
rect 14792 14504 16396 14532
rect 14792 14492 14798 14504
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 3878 14464 3884 14476
rect 3839 14436 3884 14464
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4212 14436 4445 14464
rect 4212 14424 4218 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 6089 14467 6147 14473
rect 6089 14433 6101 14467
rect 6135 14464 6147 14467
rect 6178 14464 6184 14476
rect 6135 14436 6184 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 6178 14424 6184 14436
rect 6236 14424 6242 14476
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 11146 14464 11152 14476
rect 10183 14436 11152 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11480 14436 11989 14464
rect 11480 14424 11486 14436
rect 11977 14433 11989 14436
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 13228 14436 14013 14464
rect 13228 14424 13234 14436
rect 14001 14433 14013 14436
rect 14047 14433 14059 14467
rect 14001 14427 14059 14433
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 15988 14436 16313 14464
rect 15988 14424 15994 14436
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 2884 14328 2912 14359
rect 3786 14356 3792 14408
rect 3844 14356 3850 14408
rect 4614 14396 4620 14408
rect 4575 14368 4620 14396
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 8018 14396 8024 14408
rect 7979 14368 8024 14396
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8570 14396 8576 14408
rect 8531 14368 8576 14396
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10686 14396 10692 14408
rect 10367 14368 10692 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 3142 14328 3148 14340
rect 2884 14300 3148 14328
rect 3142 14288 3148 14300
rect 3200 14328 3206 14340
rect 3804 14328 3832 14356
rect 3200 14300 3832 14328
rect 3200 14288 3206 14300
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 5350 14328 5356 14340
rect 5132 14300 5356 14328
rect 5132 14288 5138 14300
rect 5350 14288 5356 14300
rect 5408 14328 5414 14340
rect 5537 14331 5595 14337
rect 5537 14328 5549 14331
rect 5408 14300 5549 14328
rect 5408 14288 5414 14300
rect 5537 14297 5549 14300
rect 5583 14297 5595 14331
rect 5537 14291 5595 14297
rect 9398 14288 9404 14340
rect 9456 14328 9462 14340
rect 9493 14331 9551 14337
rect 9493 14328 9505 14331
rect 9456 14300 9505 14328
rect 9456 14288 9462 14300
rect 9493 14297 9505 14300
rect 9539 14328 9551 14331
rect 10336 14328 10364 14359
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 12250 14396 12256 14408
rect 12211 14368 12256 14396
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 13354 14396 13360 14408
rect 13315 14368 13360 14396
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 14182 14356 14188 14408
rect 14240 14396 14246 14408
rect 16574 14396 16580 14408
rect 14240 14368 14285 14396
rect 16535 14368 16580 14396
rect 14240 14356 14246 14368
rect 16574 14356 16580 14368
rect 16632 14396 16638 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16632 14368 16957 14396
rect 16632 14356 16638 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 9539 14300 10364 14328
rect 9539 14297 9551 14300
rect 9493 14291 9551 14297
rect 2222 14260 2228 14272
rect 2183 14232 2228 14260
rect 2222 14220 2228 14232
rect 2280 14260 2286 14272
rect 2498 14260 2504 14272
rect 2280 14232 2504 14260
rect 2280 14220 2286 14232
rect 2498 14220 2504 14232
rect 2556 14220 2562 14272
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 3970 14260 3976 14272
rect 3476 14232 3976 14260
rect 3476 14220 3482 14232
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 5258 14260 5264 14272
rect 5219 14232 5264 14260
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 9674 14260 9680 14272
rect 9635 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2593 14059 2651 14065
rect 2593 14056 2605 14059
rect 2372 14028 2605 14056
rect 2372 14016 2378 14028
rect 2593 14025 2605 14028
rect 2639 14025 2651 14059
rect 2593 14019 2651 14025
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3145 14059 3203 14065
rect 3145 14056 3157 14059
rect 2832 14028 3157 14056
rect 2832 14016 2838 14028
rect 3145 14025 3157 14028
rect 3191 14056 3203 14059
rect 3326 14056 3332 14068
rect 3191 14028 3332 14056
rect 3191 14025 3203 14028
rect 3145 14019 3203 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 7190 14056 7196 14068
rect 7147 14028 7196 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9122 14056 9128 14068
rect 9079 14028 9128 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 10192 14028 10517 14056
rect 10192 14016 10198 14028
rect 10505 14025 10517 14028
rect 10551 14025 10563 14059
rect 10505 14019 10563 14025
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11756 14028 11989 14056
rect 11756 14016 11762 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 13170 14056 13176 14068
rect 13131 14028 13176 14056
rect 11977 14019 12035 14025
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 16390 14056 16396 14068
rect 16351 14028 16396 14056
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16632 14028 16681 14056
rect 16632 14016 16638 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 3602 13948 3608 14000
rect 3660 13988 3666 14000
rect 7561 13991 7619 13997
rect 3660 13960 3740 13988
rect 3660 13948 3666 13960
rect 1854 13880 1860 13932
rect 1912 13920 1918 13932
rect 2041 13923 2099 13929
rect 2041 13920 2053 13923
rect 1912 13892 2053 13920
rect 1912 13880 1918 13892
rect 2041 13889 2053 13892
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13920 2283 13923
rect 2314 13920 2320 13932
rect 2271 13892 2320 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 3712 13929 3740 13960
rect 7561 13957 7573 13991
rect 7607 13988 7619 13991
rect 8202 13988 8208 14000
rect 7607 13960 8208 13988
rect 7607 13957 7619 13960
rect 7561 13951 7619 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5123 13892 5733 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5721 13889 5733 13892
rect 5767 13920 5779 13923
rect 6914 13920 6920 13932
rect 5767 13892 6920 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 8110 13920 8116 13932
rect 8023 13892 8116 13920
rect 8110 13880 8116 13892
rect 8168 13920 8174 13932
rect 8665 13923 8723 13929
rect 8665 13920 8677 13923
rect 8168 13892 8677 13920
rect 8168 13880 8174 13892
rect 8665 13889 8677 13892
rect 8711 13920 8723 13923
rect 11146 13920 11152 13932
rect 8711 13892 9260 13920
rect 11107 13892 11152 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 3050 13852 3056 13864
rect 2963 13824 3056 13852
rect 3050 13812 3056 13824
rect 3108 13852 3114 13864
rect 3602 13852 3608 13864
rect 3108 13824 3608 13852
rect 3108 13812 3114 13824
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 6840 13824 7389 13852
rect 3510 13784 3516 13796
rect 3471 13756 3516 13784
rect 3510 13744 3516 13756
rect 3568 13744 3574 13796
rect 5258 13744 5264 13796
rect 5316 13784 5322 13796
rect 5629 13787 5687 13793
rect 5629 13784 5641 13787
rect 5316 13756 5641 13784
rect 5316 13744 5322 13756
rect 5629 13753 5641 13756
rect 5675 13753 5687 13787
rect 5629 13747 5687 13753
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 6840 13784 6868 13824
rect 7377 13821 7389 13824
rect 7423 13852 7435 13855
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 7423 13824 8033 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 9122 13852 9128 13864
rect 9083 13824 9128 13852
rect 8021 13815 8079 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 9232 13852 9260 13892
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 9398 13861 9404 13864
rect 9392 13852 9404 13861
rect 9232 13824 9404 13852
rect 9392 13815 9404 13824
rect 9398 13812 9404 13815
rect 9456 13812 9462 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11609 13855 11667 13861
rect 11609 13852 11621 13855
rect 11480 13824 11621 13852
rect 11480 13812 11486 13824
rect 11609 13821 11621 13824
rect 11655 13821 11667 13855
rect 13722 13852 13728 13864
rect 11609 13815 11667 13821
rect 13556 13824 13728 13852
rect 6788 13756 6868 13784
rect 6788 13744 6794 13756
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7929 13787 7987 13793
rect 7929 13784 7941 13787
rect 7248 13756 7941 13784
rect 7248 13744 7254 13756
rect 7392 13728 7420 13756
rect 7929 13753 7941 13756
rect 7975 13753 7987 13787
rect 7929 13747 7987 13753
rect 12437 13787 12495 13793
rect 12437 13753 12449 13787
rect 12483 13784 12495 13787
rect 12802 13784 12808 13796
rect 12483 13756 12808 13784
rect 12483 13753 12495 13756
rect 12437 13747 12495 13753
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 1581 13719 1639 13725
rect 1581 13685 1593 13719
rect 1627 13716 1639 13719
rect 2406 13716 2412 13728
rect 1627 13688 2412 13716
rect 1627 13685 1639 13688
rect 1581 13679 1639 13685
rect 2406 13676 2412 13688
rect 2464 13676 2470 13728
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 6546 13716 6552 13728
rect 6507 13688 6552 13716
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 7374 13676 7380 13728
rect 7432 13676 7438 13728
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13556 13725 13584 13824
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 15930 13852 15936 13864
rect 15891 13824 15936 13852
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 13992 13787 14050 13793
rect 13992 13753 14004 13787
rect 14038 13784 14050 13787
rect 14090 13784 14096 13796
rect 14038 13756 14096 13784
rect 14038 13753 14050 13756
rect 13992 13747 14050 13753
rect 14090 13744 14096 13756
rect 14148 13744 14154 13796
rect 13541 13719 13599 13725
rect 13541 13716 13553 13719
rect 13228 13688 13553 13716
rect 13228 13676 13234 13688
rect 13541 13685 13553 13688
rect 13587 13685 13599 13719
rect 13541 13679 13599 13685
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 15105 13719 15163 13725
rect 15105 13716 15117 13719
rect 14240 13688 15117 13716
rect 14240 13676 14246 13688
rect 15105 13685 15117 13688
rect 15151 13685 15163 13719
rect 15105 13679 15163 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 3237 13515 3295 13521
rect 3237 13481 3249 13515
rect 3283 13512 3295 13515
rect 3510 13512 3516 13524
rect 3283 13484 3516 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4430 13512 4436 13524
rect 4391 13484 4436 13512
rect 4430 13472 4436 13484
rect 4488 13512 4494 13524
rect 4890 13512 4896 13524
rect 4488 13484 4896 13512
rect 4488 13472 4494 13484
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 6914 13512 6920 13524
rect 6875 13484 6920 13512
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8110 13512 8116 13524
rect 8071 13484 8116 13512
rect 8110 13472 8116 13484
rect 8168 13472 8174 13524
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9674 13512 9680 13524
rect 9171 13484 9680 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9674 13472 9680 13484
rect 9732 13512 9738 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 9732 13484 10057 13512
rect 9732 13472 9738 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 12584 13484 13185 13512
rect 12584 13472 12590 13484
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 13173 13475 13231 13481
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 14182 13512 14188 13524
rect 13863 13484 14188 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 14182 13472 14188 13484
rect 14240 13472 14246 13524
rect 14458 13512 14464 13524
rect 14419 13484 14464 13512
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16632 13484 16957 13512
rect 16632 13472 16638 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 16945 13475 17003 13481
rect 21085 13515 21143 13521
rect 21085 13481 21097 13515
rect 21131 13512 21143 13515
rect 21174 13512 21180 13524
rect 21131 13484 21180 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 1673 13447 1731 13453
rect 1673 13413 1685 13447
rect 1719 13444 1731 13447
rect 1854 13444 1860 13456
rect 1719 13416 1860 13444
rect 1719 13413 1731 13416
rect 1673 13407 1731 13413
rect 1854 13404 1860 13416
rect 1912 13404 1918 13456
rect 2041 13447 2099 13453
rect 2041 13413 2053 13447
rect 2087 13444 2099 13447
rect 2222 13444 2228 13456
rect 2087 13416 2228 13444
rect 2087 13413 2099 13416
rect 2041 13407 2099 13413
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 2406 13404 2412 13456
rect 2464 13444 2470 13456
rect 2593 13447 2651 13453
rect 2593 13444 2605 13447
rect 2464 13416 2605 13444
rect 2464 13404 2470 13416
rect 2593 13413 2605 13416
rect 2639 13444 2651 13447
rect 3142 13444 3148 13456
rect 2639 13416 3148 13444
rect 2639 13413 2651 13416
rect 2593 13407 2651 13413
rect 3142 13404 3148 13416
rect 3200 13404 3206 13456
rect 4525 13447 4583 13453
rect 4525 13413 4537 13447
rect 4571 13444 4583 13447
rect 4798 13444 4804 13456
rect 4571 13416 4804 13444
rect 4571 13413 4583 13416
rect 4525 13407 4583 13413
rect 4798 13404 4804 13416
rect 4856 13404 4862 13456
rect 5813 13447 5871 13453
rect 5813 13413 5825 13447
rect 5859 13444 5871 13447
rect 6270 13444 6276 13456
rect 5859 13416 6276 13444
rect 5859 13413 5871 13416
rect 5813 13407 5871 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 9398 13444 9404 13456
rect 9359 13416 9404 13444
rect 9398 13404 9404 13416
rect 9456 13404 9462 13456
rect 11238 13404 11244 13456
rect 11296 13444 11302 13456
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 11296 13416 11713 13444
rect 11296 13404 11302 13416
rect 11701 13413 11713 13416
rect 11747 13444 11759 13447
rect 12060 13447 12118 13453
rect 12060 13444 12072 13447
rect 11747 13416 12072 13444
rect 11747 13413 11759 13416
rect 11701 13407 11759 13413
rect 12060 13413 12072 13416
rect 12106 13444 12118 13447
rect 12250 13444 12256 13456
rect 12106 13416 12256 13444
rect 12106 13413 12118 13416
rect 12060 13407 12118 13413
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 4062 13376 4068 13388
rect 2547 13348 4068 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 6546 13376 6552 13388
rect 5491 13348 6552 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 4614 13308 4620 13320
rect 4575 13280 4620 13308
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 6472 13317 6500 13348
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 7466 13376 7472 13388
rect 7427 13348 7472 13376
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 15838 13385 15844 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 8352 13348 10149 13376
rect 8352 13336 8358 13348
rect 10137 13345 10149 13348
rect 10183 13345 10195 13379
rect 15832 13376 15844 13385
rect 15799 13348 15844 13376
rect 10137 13339 10195 13345
rect 15832 13339 15844 13348
rect 15838 13336 15844 13339
rect 15896 13336 15902 13388
rect 18316 13379 18374 13385
rect 18316 13345 18328 13379
rect 18362 13376 18374 13379
rect 19150 13376 19156 13388
rect 18362 13348 19156 13376
rect 18362 13345 18374 13348
rect 18316 13339 18374 13345
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 20898 13376 20904 13388
rect 20859 13348 20904 13376
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 9122 13308 9128 13320
rect 8619 13280 9128 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 10226 13308 10232 13320
rect 10187 13280 10232 13308
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15528 13280 15577 13308
rect 15528 13268 15534 13280
rect 15565 13277 15577 13280
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 17828 13280 18061 13308
rect 17828 13268 17834 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 5258 13240 5264 13252
rect 3927 13212 5264 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 5905 13243 5963 13249
rect 5905 13209 5917 13243
rect 5951 13240 5963 13243
rect 5994 13240 6000 13252
rect 5951 13212 6000 13240
rect 5951 13209 5963 13212
rect 5905 13203 5963 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 7650 13240 7656 13252
rect 7611 13212 7656 13240
rect 7650 13200 7656 13212
rect 7708 13200 7714 13252
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 9766 13240 9772 13252
rect 9723 13212 9772 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 19426 13240 19432 13252
rect 19387 13212 19432 13240
rect 19426 13200 19432 13212
rect 19484 13200 19490 13252
rect 2133 13175 2191 13181
rect 2133 13141 2145 13175
rect 2179 13172 2191 13175
rect 2222 13172 2228 13184
rect 2179 13144 2228 13172
rect 2179 13141 2191 13144
rect 2133 13135 2191 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 4062 13172 4068 13184
rect 4023 13144 4068 13172
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 5592 13144 7297 13172
rect 5592 13132 5598 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 7285 13135 7343 13141
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14884 13144 14933 13172
rect 14884 13132 14890 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 14921 13135 14979 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 2590 12968 2596 12980
rect 2547 12940 2596 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 3936 12940 3985 12968
rect 3936 12928 3942 12940
rect 3973 12937 3985 12940
rect 4019 12968 4031 12971
rect 4614 12968 4620 12980
rect 4019 12940 4620 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5258 12968 5264 12980
rect 5215 12940 5264 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6273 12971 6331 12977
rect 6273 12968 6285 12971
rect 6236 12940 6285 12968
rect 6236 12928 6242 12940
rect 6273 12937 6285 12940
rect 6319 12968 6331 12971
rect 6362 12968 6368 12980
rect 6319 12940 6368 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 8294 12928 8300 12980
rect 8352 12968 8358 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8352 12940 8769 12968
rect 8352 12928 8358 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 9122 12968 9128 12980
rect 9083 12940 9128 12968
rect 8757 12931 8815 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9306 12968 9312 12980
rect 9267 12940 9312 12968
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 10284 12940 10333 12968
rect 10284 12928 10290 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 11238 12968 11244 12980
rect 11199 12940 11244 12968
rect 10321 12931 10379 12937
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 12710 12968 12716 12980
rect 11624 12940 12716 12968
rect 1946 12792 1952 12844
rect 2004 12832 2010 12844
rect 2608 12841 2636 12928
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 9640 12872 9996 12900
rect 9640 12860 9646 12872
rect 2593 12835 2651 12841
rect 2593 12832 2605 12835
rect 2004 12804 2605 12832
rect 2004 12792 2010 12804
rect 2593 12801 2605 12804
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4798 12832 4804 12844
rect 4663 12804 4804 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 5350 12792 5356 12844
rect 5408 12832 5414 12844
rect 5810 12832 5816 12844
rect 5408 12804 5816 12832
rect 5408 12792 5414 12804
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6328 12804 6561 12832
rect 6328 12792 6334 12804
rect 6549 12801 6561 12804
rect 6595 12832 6607 12835
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6595 12804 6837 12832
rect 6595 12801 6607 12804
rect 6549 12795 6607 12801
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 9766 12832 9772 12844
rect 8536 12804 9772 12832
rect 8536 12792 8542 12804
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 9968 12841 9996 12872
rect 9953 12835 10011 12841
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10244 12832 10272 12928
rect 10873 12903 10931 12909
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 11330 12900 11336 12912
rect 10919 12872 11336 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 11330 12860 11336 12872
rect 11388 12900 11394 12912
rect 11624 12900 11652 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 16264 12940 16405 12968
rect 16264 12928 16270 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 16393 12931 16451 12937
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 22278 12928 22284 12980
rect 22336 12968 22342 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 22336 12940 22477 12968
rect 22336 12928 22342 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 22465 12931 22523 12937
rect 13814 12900 13820 12912
rect 11388 12872 11652 12900
rect 13775 12872 13820 12900
rect 11388 12860 11394 12872
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 15102 12900 15108 12912
rect 15063 12872 15108 12900
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 9999 12804 10272 12832
rect 17037 12835 17095 12841
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17313 12835 17371 12841
rect 17313 12832 17325 12835
rect 17083 12804 17325 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17313 12801 17325 12804
rect 17359 12801 17371 12835
rect 17313 12795 17371 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2498 12764 2504 12776
rect 1443 12736 2504 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2498 12724 2504 12736
rect 2556 12724 2562 12776
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12764 5595 12767
rect 5626 12764 5632 12776
rect 5583 12736 5632 12764
rect 5583 12733 5595 12736
rect 5537 12727 5595 12733
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 2133 12699 2191 12705
rect 2133 12665 2145 12699
rect 2179 12696 2191 12699
rect 2838 12699 2896 12705
rect 2838 12696 2850 12699
rect 2179 12668 2850 12696
rect 2179 12665 2191 12668
rect 2133 12659 2191 12665
rect 2838 12665 2850 12668
rect 2884 12696 2896 12699
rect 2958 12696 2964 12708
rect 2884 12668 2964 12696
rect 2884 12665 2896 12668
rect 2838 12659 2896 12665
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 5442 12656 5448 12708
rect 5500 12696 5506 12708
rect 6288 12696 6316 12792
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7081 12767 7139 12773
rect 7081 12764 7093 12767
rect 6972 12736 7093 12764
rect 6972 12724 6978 12736
rect 7081 12733 7093 12736
rect 7127 12733 7139 12767
rect 7081 12727 7139 12733
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 11330 12773 11336 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 9180 12736 9689 12764
rect 9180 12724 9186 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 11325 12727 11336 12773
rect 11388 12764 11394 12776
rect 12437 12767 12495 12773
rect 11388 12736 11425 12764
rect 11330 12724 11336 12727
rect 11388 12724 11394 12736
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 5500 12668 6316 12696
rect 5500 12656 5506 12668
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12628 5046 12640
rect 5629 12631 5687 12637
rect 5629 12628 5641 12631
rect 5040 12600 5641 12628
rect 5040 12588 5046 12600
rect 5629 12597 5641 12600
rect 5675 12628 5687 12631
rect 6730 12628 6736 12640
rect 5675 12600 6736 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 8202 12628 8208 12640
rect 8163 12600 8208 12628
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 11885 12631 11943 12637
rect 11885 12628 11897 12631
rect 11848 12600 11897 12628
rect 11848 12588 11854 12600
rect 11885 12597 11897 12600
rect 11931 12628 11943 12631
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11931 12600 12265 12628
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 12253 12597 12265 12600
rect 12299 12628 12311 12631
rect 12452 12628 12480 12727
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14826 12764 14832 12776
rect 13872 12736 14832 12764
rect 13872 12724 13878 12736
rect 14826 12724 14832 12736
rect 14884 12764 14890 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14884 12736 14933 12764
rect 14884 12724 14890 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16347 12736 16773 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16761 12733 16773 12736
rect 16807 12764 16819 12767
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 16807 12736 18061 12764
rect 16807 12733 16819 12736
rect 16761 12727 16819 12733
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 22278 12764 22284 12776
rect 22239 12736 22284 12764
rect 18049 12727 18107 12733
rect 22278 12724 22284 12736
rect 22336 12764 22342 12776
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22336 12736 22753 12764
rect 22336 12724 22342 12736
rect 22741 12733 22753 12736
rect 22787 12733 22799 12767
rect 22741 12727 22799 12733
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12710 12705 12716 12708
rect 12682 12699 12716 12705
rect 12682 12696 12694 12699
rect 12584 12668 12694 12696
rect 12584 12656 12590 12668
rect 12682 12665 12694 12668
rect 12768 12696 12774 12708
rect 15194 12696 15200 12708
rect 12768 12668 12830 12696
rect 14568 12668 15200 12696
rect 12682 12659 12716 12665
rect 12710 12656 12716 12659
rect 12768 12656 12774 12668
rect 13170 12628 13176 12640
rect 12299 12600 13176 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 13170 12588 13176 12600
rect 13228 12628 13234 12640
rect 14568 12628 14596 12668
rect 15194 12656 15200 12668
rect 15252 12696 15258 12708
rect 15470 12696 15476 12708
rect 15252 12668 15476 12696
rect 15252 12656 15258 12668
rect 15470 12656 15476 12668
rect 15528 12696 15534 12708
rect 15565 12699 15623 12705
rect 15565 12696 15577 12699
rect 15528 12668 15577 12696
rect 15528 12656 15534 12668
rect 15565 12665 15577 12668
rect 15611 12665 15623 12699
rect 15565 12659 15623 12665
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 17828 12668 18521 12696
rect 17828 12656 17834 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 14826 12628 14832 12640
rect 13228 12600 14596 12628
rect 14787 12600 14832 12628
rect 13228 12588 13234 12600
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 16853 12631 16911 12637
rect 16853 12597 16865 12631
rect 16899 12628 16911 12631
rect 17218 12628 17224 12640
rect 16899 12600 17224 12628
rect 16899 12597 16911 12600
rect 16853 12591 16911 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12628 17371 12631
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17359 12600 17509 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17497 12597 17509 12600
rect 17543 12628 17555 12631
rect 18969 12631 19027 12637
rect 18969 12628 18981 12631
rect 17543 12600 18981 12628
rect 17543 12597 17555 12600
rect 17497 12591 17555 12597
rect 18969 12597 18981 12600
rect 19015 12628 19027 12631
rect 19150 12628 19156 12640
rect 19015 12600 19156 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 2314 12424 2320 12436
rect 1719 12396 2320 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 2314 12384 2320 12396
rect 2372 12424 2378 12436
rect 3878 12424 3884 12436
rect 2372 12396 3884 12424
rect 2372 12384 2378 12396
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4246 12424 4252 12436
rect 4207 12396 4252 12424
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4709 12427 4767 12433
rect 4709 12393 4721 12427
rect 4755 12424 4767 12427
rect 4890 12424 4896 12436
rect 4755 12396 4896 12424
rect 4755 12393 4767 12396
rect 4709 12387 4767 12393
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 6822 12424 6828 12436
rect 6783 12396 6828 12424
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9582 12424 9588 12436
rect 9447 12396 9588 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9766 12424 9772 12436
rect 9723 12396 9772 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11238 12424 11244 12436
rect 11199 12396 11244 12424
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11609 12427 11667 12433
rect 11609 12393 11621 12427
rect 11655 12424 11667 12427
rect 11698 12424 11704 12436
rect 11655 12396 11704 12424
rect 11655 12393 11667 12396
rect 11609 12387 11667 12393
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12710 12424 12716 12436
rect 12575 12396 12716 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 19150 12424 19156 12436
rect 19111 12396 19156 12424
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 22002 12424 22008 12436
rect 21963 12396 22008 12424
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 2832 12328 2877 12356
rect 2832 12316 2838 12328
rect 15286 12316 15292 12368
rect 15344 12356 15350 12368
rect 15534 12359 15592 12365
rect 15534 12356 15546 12359
rect 15344 12328 15546 12356
rect 15344 12316 15350 12328
rect 15534 12325 15546 12328
rect 15580 12325 15592 12359
rect 15534 12319 15592 12325
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12257 2191 12291
rect 2133 12251 2191 12257
rect 1762 12152 1768 12164
rect 1723 12124 1768 12152
rect 1762 12112 1768 12124
rect 1820 12112 1826 12164
rect 2148 12152 2176 12251
rect 2222 12248 2228 12300
rect 2280 12288 2286 12300
rect 2682 12288 2688 12300
rect 2280 12260 2688 12288
rect 2280 12248 2286 12260
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 5712 12291 5770 12297
rect 5712 12288 5724 12291
rect 5408 12260 5724 12288
rect 5408 12248 5414 12260
rect 5712 12257 5724 12260
rect 5758 12288 5770 12291
rect 5994 12288 6000 12300
rect 5758 12260 6000 12288
rect 5758 12257 5770 12260
rect 5712 12251 5770 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 8294 12288 8300 12300
rect 8255 12260 8300 12288
rect 8294 12248 8300 12260
rect 8352 12248 8358 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 10137 12291 10195 12297
rect 10137 12257 10149 12291
rect 10183 12288 10195 12291
rect 10778 12288 10784 12300
rect 10183 12260 10784 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 11701 12291 11759 12297
rect 11701 12288 11713 12291
rect 11572 12260 11713 12288
rect 11572 12248 11578 12260
rect 11701 12257 11713 12260
rect 11747 12257 11759 12291
rect 13998 12288 14004 12300
rect 13959 12260 14004 12288
rect 11701 12251 11759 12257
rect 13998 12248 14004 12260
rect 14056 12248 14062 12300
rect 17770 12288 17776 12300
rect 15304 12260 17776 12288
rect 2314 12220 2320 12232
rect 2275 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 5442 12220 5448 12232
rect 5403 12192 5448 12220
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 8386 12220 8392 12232
rect 8347 12192 8392 12220
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8662 12220 8668 12232
rect 8619 12192 8668 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8662 12180 8668 12192
rect 8720 12220 8726 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8720 12192 8953 12220
rect 8720 12180 8726 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 8941 12183 8999 12189
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10686 12220 10692 12232
rect 10367 12192 10692 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10686 12180 10692 12192
rect 10744 12220 10750 12232
rect 10962 12220 10968 12232
rect 10744 12192 10968 12220
rect 10744 12180 10750 12192
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 11790 12220 11796 12232
rect 11751 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12180 11854 12232
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 14458 12220 14464 12232
rect 14323 12192 14464 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 2222 12152 2228 12164
rect 2148 12124 2228 12152
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 2648 12056 3157 12084
rect 2648 12044 2654 12056
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3145 12047 3203 12053
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5169 12087 5227 12093
rect 5169 12084 5181 12087
rect 4764 12056 5181 12084
rect 4764 12044 4770 12056
rect 5169 12053 5181 12056
rect 5215 12084 5227 12087
rect 5258 12084 5264 12096
rect 5215 12056 5264 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 7466 12084 7472 12096
rect 7427 12056 7472 12084
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 7926 12084 7932 12096
rect 7887 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 13078 12084 13084 12096
rect 13039 12056 13084 12084
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13446 12084 13452 12096
rect 13407 12056 13452 12084
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 13630 12084 13636 12096
rect 13591 12056 13636 12084
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 14108 12084 14136 12183
rect 14458 12180 14464 12192
rect 14516 12220 14522 12232
rect 14826 12220 14832 12232
rect 14516 12192 14832 12220
rect 14516 12180 14522 12192
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15304 12229 15332 12260
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 18046 12297 18052 12300
rect 18040 12288 18052 12297
rect 18007 12260 18052 12288
rect 18040 12251 18052 12260
rect 18046 12248 18052 12251
rect 18104 12248 18110 12300
rect 21821 12291 21879 12297
rect 21821 12257 21833 12291
rect 21867 12288 21879 12291
rect 21867 12260 22048 12288
rect 21867 12257 21879 12260
rect 21821 12251 21879 12257
rect 22020 12232 22048 12260
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 15252 12192 15301 12220
rect 15252 12180 15258 12192
rect 15289 12189 15301 12192
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 22002 12180 22008 12232
rect 22060 12180 22066 12232
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 16669 12155 16727 12161
rect 16669 12152 16681 12155
rect 16632 12124 16681 12152
rect 16632 12112 16638 12124
rect 16669 12121 16681 12124
rect 16715 12121 16727 12155
rect 16669 12115 16727 12121
rect 14734 12084 14740 12096
rect 14108 12056 14740 12084
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 17218 12084 17224 12096
rect 17179 12056 17224 12084
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1673 11883 1731 11889
rect 1673 11849 1685 11883
rect 1719 11880 1731 11883
rect 2314 11880 2320 11892
rect 1719 11852 2320 11880
rect 1719 11849 1731 11852
rect 1673 11843 1731 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 3510 11880 3516 11892
rect 2832 11852 3516 11880
rect 2832 11840 2838 11852
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 5169 11883 5227 11889
rect 5169 11849 5181 11883
rect 5215 11880 5227 11883
rect 5534 11880 5540 11892
rect 5215 11852 5540 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8294 11880 8300 11892
rect 7975 11852 8300 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 1946 11812 1952 11824
rect 1907 11784 1952 11812
rect 1946 11772 1952 11784
rect 2004 11812 2010 11824
rect 2004 11784 2176 11812
rect 2004 11772 2010 11784
rect 2148 11753 2176 11784
rect 2133 11747 2191 11753
rect 2133 11713 2145 11747
rect 2179 11713 2191 11747
rect 2133 11707 2191 11713
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 4755 11716 5825 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 5813 11713 5825 11716
rect 5859 11744 5871 11747
rect 5994 11744 6000 11756
rect 5859 11716 6000 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 5994 11704 6000 11716
rect 6052 11744 6058 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6052 11716 6561 11744
rect 6052 11704 6058 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6549 11707 6607 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 7944 11744 7972 11843
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 10778 11880 10784 11892
rect 10739 11852 10784 11880
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11238 11880 11244 11892
rect 11151 11852 11244 11880
rect 11238 11840 11244 11852
rect 11296 11880 11302 11892
rect 11790 11880 11796 11892
rect 11296 11852 11796 11880
rect 11296 11840 11302 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 15289 11883 15347 11889
rect 15289 11849 15301 11883
rect 15335 11880 15347 11883
rect 15470 11880 15476 11892
rect 15335 11852 15476 11880
rect 15335 11849 15347 11852
rect 15289 11843 15347 11849
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 16025 11883 16083 11889
rect 16025 11849 16037 11883
rect 16071 11880 16083 11883
rect 17218 11880 17224 11892
rect 16071 11852 17224 11880
rect 16071 11849 16083 11852
rect 16025 11843 16083 11849
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 21361 11883 21419 11889
rect 21361 11849 21373 11883
rect 21407 11880 21419 11883
rect 22186 11880 22192 11892
rect 21407 11852 22192 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 7423 11716 7972 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16448 11716 16497 11744
rect 16448 11704 16454 11716
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11744 16727 11747
rect 17126 11744 17132 11756
rect 16715 11716 17132 11744
rect 16715 11713 16727 11716
rect 16669 11707 16727 11713
rect 17126 11704 17132 11716
rect 17184 11744 17190 11756
rect 18046 11744 18052 11756
rect 17184 11716 18052 11744
rect 17184 11704 17190 11716
rect 18046 11704 18052 11716
rect 18104 11744 18110 11756
rect 18509 11747 18567 11753
rect 18509 11744 18521 11747
rect 18104 11716 18521 11744
rect 18104 11704 18110 11716
rect 18509 11713 18521 11716
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 2406 11685 2412 11688
rect 2400 11676 2412 11685
rect 2367 11648 2412 11676
rect 2400 11639 2412 11648
rect 2406 11636 2412 11639
rect 2464 11636 2470 11688
rect 8662 11685 8668 11688
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8159 11648 8401 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8656 11676 8668 11685
rect 8389 11639 8447 11645
rect 8496 11648 8668 11676
rect 2498 11568 2504 11620
rect 2556 11608 2562 11620
rect 4062 11608 4068 11620
rect 2556 11580 4068 11608
rect 2556 11568 2562 11580
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 4154 11568 4160 11620
rect 4212 11608 4218 11620
rect 4985 11611 5043 11617
rect 4985 11608 4997 11611
rect 4212 11580 4997 11608
rect 4212 11568 4218 11580
rect 4985 11577 4997 11580
rect 5031 11608 5043 11611
rect 5629 11611 5687 11617
rect 5629 11608 5641 11611
rect 5031 11580 5641 11608
rect 5031 11577 5043 11580
rect 4985 11571 5043 11577
rect 5629 11577 5641 11580
rect 5675 11577 5687 11611
rect 5629 11571 5687 11577
rect 7285 11611 7343 11617
rect 7285 11577 7297 11611
rect 7331 11608 7343 11611
rect 8496 11608 8524 11648
rect 8656 11639 8668 11648
rect 8662 11636 8668 11639
rect 8720 11636 8726 11688
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11514 11676 11520 11688
rect 10928 11648 11520 11676
rect 10928 11636 10934 11648
rect 11514 11636 11520 11648
rect 11572 11676 11578 11688
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 11572 11648 12173 11676
rect 11572 11636 11578 11648
rect 12161 11645 12173 11648
rect 12207 11645 12219 11679
rect 13170 11676 13176 11688
rect 13131 11648 13176 11676
rect 12161 11639 12219 11645
rect 13170 11636 13176 11648
rect 13228 11676 13234 11688
rect 13357 11679 13415 11685
rect 13357 11676 13369 11679
rect 13228 11648 13369 11676
rect 13228 11636 13234 11648
rect 13357 11645 13369 11648
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13613 11679 13671 11685
rect 13613 11676 13625 11679
rect 13504 11648 13625 11676
rect 13504 11636 13510 11648
rect 13613 11645 13625 11648
rect 13659 11645 13671 11679
rect 21174 11676 21180 11688
rect 21135 11648 21180 11676
rect 13613 11639 13671 11645
rect 21174 11636 21180 11648
rect 21232 11676 21238 11688
rect 21637 11679 21695 11685
rect 21637 11676 21649 11679
rect 21232 11648 21649 11676
rect 21232 11636 21238 11648
rect 21637 11645 21649 11648
rect 21683 11645 21695 11679
rect 21637 11639 21695 11645
rect 7331 11580 8524 11608
rect 11333 11611 11391 11617
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 11333 11577 11345 11611
rect 11379 11608 11391 11611
rect 13722 11608 13728 11620
rect 11379 11580 13728 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18049 11611 18107 11617
rect 18049 11608 18061 11611
rect 18012 11580 18061 11608
rect 18012 11568 18018 11580
rect 18049 11577 18061 11580
rect 18095 11577 18107 11611
rect 18049 11571 18107 11577
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 4706 11540 4712 11552
rect 2832 11512 4712 11540
rect 2832 11500 2838 11512
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 7892 11512 8125 11540
rect 7892 11500 7898 11512
rect 8113 11509 8125 11512
rect 8159 11540 8171 11543
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 8159 11512 8217 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 8205 11503 8263 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 10100 11512 10333 11540
rect 10100 11500 10106 11512
rect 10321 11509 10333 11512
rect 10367 11509 10379 11543
rect 11790 11540 11796 11552
rect 11751 11512 11796 11540
rect 10321 11503 10379 11509
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 13998 11540 14004 11552
rect 12943 11512 14004 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15102 11540 15108 11552
rect 14783 11512 15108 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15838 11540 15844 11552
rect 15799 11512 15844 11540
rect 15838 11500 15844 11512
rect 15896 11540 15902 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 15896 11512 16405 11540
rect 15896 11500 15902 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 17126 11540 17132 11552
rect 17087 11512 17132 11540
rect 16393 11503 16451 11509
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 22002 11540 22008 11552
rect 21963 11512 22008 11540
rect 22002 11500 22008 11512
rect 22060 11500 22066 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3234 11336 3240 11348
rect 2915 11308 3240 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5534 11336 5540 11348
rect 5307 11308 5540 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5534 11296 5540 11308
rect 5592 11336 5598 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 5592 11308 5641 11336
rect 5592 11296 5598 11308
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 6086 11336 6092 11348
rect 6047 11308 6092 11336
rect 5629 11299 5687 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7098 11336 7104 11348
rect 6963 11308 7104 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 8662 11336 8668 11348
rect 8527 11308 8668 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9861 11339 9919 11345
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 11790 11336 11796 11348
rect 9907 11308 11796 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13446 11336 13452 11348
rect 13311 11308 13452 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13722 11336 13728 11348
rect 13683 11308 13728 11336
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 14458 11336 14464 11348
rect 14419 11308 14464 11336
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15289 11339 15347 11345
rect 15289 11336 15301 11339
rect 14792 11308 15301 11336
rect 14792 11296 14798 11308
rect 15289 11305 15301 11308
rect 15335 11305 15347 11339
rect 16390 11336 16396 11348
rect 16351 11308 16396 11336
rect 15289 11299 15347 11305
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 17770 11336 17776 11348
rect 17731 11308 17776 11336
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 7374 11277 7380 11280
rect 7368 11268 7380 11277
rect 7287 11240 7380 11268
rect 7368 11231 7380 11240
rect 7432 11268 7438 11280
rect 8202 11268 8208 11280
rect 7432 11240 8208 11268
rect 7374 11228 7380 11231
rect 7432 11228 7438 11240
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 11140 11271 11198 11277
rect 11140 11237 11152 11271
rect 11186 11268 11198 11271
rect 11238 11268 11244 11280
rect 11186 11240 11244 11268
rect 11186 11237 11198 11240
rect 11140 11231 11198 11237
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 13464 11268 13492 11296
rect 13464 11240 13860 11268
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11200 2375 11203
rect 2406 11200 2412 11212
rect 2363 11172 2412 11200
rect 2363 11169 2375 11172
rect 2317 11163 2375 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4028 11172 4445 11200
rect 4028 11160 4034 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 4571 11172 6469 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1762 11132 1768 11144
rect 1443 11104 1768 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3421 11135 3479 11141
rect 3421 11132 3433 11135
rect 3099 11104 3433 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3421 11101 3433 11104
rect 3467 11132 3479 11135
rect 3602 11132 3608 11144
rect 3467 11104 3608 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4396 11104 4629 11132
rect 4396 11092 4402 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4062 11064 4068 11076
rect 4023 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 2409 10999 2467 11005
rect 2409 10965 2421 10999
rect 2455 10996 2467 10999
rect 4724 10996 4752 11172
rect 6457 11169 6469 11172
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10962 11200 10968 11212
rect 10459 11172 10968 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 13832 11200 13860 11240
rect 13832 11172 13952 11200
rect 13924 11144 13952 11172
rect 15286 11160 15292 11212
rect 15344 11200 15350 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15344 11172 15669 11200
rect 15344 11160 15350 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 17586 11200 17592 11212
rect 17547 11172 17592 11200
rect 15657 11163 15715 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 6914 11132 6920 11144
rect 6328 11104 6920 11132
rect 6328 11092 6334 11104
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6972 11104 7113 11132
rect 6972 11092 6978 11104
rect 7101 11101 7113 11104
rect 7147 11101 7159 11135
rect 7101 11095 7159 11101
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10836 11104 10885 11132
rect 10836 11092 10842 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 13078 11132 13084 11144
rect 12308 11104 13084 11132
rect 12308 11092 12314 11104
rect 13078 11092 13084 11104
rect 13136 11132 13142 11144
rect 13817 11135 13875 11141
rect 13817 11132 13829 11135
rect 13136 11104 13829 11132
rect 13136 11092 13142 11104
rect 13817 11101 13829 11104
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 13964 11104 14057 11132
rect 14936 11104 15761 11132
rect 13964 11092 13970 11104
rect 13354 11064 13360 11076
rect 13315 11036 13360 11064
rect 13354 11024 13360 11036
rect 13412 11024 13418 11076
rect 2455 10968 4752 10996
rect 2455 10965 2467 10968
rect 2409 10959 2467 10965
rect 11974 10956 11980 11008
rect 12032 10996 12038 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 12032 10968 12265 10996
rect 12032 10956 12038 10968
rect 12253 10965 12265 10968
rect 12299 10996 12311 10999
rect 12805 10999 12863 11005
rect 12805 10996 12817 10999
rect 12299 10968 12817 10996
rect 12299 10965 12311 10968
rect 12253 10959 12311 10965
rect 12805 10965 12817 10968
rect 12851 10965 12863 10999
rect 12805 10959 12863 10965
rect 13998 10956 14004 11008
rect 14056 10996 14062 11008
rect 14936 10996 14964 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16482 11132 16488 11144
rect 15979 11104 16488 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 15102 11064 15108 11076
rect 15015 11036 15108 11064
rect 15102 11024 15108 11036
rect 15160 11064 15166 11076
rect 15948 11064 15976 11095
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 15160 11036 15976 11064
rect 15160 11024 15166 11036
rect 14056 10968 14964 10996
rect 14056 10956 14062 10968
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1946 10792 1952 10804
rect 1688 10764 1952 10792
rect 1688 10665 1716 10764
rect 1946 10752 1952 10764
rect 2004 10752 2010 10804
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 2372 10764 3065 10792
rect 2372 10752 2378 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 3053 10755 3111 10761
rect 3697 10795 3755 10801
rect 3697 10761 3709 10795
rect 3743 10792 3755 10795
rect 4338 10792 4344 10804
rect 3743 10764 4344 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 3068 10656 3096 10755
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 6825 10795 6883 10801
rect 6825 10761 6837 10795
rect 6871 10792 6883 10795
rect 8297 10795 8355 10801
rect 8297 10792 8309 10795
rect 6871 10764 8309 10792
rect 6871 10761 6883 10764
rect 6825 10755 6883 10761
rect 8297 10761 8309 10764
rect 8343 10792 8355 10795
rect 8386 10792 8392 10804
rect 8343 10764 8392 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11238 10792 11244 10804
rect 11103 10764 11244 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 13906 10792 13912 10804
rect 13863 10764 13912 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15562 10792 15568 10804
rect 15243 10764 15568 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 16574 10792 16580 10804
rect 16535 10764 16580 10792
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17310 10792 17316 10804
rect 16991 10764 17316 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 19242 10792 19248 10804
rect 18555 10764 19248 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 6273 10727 6331 10733
rect 6273 10693 6285 10727
rect 6319 10724 6331 10727
rect 6319 10696 7420 10724
rect 6319 10693 6331 10696
rect 6273 10687 6331 10693
rect 7392 10668 7420 10696
rect 3068 10628 4292 10656
rect 1673 10619 1731 10625
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 3936 10560 4077 10588
rect 3936 10548 3942 10560
rect 4065 10557 4077 10560
rect 4111 10588 4123 10591
rect 4157 10591 4215 10597
rect 4157 10588 4169 10591
rect 4111 10560 4169 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4157 10557 4169 10560
rect 4203 10557 4215 10591
rect 4264 10588 4292 10628
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 7098 10656 7104 10668
rect 6788 10628 7104 10656
rect 6788 10616 6794 10628
rect 7098 10616 7104 10628
rect 7156 10656 7162 10668
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 7156 10628 7297 10656
rect 7156 10616 7162 10628
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7432 10628 7477 10656
rect 7432 10616 7438 10628
rect 13998 10616 14004 10668
rect 14056 10656 14062 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14056 10628 14657 10656
rect 14056 10616 14062 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 14645 10619 14703 10625
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10656 15899 10659
rect 16022 10656 16028 10668
rect 15887 10628 16028 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 16022 10616 16028 10628
rect 16080 10656 16086 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 16080 10628 16221 10656
rect 16080 10616 16086 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 4430 10597 4436 10600
rect 4413 10591 4436 10597
rect 4413 10588 4425 10591
rect 4264 10560 4425 10588
rect 4157 10551 4215 10557
rect 4413 10557 4425 10560
rect 4488 10588 4494 10600
rect 4488 10560 4561 10588
rect 4413 10551 4436 10557
rect 4430 10548 4436 10551
rect 4488 10548 4494 10560
rect 6638 10548 6644 10600
rect 6696 10588 6702 10600
rect 6914 10588 6920 10600
rect 6696 10560 6920 10588
rect 6696 10548 6702 10560
rect 6914 10548 6920 10560
rect 6972 10588 6978 10600
rect 7834 10588 7840 10600
rect 6972 10560 7840 10588
rect 6972 10548 6978 10560
rect 7834 10548 7840 10560
rect 7892 10588 7898 10600
rect 9490 10588 9496 10600
rect 7892 10560 9496 10588
rect 7892 10548 7898 10560
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10778 10588 10784 10600
rect 9732 10560 10784 10588
rect 9732 10548 9738 10560
rect 10778 10548 10784 10560
rect 10836 10588 10842 10600
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 10836 10560 11621 10588
rect 10836 10548 10842 10560
rect 11609 10557 11621 10560
rect 11655 10588 11667 10591
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 11655 10560 12173 10588
rect 11655 10557 11667 10560
rect 11609 10551 11667 10557
rect 12161 10557 12173 10560
rect 12207 10588 12219 10591
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 12207 10560 12449 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12437 10557 12449 10560
rect 12483 10588 12495 10591
rect 13170 10588 13176 10600
rect 12483 10560 13176 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 13170 10548 13176 10560
rect 13228 10548 13234 10600
rect 16758 10588 16764 10600
rect 16719 10560 16764 10588
rect 16758 10548 16764 10560
rect 16816 10588 16822 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 16816 10560 17233 10588
rect 16816 10548 16822 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17221 10551 17279 10557
rect 18230 10548 18236 10600
rect 18288 10588 18294 10600
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 18288 10560 18337 10588
rect 18288 10548 18294 10560
rect 18325 10557 18337 10560
rect 18371 10588 18383 10591
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18371 10560 18889 10588
rect 18371 10557 18383 10560
rect 18325 10551 18383 10557
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 1946 10529 1952 10532
rect 1940 10520 1952 10529
rect 1907 10492 1952 10520
rect 1940 10483 1952 10492
rect 1946 10480 1952 10483
rect 2004 10480 2010 10532
rect 9217 10523 9275 10529
rect 9217 10489 9229 10523
rect 9263 10520 9275 10523
rect 9766 10520 9772 10532
rect 9263 10492 9772 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 9766 10480 9772 10492
rect 9824 10520 9830 10532
rect 9944 10523 10002 10529
rect 9944 10520 9956 10523
rect 9824 10492 9956 10520
rect 9824 10480 9830 10492
rect 9944 10489 9956 10492
rect 9990 10520 10002 10523
rect 10134 10520 10140 10532
rect 9990 10492 10140 10520
rect 9990 10489 10002 10492
rect 9944 10483 10002 10489
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12682 10523 12740 10529
rect 12682 10520 12694 10523
rect 12032 10492 12694 10520
rect 12032 10480 12038 10492
rect 12682 10489 12694 10492
rect 12728 10489 12740 10523
rect 12682 10483 12740 10489
rect 15102 10480 15108 10532
rect 15160 10520 15166 10532
rect 15657 10523 15715 10529
rect 15657 10520 15669 10523
rect 15160 10492 15669 10520
rect 15160 10480 15166 10492
rect 15657 10489 15669 10492
rect 15703 10489 15715 10523
rect 15657 10483 15715 10489
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10452 6610 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 6604 10424 7205 10452
rect 6604 10412 6610 10424
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 7193 10415 7251 10421
rect 14826 10412 14832 10464
rect 14884 10452 14890 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14884 10424 15025 10452
rect 14884 10412 14890 10424
rect 15013 10421 15025 10424
rect 15059 10452 15071 10455
rect 15286 10452 15292 10464
rect 15059 10424 15292 10452
rect 15059 10421 15071 10424
rect 15013 10415 15071 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 17586 10452 17592 10464
rect 17547 10424 17592 10452
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 2832 10220 2877 10248
rect 2832 10208 2838 10220
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3200 10220 3801 10248
rect 3200 10208 3206 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 4488 10220 4537 10248
rect 4488 10208 4494 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 7193 10251 7251 10257
rect 7193 10217 7205 10251
rect 7239 10248 7251 10251
rect 7374 10248 7380 10260
rect 7239 10220 7380 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7650 10248 7656 10260
rect 7611 10220 7656 10248
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 7834 10208 7840 10260
rect 7892 10248 7898 10260
rect 8110 10248 8116 10260
rect 7892 10220 8116 10248
rect 7892 10208 7898 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10870 10248 10876 10260
rect 9723 10220 10876 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11241 10251 11299 10257
rect 11241 10217 11253 10251
rect 11287 10248 11299 10251
rect 12250 10248 12256 10260
rect 11287 10220 12256 10248
rect 11287 10217 11299 10220
rect 11241 10211 11299 10217
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 13541 10251 13599 10257
rect 13541 10217 13553 10251
rect 13587 10248 13599 10251
rect 15102 10248 15108 10260
rect 13587 10220 15108 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15562 10248 15568 10260
rect 15523 10220 15568 10248
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 17126 10248 17132 10260
rect 17087 10220 17132 10248
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 1762 10180 1768 10192
rect 1723 10152 1768 10180
rect 1762 10140 1768 10152
rect 1820 10140 1826 10192
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10180 2559 10183
rect 3234 10180 3240 10192
rect 2547 10152 3240 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 3510 10180 3516 10192
rect 3471 10152 3516 10180
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 4338 10140 4344 10192
rect 4396 10180 4402 10192
rect 5350 10180 5356 10192
rect 4396 10152 5356 10180
rect 4396 10140 4402 10152
rect 5350 10140 5356 10152
rect 5408 10189 5414 10192
rect 5408 10183 5472 10189
rect 5408 10149 5426 10183
rect 5460 10149 5472 10183
rect 5408 10143 5472 10149
rect 5408 10140 5414 10143
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 8846 10140 8852 10192
rect 8904 10180 8910 10192
rect 11698 10180 11704 10192
rect 8904 10152 11704 10180
rect 8904 10140 8910 10152
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 13449 10183 13507 10189
rect 13449 10149 13461 10183
rect 13495 10180 13507 10183
rect 13722 10180 13728 10192
rect 13495 10152 13728 10180
rect 13495 10149 13507 10152
rect 13449 10143 13507 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 13998 10180 14004 10192
rect 13959 10152 14004 10180
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 16022 10189 16028 10192
rect 16016 10180 16028 10189
rect 15983 10152 16028 10180
rect 16016 10143 16028 10152
rect 16022 10140 16028 10143
rect 16080 10140 16086 10192
rect 2958 10112 2964 10124
rect 2871 10084 2964 10112
rect 2958 10072 2964 10084
rect 3016 10112 3022 10124
rect 3418 10112 3424 10124
rect 3016 10084 3424 10112
rect 3016 10072 3022 10084
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 8018 10112 8024 10124
rect 7979 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8220 10112 8248 10140
rect 8665 10115 8723 10121
rect 8665 10112 8677 10115
rect 8220 10084 8677 10112
rect 8665 10081 8677 10084
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9732 10084 10057 10112
rect 9732 10072 9738 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 11238 10112 11244 10124
rect 11011 10084 11244 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 11609 10115 11667 10121
rect 11609 10112 11621 10115
rect 11572 10084 11621 10112
rect 11572 10072 11578 10084
rect 11609 10081 11621 10084
rect 11655 10081 11667 10115
rect 11609 10075 11667 10081
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 13872 10084 13921 10112
rect 13872 10072 13878 10084
rect 13909 10081 13921 10084
rect 13955 10081 13967 10115
rect 13909 10075 13967 10081
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15746 10112 15752 10124
rect 15528 10084 15752 10112
rect 15528 10072 15534 10084
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 1946 10044 1952 10056
rect 1907 10016 1952 10044
rect 1946 10004 1952 10016
rect 2004 10044 2010 10056
rect 3142 10044 3148 10056
rect 2004 10016 3148 10044
rect 2004 10004 2010 10016
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 4154 10044 4160 10056
rect 4111 10016 4160 10044
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 5166 10044 5172 10056
rect 5127 10016 5172 10044
rect 5166 10004 5172 10016
rect 5224 10004 5230 10056
rect 8202 10044 8208 10056
rect 8115 10016 8208 10044
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 9456 10016 10149 10044
rect 9456 10004 9462 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10137 10007 10195 10013
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 11974 10044 11980 10056
rect 11931 10016 11980 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 1397 9979 1455 9985
rect 1397 9945 1409 9979
rect 1443 9976 1455 9979
rect 2222 9976 2228 9988
rect 1443 9948 2228 9976
rect 1443 9945 1455 9948
rect 1397 9939 1455 9945
rect 2222 9936 2228 9948
rect 2280 9976 2286 9988
rect 4893 9979 4951 9985
rect 4893 9976 4905 9979
rect 2280 9948 4905 9976
rect 2280 9936 2286 9948
rect 4893 9945 4905 9948
rect 4939 9945 4951 9979
rect 4893 9939 4951 9945
rect 7561 9979 7619 9985
rect 7561 9945 7573 9979
rect 7607 9976 7619 9979
rect 8211 9976 8239 10004
rect 7607 9948 8239 9976
rect 13081 9979 13139 9985
rect 7607 9945 7619 9948
rect 7561 9939 7619 9945
rect 13081 9945 13093 9979
rect 13127 9976 13139 9979
rect 14108 9976 14136 10007
rect 14550 9976 14556 9988
rect 13127 9948 14556 9976
rect 13127 9945 13139 9948
rect 13081 9939 13139 9945
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 3145 9911 3203 9917
rect 3145 9877 3157 9911
rect 3191 9908 3203 9911
rect 5074 9908 5080 9920
rect 3191 9880 5080 9908
rect 3191 9877 3203 9880
rect 3145 9871 3203 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 6546 9908 6552 9920
rect 6507 9880 6552 9908
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12802 9908 12808 9920
rect 12575 9880 12808 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 1949 9707 2007 9713
rect 1949 9704 1961 9707
rect 1912 9676 1961 9704
rect 1912 9664 1918 9676
rect 1949 9673 1961 9676
rect 1995 9673 2007 9707
rect 1949 9667 2007 9673
rect 3513 9707 3571 9713
rect 3513 9673 3525 9707
rect 3559 9704 3571 9707
rect 3602 9704 3608 9716
rect 3559 9676 3608 9704
rect 3559 9673 3571 9676
rect 3513 9667 3571 9673
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 3878 9704 3884 9716
rect 3839 9676 3884 9704
rect 3878 9664 3884 9676
rect 3936 9704 3942 9716
rect 4706 9704 4712 9716
rect 3936 9676 4712 9704
rect 3936 9664 3942 9676
rect 4706 9664 4712 9676
rect 4764 9704 4770 9716
rect 5166 9704 5172 9716
rect 4764 9676 5172 9704
rect 4764 9664 4770 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5350 9704 5356 9716
rect 5311 9676 5356 9704
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 8202 9704 8208 9716
rect 8163 9676 8208 9704
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 10318 9664 10324 9716
rect 10376 9704 10382 9716
rect 11057 9707 11115 9713
rect 11057 9704 11069 9707
rect 10376 9676 11069 9704
rect 10376 9664 10382 9676
rect 11057 9673 11069 9676
rect 11103 9673 11115 9707
rect 11057 9667 11115 9673
rect 11698 9664 11704 9716
rect 11756 9704 11762 9716
rect 12069 9707 12127 9713
rect 12069 9704 12081 9707
rect 11756 9676 12081 9704
rect 11756 9664 11762 9676
rect 12069 9673 12081 9676
rect 12115 9673 12127 9707
rect 13998 9704 14004 9716
rect 13959 9676 14004 9704
rect 12069 9667 12127 9673
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 15841 9707 15899 9713
rect 15841 9673 15853 9707
rect 15887 9704 15899 9707
rect 16022 9704 16028 9716
rect 15887 9676 16028 9704
rect 15887 9673 15899 9676
rect 15841 9667 15899 9673
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 17129 9707 17187 9713
rect 17129 9673 17141 9707
rect 17175 9704 17187 9707
rect 17586 9704 17592 9716
rect 17175 9676 17592 9704
rect 17175 9673 17187 9676
rect 17129 9667 17187 9673
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 18230 9704 18236 9716
rect 18191 9676 18236 9704
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 1486 9596 1492 9648
rect 1544 9636 1550 9648
rect 1581 9639 1639 9645
rect 1581 9636 1593 9639
rect 1544 9608 1593 9636
rect 1544 9596 1550 9608
rect 1581 9605 1593 9608
rect 1627 9605 1639 9639
rect 1581 9599 1639 9605
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 2317 9639 2375 9645
rect 2317 9636 2329 9639
rect 1820 9608 2329 9636
rect 1820 9596 1826 9608
rect 2317 9605 2329 9608
rect 2363 9605 2375 9639
rect 2317 9599 2375 9605
rect 2406 9596 2412 9648
rect 2464 9636 2470 9648
rect 2685 9639 2743 9645
rect 2685 9636 2697 9639
rect 2464 9608 2697 9636
rect 2464 9596 2470 9608
rect 2685 9605 2697 9608
rect 2731 9605 2743 9639
rect 2685 9599 2743 9605
rect 3620 9568 3648 9664
rect 5184 9568 5212 9664
rect 9674 9636 9680 9648
rect 9635 9608 9680 9636
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 12342 9636 12348 9648
rect 11204 9608 12348 9636
rect 11204 9596 11210 9608
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 12860 9608 13032 9636
rect 12860 9596 12866 9608
rect 10321 9571 10379 9577
rect 2424 9540 3096 9568
rect 3620 9540 4108 9568
rect 5184 9540 6040 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 2314 9500 2320 9512
rect 1443 9472 2320 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2424 9500 2452 9540
rect 2493 9503 2551 9509
rect 2493 9500 2505 9503
rect 2424 9472 2505 9500
rect 2493 9469 2505 9472
rect 2539 9469 2551 9503
rect 2493 9463 2551 9469
rect 3068 9441 3096 9540
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3936 9472 3985 9500
rect 3936 9460 3942 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 4080 9500 4108 9540
rect 4229 9503 4287 9509
rect 4229 9500 4241 9503
rect 4080 9472 4241 9500
rect 3973 9463 4031 9469
rect 4229 9469 4241 9472
rect 4275 9500 4287 9503
rect 4614 9500 4620 9512
rect 4275 9472 4620 9500
rect 4275 9469 4287 9472
rect 4229 9463 4287 9469
rect 4614 9460 4620 9472
rect 4672 9500 4678 9512
rect 5442 9500 5448 9512
rect 4672 9472 5448 9500
rect 4672 9460 4678 9472
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6012 9509 6040 9540
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10686 9568 10692 9580
rect 10367 9540 10692 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 13004 9577 13032 9608
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 16393 9639 16451 9645
rect 16393 9636 16405 9639
rect 15804 9608 16405 9636
rect 15804 9596 15810 9608
rect 16393 9605 16405 9608
rect 16439 9605 16451 9639
rect 16393 9599 16451 9605
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9500 6055 9503
rect 6638 9500 6644 9512
rect 6043 9472 6644 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6638 9460 6644 9472
rect 6696 9500 6702 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6696 9472 6837 9500
rect 6696 9460 6702 9472
rect 6825 9469 6837 9472
rect 6871 9500 6883 9503
rect 7926 9500 7932 9512
rect 6871 9472 7932 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 12894 9500 12900 9512
rect 12851 9472 12900 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 3053 9435 3111 9441
rect 3053 9401 3065 9435
rect 3099 9432 3111 9435
rect 3099 9404 4292 9432
rect 3099 9401 3111 9404
rect 3053 9395 3111 9401
rect 4264 9376 4292 9404
rect 7006 9392 7012 9444
rect 7064 9441 7070 9444
rect 7064 9435 7128 9441
rect 7064 9401 7082 9435
rect 7116 9401 7128 9435
rect 7064 9395 7128 9401
rect 8849 9435 8907 9441
rect 8849 9401 8861 9435
rect 8895 9432 8907 9435
rect 10045 9435 10103 9441
rect 10045 9432 10057 9435
rect 8895 9404 10057 9432
rect 8895 9401 8907 9404
rect 8849 9395 8907 9401
rect 10045 9401 10057 9404
rect 10091 9432 10103 9435
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 10091 9404 11253 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 11241 9401 11253 9404
rect 11287 9401 11299 9435
rect 11241 9395 11299 9401
rect 7064 9392 7070 9395
rect 12710 9392 12716 9444
rect 12768 9432 12774 9444
rect 14369 9435 14427 9441
rect 14369 9432 14381 9435
rect 12768 9404 14381 9432
rect 12768 9392 12774 9404
rect 14369 9401 14381 9404
rect 14415 9432 14427 9435
rect 14476 9432 14504 9463
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 14717 9503 14775 9509
rect 14717 9500 14729 9503
rect 14608 9472 14729 9500
rect 14608 9460 14614 9472
rect 14717 9469 14729 9472
rect 14763 9469 14775 9503
rect 16942 9500 16948 9512
rect 16903 9472 16948 9500
rect 14717 9463 14775 9469
rect 16942 9460 16948 9472
rect 17000 9500 17006 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 17000 9472 17417 9500
rect 17000 9460 17006 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 17405 9463 17463 9469
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18509 9503 18567 9509
rect 18509 9500 18521 9503
rect 18104 9472 18521 9500
rect 18104 9460 18110 9472
rect 18509 9469 18521 9472
rect 18555 9469 18567 9503
rect 18509 9463 18567 9469
rect 15746 9432 15752 9444
rect 14415 9404 15752 9432
rect 14415 9401 14427 9404
rect 14369 9395 14427 9401
rect 15746 9392 15752 9404
rect 15804 9392 15810 9444
rect 4246 9324 4252 9376
rect 4304 9324 4310 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 9125 9367 9183 9373
rect 9125 9364 9137 9367
rect 8536 9336 9137 9364
rect 8536 9324 8542 9336
rect 9125 9333 9137 9336
rect 9171 9364 9183 9367
rect 9398 9364 9404 9376
rect 9171 9336 9404 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 10134 9364 10140 9376
rect 9548 9336 9593 9364
rect 10095 9336 10140 9364
rect 9548 9324 9554 9336
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10686 9364 10692 9376
rect 10647 9336 10692 9364
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 11572 9336 11713 9364
rect 11572 9324 11578 9336
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 11701 9327 11759 9333
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12897 9367 12955 9373
rect 12492 9336 12537 9364
rect 12492 9324 12498 9336
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 12986 9364 12992 9376
rect 12943 9336 12992 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13504 9336 13553 9364
rect 13504 9324 13510 9336
rect 13541 9333 13553 9336
rect 13587 9364 13599 9367
rect 13814 9364 13820 9376
rect 13587 9336 13820 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1854 9160 1860 9172
rect 1815 9132 1860 9160
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2590 9160 2596 9172
rect 2551 9132 2596 9160
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3329 9163 3387 9169
rect 3329 9160 3341 9163
rect 2740 9132 3341 9160
rect 2740 9120 2746 9132
rect 3329 9129 3341 9132
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 3881 9163 3939 9169
rect 3881 9129 3893 9163
rect 3927 9160 3939 9163
rect 3970 9160 3976 9172
rect 3927 9132 3976 9160
rect 3927 9129 3939 9132
rect 3881 9123 3939 9129
rect 3970 9120 3976 9132
rect 4028 9160 4034 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 4028 9132 4077 9160
rect 4028 9120 4034 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4212 9132 4445 9160
rect 4212 9120 4218 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 5261 9163 5319 9169
rect 4580 9132 4625 9160
rect 4580 9120 4586 9132
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 5350 9160 5356 9172
rect 5307 9132 5356 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 6972 9132 7757 9160
rect 6972 9120 6978 9132
rect 7745 9129 7757 9132
rect 7791 9160 7803 9163
rect 8018 9160 8024 9172
rect 7791 9132 8024 9160
rect 7791 9129 7803 9132
rect 7745 9123 7803 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 10134 9160 10140 9172
rect 9539 9132 10140 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 2958 9092 2964 9104
rect 2919 9064 2964 9092
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 6362 9092 6368 9104
rect 6323 9064 6368 9092
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 6457 9095 6515 9101
rect 6457 9061 6469 9095
rect 6503 9092 6515 9095
rect 6730 9092 6736 9104
rect 6503 9064 6736 9092
rect 6503 9061 6515 9064
rect 6457 9055 6515 9061
rect 6730 9052 6736 9064
rect 6788 9052 6794 9104
rect 7466 9052 7472 9104
rect 7524 9092 7530 9104
rect 8478 9092 8484 9104
rect 7524 9064 8484 9092
rect 7524 9052 7530 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 9508 9092 9536 9123
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 14645 9163 14703 9169
rect 14645 9160 14657 9163
rect 13044 9132 14657 9160
rect 13044 9120 13050 9132
rect 14645 9129 14657 9132
rect 14691 9129 14703 9163
rect 14645 9123 14703 9129
rect 15381 9163 15439 9169
rect 15381 9129 15393 9163
rect 15427 9160 15439 9163
rect 15562 9160 15568 9172
rect 15427 9132 15568 9160
rect 15427 9129 15439 9132
rect 15381 9123 15439 9129
rect 15562 9120 15568 9132
rect 15620 9120 15626 9172
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16022 9160 16028 9172
rect 15979 9132 16028 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 16666 9160 16672 9172
rect 16623 9132 16672 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 8588 9064 9536 9092
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1946 9024 1952 9036
rect 1443 8996 1952 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 2130 8984 2136 9036
rect 2188 9024 2194 9036
rect 2409 9027 2467 9033
rect 2409 9024 2421 9027
rect 2188 8996 2421 9024
rect 2188 8984 2194 8996
rect 2409 8993 2421 8996
rect 2455 8993 2467 9027
rect 2409 8987 2467 8993
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 7800 8996 8401 9024
rect 7800 8984 7806 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 4614 8956 4620 8968
rect 4575 8928 4620 8956
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 7006 8956 7012 8968
rect 6604 8928 7012 8956
rect 6604 8916 6610 8928
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 1581 8891 1639 8897
rect 1581 8857 1593 8891
rect 1627 8888 1639 8891
rect 2498 8888 2504 8900
rect 1627 8860 2504 8888
rect 1627 8857 1639 8860
rect 1581 8851 1639 8857
rect 2498 8848 2504 8860
rect 2556 8848 2562 8900
rect 5997 8891 6055 8897
rect 5997 8857 6009 8891
rect 6043 8888 6055 8891
rect 7834 8888 7840 8900
rect 6043 8860 7840 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 8021 8891 8079 8897
rect 8021 8857 8033 8891
rect 8067 8888 8079 8891
rect 8588 8888 8616 9064
rect 9950 9033 9956 9036
rect 9944 9024 9956 9033
rect 8680 8996 9956 9024
rect 8680 8965 8708 8996
rect 9944 8987 9956 8996
rect 10008 9024 10014 9036
rect 10008 8996 10044 9024
rect 9950 8984 9956 8987
rect 10008 8984 10014 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12710 9024 12716 9036
rect 12492 8996 12716 9024
rect 12492 8984 12498 8996
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 12969 9027 13027 9033
rect 12969 9024 12981 9027
rect 12860 8996 12981 9024
rect 12860 8984 12866 8996
rect 12969 8993 12981 8996
rect 13015 8993 13027 9027
rect 16390 9024 16396 9036
rect 16351 8996 16396 9024
rect 12969 8987 13027 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 8665 8959 8723 8965
rect 8665 8925 8677 8959
rect 8711 8925 8723 8959
rect 8665 8919 8723 8925
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9732 8928 9777 8956
rect 9732 8916 9738 8928
rect 8067 8860 8616 8888
rect 14093 8891 14151 8897
rect 8067 8857 8079 8860
rect 8021 8851 8079 8857
rect 14093 8857 14105 8891
rect 14139 8888 14151 8891
rect 14550 8888 14556 8900
rect 14139 8860 14556 8888
rect 14139 8857 14151 8860
rect 14093 8851 14151 8857
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10744 8792 11069 8820
rect 10744 8780 10750 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11606 8820 11612 8832
rect 11567 8792 11612 8820
rect 11057 8783 11115 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12529 8823 12587 8829
rect 12529 8789 12541 8823
rect 12575 8820 12587 8823
rect 12894 8820 12900 8832
rect 12575 8792 12900 8820
rect 12575 8789 12587 8792
rect 12529 8783 12587 8789
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2188 8588 2421 8616
rect 2188 8576 2194 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4212 8588 4445 8616
rect 4212 8576 4218 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4672 8588 4813 8616
rect 4672 8576 4678 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 6546 8616 6552 8628
rect 5767 8588 6552 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7466 8616 7472 8628
rect 7427 8588 7472 8616
rect 7466 8576 7472 8588
rect 7524 8576 7530 8628
rect 7742 8616 7748 8628
rect 7703 8588 7748 8616
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12802 8616 12808 8628
rect 11931 8588 12808 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12802 8576 12808 8588
rect 12860 8616 12866 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 12860 8588 13829 8616
rect 12860 8576 12866 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 16390 8616 16396 8628
rect 16351 8588 16396 8616
rect 13817 8579 13875 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 1670 8548 1676 8560
rect 1631 8520 1676 8548
rect 1670 8508 1676 8520
rect 1728 8508 1734 8560
rect 6089 8551 6147 8557
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 6362 8548 6368 8560
rect 6135 8520 6368 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 6362 8508 6368 8520
rect 6420 8508 6426 8560
rect 6457 8551 6515 8557
rect 6457 8517 6469 8551
rect 6503 8548 6515 8551
rect 6730 8548 6736 8560
rect 6503 8520 6736 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 9950 8548 9956 8560
rect 9355 8520 9956 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 10321 8551 10379 8557
rect 10321 8517 10333 8551
rect 10367 8548 10379 8551
rect 11698 8548 11704 8560
rect 10367 8520 11704 8548
rect 10367 8517 10379 8520
rect 10321 8511 10379 8517
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4522 8480 4528 8492
rect 4203 8452 4528 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 11256 8489 11284 8520
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8480 11299 8483
rect 11425 8483 11483 8489
rect 11287 8452 11321 8480
rect 11287 8449 11299 8452
rect 11241 8443 11299 8449
rect 11425 8449 11437 8483
rect 11471 8480 11483 8483
rect 11606 8480 11612 8492
rect 11471 8452 11612 8480
rect 11471 8449 11483 8452
rect 11425 8443 11483 8449
rect 11606 8440 11612 8452
rect 11664 8480 11670 8492
rect 11664 8452 12572 8480
rect 11664 8440 11670 8452
rect 1489 8415 1547 8421
rect 1489 8381 1501 8415
rect 1535 8412 1547 8415
rect 2038 8412 2044 8424
rect 1535 8384 2044 8412
rect 1535 8381 1547 8384
rect 1489 8375 1547 8381
rect 2038 8372 2044 8384
rect 2096 8372 2102 8424
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8202 8421 8208 8424
rect 8196 8412 8208 8421
rect 8163 8384 8208 8412
rect 8196 8375 8208 8384
rect 8202 8372 8208 8375
rect 8260 8372 8266 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12434 8412 12440 8424
rect 12299 8384 12440 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12544 8412 12572 8452
rect 12693 8415 12751 8421
rect 12693 8412 12705 8415
rect 12544 8384 12705 8412
rect 12693 8381 12705 8384
rect 12739 8381 12751 8415
rect 12693 8375 12751 8381
rect 10594 8344 10600 8356
rect 10555 8316 10600 8344
rect 10594 8304 10600 8316
rect 10652 8344 10658 8356
rect 11149 8347 11207 8353
rect 11149 8344 11161 8347
rect 10652 8316 11161 8344
rect 10652 8304 10658 8316
rect 11149 8313 11161 8316
rect 11195 8313 11207 8347
rect 11149 8307 11207 8313
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9732 8248 9965 8276
rect 9732 8236 9738 8248
rect 9953 8245 9965 8248
rect 9999 8276 10011 8279
rect 10134 8276 10140 8288
rect 9999 8248 10140 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 1946 8072 1952 8084
rect 1719 8044 1952 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 7926 8072 7932 8084
rect 7887 8044 7932 8072
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8294 8072 8300 8084
rect 8255 8044 8300 8072
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9950 8072 9956 8084
rect 8803 8044 9956 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 11793 8075 11851 8081
rect 11793 8072 11805 8075
rect 11664 8044 11805 8072
rect 11664 8032 11670 8044
rect 11793 8041 11805 8044
rect 11839 8072 11851 8075
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11839 8044 12357 8072
rect 11839 8041 11851 8044
rect 11793 8035 11851 8041
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12492 8044 12725 8072
rect 12492 8032 12498 8044
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 12894 8072 12900 8084
rect 12855 8044 12900 8072
rect 12713 8035 12771 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 10134 7964 10140 8016
rect 10192 8004 10198 8016
rect 12452 8004 12480 8032
rect 10192 7976 12480 8004
rect 10192 7964 10198 7976
rect 10428 7948 10456 7976
rect 10410 7936 10416 7948
rect 10323 7908 10416 7936
rect 10410 7896 10416 7908
rect 10468 7896 10474 7948
rect 10686 7945 10692 7948
rect 10680 7936 10692 7945
rect 10647 7908 10692 7936
rect 10680 7899 10692 7908
rect 10686 7896 10692 7899
rect 10744 7896 10750 7948
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 10410 7528 10416 7540
rect 10371 7500 10416 7528
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 10781 7531 10839 7537
rect 10781 7528 10793 7531
rect 10744 7500 10793 7528
rect 10744 7488 10750 7500
rect 10781 7497 10793 7500
rect 10827 7497 10839 7531
rect 10781 7491 10839 7497
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 9490 6440 9496 6452
rect 4856 6412 9496 6440
rect 4856 6400 4862 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9950 5769 9956 5772
rect 9944 5760 9956 5769
rect 9732 5732 9777 5760
rect 9911 5732 9956 5760
rect 9732 5720 9738 5732
rect 9944 5723 9956 5732
rect 9950 5720 9956 5723
rect 10008 5720 10014 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9732 5324 10057 5352
rect 9732 5312 9738 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 9950 5012 9956 5024
rect 9815 4984 9956 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9950 4972 9956 4984
rect 10008 5012 10014 5024
rect 13906 5012 13912 5024
rect 10008 4984 13912 5012
rect 10008 4972 10014 4984
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 3332 25372 3384 25424
rect 1860 25304 1912 25356
rect 2320 25304 2372 25356
rect 3056 25347 3108 25356
rect 3056 25313 3065 25347
rect 3065 25313 3099 25347
rect 3099 25313 3108 25347
rect 3056 25304 3108 25313
rect 4712 25347 4764 25356
rect 4712 25313 4721 25347
rect 4721 25313 4755 25347
rect 4755 25313 4764 25347
rect 4712 25304 4764 25313
rect 4804 25279 4856 25288
rect 4804 25245 4813 25279
rect 4813 25245 4847 25279
rect 4847 25245 4856 25279
rect 4804 25236 4856 25245
rect 4988 25279 5040 25288
rect 4988 25245 4997 25279
rect 4997 25245 5031 25279
rect 5031 25245 5040 25279
rect 4988 25236 5040 25245
rect 6920 25279 6972 25288
rect 6920 25245 6929 25279
rect 6929 25245 6963 25279
rect 6963 25245 6972 25279
rect 6920 25236 6972 25245
rect 2964 25168 3016 25220
rect 9128 25168 9180 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 2872 25100 2924 25152
rect 8392 25143 8444 25152
rect 8392 25109 8401 25143
rect 8401 25109 8435 25143
rect 8435 25109 8444 25143
rect 8392 25100 8444 25109
rect 13084 25100 13136 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 1860 24871 1912 24880
rect 1860 24837 1869 24871
rect 1869 24837 1903 24871
rect 1903 24837 1912 24871
rect 1860 24828 1912 24837
rect 2320 24871 2372 24880
rect 2320 24837 2329 24871
rect 2329 24837 2363 24871
rect 2363 24837 2372 24871
rect 2320 24828 2372 24837
rect 5356 24828 5408 24880
rect 2964 24760 3016 24812
rect 1676 24692 1728 24744
rect 2780 24735 2832 24744
rect 2780 24701 2789 24735
rect 2789 24701 2823 24735
rect 2823 24701 2832 24735
rect 2780 24692 2832 24701
rect 3240 24692 3292 24744
rect 3424 24692 3476 24744
rect 4712 24760 4764 24812
rect 8208 24760 8260 24812
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 12256 24803 12308 24812
rect 8392 24760 8444 24769
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 3056 24624 3108 24676
rect 6184 24735 6236 24744
rect 6184 24701 6193 24735
rect 6193 24701 6227 24735
rect 6227 24701 6236 24735
rect 6184 24692 6236 24701
rect 9312 24692 9364 24744
rect 9496 24624 9548 24676
rect 11796 24667 11848 24676
rect 11796 24633 11805 24667
rect 11805 24633 11839 24667
rect 11839 24633 11848 24667
rect 11796 24624 11848 24633
rect 1768 24556 1820 24608
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 3976 24599 4028 24608
rect 3976 24565 3985 24599
rect 3985 24565 4019 24599
rect 4019 24565 4028 24599
rect 3976 24556 4028 24565
rect 4436 24599 4488 24608
rect 4436 24565 4445 24599
rect 4445 24565 4479 24599
rect 4479 24565 4488 24599
rect 4436 24556 4488 24565
rect 5540 24556 5592 24608
rect 7840 24599 7892 24608
rect 7840 24565 7849 24599
rect 7849 24565 7883 24599
rect 7883 24565 7892 24599
rect 7840 24556 7892 24565
rect 7932 24556 7984 24608
rect 9312 24556 9364 24608
rect 9680 24556 9732 24608
rect 12532 24556 12584 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 2412 24352 2464 24404
rect 2596 24395 2648 24404
rect 2596 24361 2605 24395
rect 2605 24361 2639 24395
rect 2639 24361 2648 24395
rect 2596 24352 2648 24361
rect 3976 24352 4028 24404
rect 8024 24395 8076 24404
rect 8024 24361 8033 24395
rect 8033 24361 8067 24395
rect 8067 24361 8076 24395
rect 8024 24352 8076 24361
rect 9772 24352 9824 24404
rect 10968 24352 11020 24404
rect 15660 24395 15712 24404
rect 15660 24361 15669 24395
rect 15669 24361 15703 24395
rect 15703 24361 15712 24395
rect 15660 24352 15712 24361
rect 17316 24395 17368 24404
rect 17316 24361 17325 24395
rect 17325 24361 17359 24395
rect 17359 24361 17368 24395
rect 17316 24352 17368 24361
rect 21824 24395 21876 24404
rect 21824 24361 21833 24395
rect 21833 24361 21867 24395
rect 21867 24361 21876 24395
rect 21824 24352 21876 24361
rect 25320 24352 25372 24404
rect 3240 24327 3292 24336
rect 3240 24293 3249 24327
rect 3249 24293 3283 24327
rect 3283 24293 3292 24327
rect 3240 24284 3292 24293
rect 4804 24284 4856 24336
rect 11612 24284 11664 24336
rect 5080 24259 5132 24268
rect 5080 24225 5114 24259
rect 5114 24225 5132 24259
rect 5080 24216 5132 24225
rect 7012 24216 7064 24268
rect 9588 24216 9640 24268
rect 15384 24216 15436 24268
rect 17132 24259 17184 24268
rect 17132 24225 17141 24259
rect 17141 24225 17175 24259
rect 17175 24225 17184 24259
rect 17132 24216 17184 24225
rect 21640 24259 21692 24268
rect 21640 24225 21649 24259
rect 21649 24225 21683 24259
rect 21683 24225 21692 24259
rect 21640 24216 21692 24225
rect 23296 24259 23348 24268
rect 23296 24225 23305 24259
rect 23305 24225 23339 24259
rect 23339 24225 23348 24259
rect 23296 24216 23348 24225
rect 4620 24148 4672 24200
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 8392 24148 8444 24200
rect 10324 24191 10376 24200
rect 10324 24157 10333 24191
rect 10333 24157 10367 24191
rect 10367 24157 10376 24191
rect 11428 24191 11480 24200
rect 10324 24148 10376 24157
rect 2688 24080 2740 24132
rect 7564 24123 7616 24132
rect 7564 24089 7573 24123
rect 7573 24089 7607 24123
rect 7607 24089 7616 24123
rect 7564 24080 7616 24089
rect 1676 24055 1728 24064
rect 1676 24021 1685 24055
rect 1685 24021 1719 24055
rect 1719 24021 1728 24055
rect 1676 24012 1728 24021
rect 2228 24055 2280 24064
rect 2228 24021 2237 24055
rect 2237 24021 2271 24055
rect 2271 24021 2280 24055
rect 2228 24012 2280 24021
rect 4712 24012 4764 24064
rect 4988 24012 5040 24064
rect 7748 24012 7800 24064
rect 10140 24012 10192 24064
rect 11428 24157 11437 24191
rect 11437 24157 11471 24191
rect 11471 24157 11480 24191
rect 11428 24148 11480 24157
rect 13912 24055 13964 24064
rect 13912 24021 13921 24055
rect 13921 24021 13955 24055
rect 13955 24021 13964 24055
rect 13912 24012 13964 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 4160 23808 4212 23860
rect 2412 23604 2464 23656
rect 4160 23604 4212 23656
rect 2688 23536 2740 23588
rect 4804 23808 4856 23860
rect 6460 23851 6512 23860
rect 6460 23817 6469 23851
rect 6469 23817 6503 23851
rect 6503 23817 6512 23851
rect 6460 23808 6512 23817
rect 7012 23851 7064 23860
rect 7012 23817 7021 23851
rect 7021 23817 7055 23851
rect 7055 23817 7064 23851
rect 7012 23808 7064 23817
rect 9588 23808 9640 23860
rect 9772 23851 9824 23860
rect 9772 23817 9781 23851
rect 9781 23817 9815 23851
rect 9815 23817 9824 23851
rect 9772 23808 9824 23817
rect 16488 23851 16540 23860
rect 16488 23817 16497 23851
rect 16497 23817 16531 23851
rect 16531 23817 16540 23851
rect 16488 23808 16540 23817
rect 18420 23851 18472 23860
rect 18420 23817 18429 23851
rect 18429 23817 18463 23851
rect 18463 23817 18472 23851
rect 18420 23808 18472 23817
rect 19524 23851 19576 23860
rect 19524 23817 19533 23851
rect 19533 23817 19567 23851
rect 19567 23817 19576 23851
rect 19524 23808 19576 23817
rect 20628 23851 20680 23860
rect 20628 23817 20637 23851
rect 20637 23817 20671 23851
rect 20671 23817 20680 23851
rect 20628 23808 20680 23817
rect 21732 23851 21784 23860
rect 21732 23817 21741 23851
rect 21741 23817 21775 23851
rect 21775 23817 21784 23851
rect 21732 23808 21784 23817
rect 24768 23808 24820 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 5080 23672 5132 23724
rect 8024 23740 8076 23792
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 8668 23672 8720 23724
rect 9312 23672 9364 23724
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 15476 23672 15528 23724
rect 16212 23672 16264 23724
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 7564 23647 7616 23656
rect 7564 23613 7573 23647
rect 7573 23613 7607 23647
rect 7607 23613 7616 23647
rect 7564 23604 7616 23613
rect 7840 23604 7892 23656
rect 8208 23604 8260 23656
rect 9680 23604 9732 23656
rect 5264 23536 5316 23588
rect 9588 23536 9640 23588
rect 10324 23536 10376 23588
rect 11060 23536 11112 23588
rect 11612 23536 11664 23588
rect 12348 23536 12400 23588
rect 13912 23536 13964 23588
rect 14832 23536 14884 23588
rect 15384 23536 15436 23588
rect 1768 23511 1820 23520
rect 1768 23477 1777 23511
rect 1777 23477 1811 23511
rect 1811 23477 1820 23511
rect 1768 23468 1820 23477
rect 2412 23468 2464 23520
rect 3884 23468 3936 23520
rect 4620 23468 4672 23520
rect 6828 23468 6880 23520
rect 7104 23468 7156 23520
rect 10968 23468 11020 23520
rect 11428 23468 11480 23520
rect 12808 23511 12860 23520
rect 12808 23477 12817 23511
rect 12817 23477 12851 23511
rect 12851 23477 12860 23511
rect 12808 23468 12860 23477
rect 13636 23511 13688 23520
rect 13636 23477 13645 23511
rect 13645 23477 13679 23511
rect 13679 23477 13688 23511
rect 13636 23468 13688 23477
rect 15200 23511 15252 23520
rect 15200 23477 15209 23511
rect 15209 23477 15243 23511
rect 15243 23477 15252 23511
rect 15200 23468 15252 23477
rect 16028 23468 16080 23520
rect 18236 23647 18288 23656
rect 18236 23613 18245 23647
rect 18245 23613 18279 23647
rect 18279 23613 18288 23647
rect 18236 23604 18288 23613
rect 19432 23604 19484 23656
rect 21180 23604 21232 23656
rect 24768 23647 24820 23656
rect 21640 23536 21692 23588
rect 24768 23613 24777 23647
rect 24777 23613 24811 23647
rect 24811 23613 24820 23647
rect 24768 23604 24820 23613
rect 16580 23468 16632 23520
rect 17132 23511 17184 23520
rect 17132 23477 17141 23511
rect 17141 23477 17175 23511
rect 17175 23477 17184 23511
rect 17132 23468 17184 23477
rect 19340 23468 19392 23520
rect 22284 23468 22336 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 24216 23511 24268 23520
rect 24216 23477 24225 23511
rect 24225 23477 24259 23511
rect 24259 23477 24268 23511
rect 24216 23468 24268 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2596 23264 2648 23316
rect 2780 23264 2832 23316
rect 4988 23264 5040 23316
rect 7840 23264 7892 23316
rect 3240 23196 3292 23248
rect 7748 23196 7800 23248
rect 9588 23264 9640 23316
rect 9680 23264 9732 23316
rect 10140 23307 10192 23316
rect 10140 23273 10149 23307
rect 10149 23273 10183 23307
rect 10183 23273 10192 23307
rect 10140 23264 10192 23273
rect 12440 23264 12492 23316
rect 16488 23264 16540 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 19248 23264 19300 23316
rect 21640 23264 21692 23316
rect 22376 23307 22428 23316
rect 22376 23273 22385 23307
rect 22385 23273 22419 23307
rect 22419 23273 22428 23307
rect 22376 23264 22428 23273
rect 24032 23307 24084 23316
rect 24032 23273 24041 23307
rect 24041 23273 24075 23307
rect 24075 23273 24084 23307
rect 24032 23264 24084 23273
rect 9864 23196 9916 23248
rect 11428 23196 11480 23248
rect 12256 23239 12308 23248
rect 12256 23205 12290 23239
rect 12290 23205 12308 23239
rect 12256 23196 12308 23205
rect 2320 23128 2372 23180
rect 3056 23128 3108 23180
rect 3424 23128 3476 23180
rect 4160 23128 4212 23180
rect 4620 23171 4672 23180
rect 4620 23137 4629 23171
rect 4629 23137 4663 23171
rect 4663 23137 4672 23171
rect 4620 23128 4672 23137
rect 4712 23128 4764 23180
rect 7196 23128 7248 23180
rect 11980 23171 12032 23180
rect 11980 23137 11989 23171
rect 11989 23137 12023 23171
rect 12023 23137 12032 23171
rect 11980 23128 12032 23137
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 17316 23128 17368 23180
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 18880 23171 18932 23180
rect 18880 23137 18889 23171
rect 18889 23137 18923 23171
rect 18923 23137 18932 23171
rect 18880 23128 18932 23137
rect 20812 23128 20864 23180
rect 22192 23171 22244 23180
rect 22192 23137 22201 23171
rect 22201 23137 22235 23171
rect 22235 23137 22244 23171
rect 22192 23128 22244 23137
rect 23848 23171 23900 23180
rect 23848 23137 23857 23171
rect 23857 23137 23891 23171
rect 23891 23137 23900 23171
rect 23848 23128 23900 23137
rect 1768 23060 1820 23112
rect 3056 22992 3108 23044
rect 6828 23060 6880 23112
rect 7012 23060 7064 23112
rect 9496 23060 9548 23112
rect 10968 23060 11020 23112
rect 19340 22992 19392 23044
rect 2044 22967 2096 22976
rect 2044 22933 2053 22967
rect 2053 22933 2087 22967
rect 2087 22933 2096 22967
rect 2044 22924 2096 22933
rect 3240 22924 3292 22976
rect 6276 22924 6328 22976
rect 6644 22967 6696 22976
rect 6644 22933 6653 22967
rect 6653 22933 6687 22967
rect 6687 22933 6696 22967
rect 6644 22924 6696 22933
rect 10048 22924 10100 22976
rect 10968 22924 11020 22976
rect 11152 22924 11204 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2412 22720 2464 22772
rect 3240 22720 3292 22772
rect 4160 22720 4212 22772
rect 4620 22763 4672 22772
rect 4620 22729 4629 22763
rect 4629 22729 4663 22763
rect 4663 22729 4672 22763
rect 4620 22720 4672 22729
rect 7196 22720 7248 22772
rect 8116 22720 8168 22772
rect 9680 22763 9732 22772
rect 9680 22729 9689 22763
rect 9689 22729 9723 22763
rect 9723 22729 9732 22763
rect 9680 22720 9732 22729
rect 11336 22720 11388 22772
rect 12256 22720 12308 22772
rect 16396 22720 16448 22772
rect 7012 22652 7064 22704
rect 11980 22695 12032 22704
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 6276 22584 6328 22636
rect 11980 22661 11989 22695
rect 11989 22661 12023 22695
rect 12023 22661 12032 22695
rect 11980 22652 12032 22661
rect 12348 22652 12400 22704
rect 23848 22695 23900 22704
rect 23848 22661 23857 22695
rect 23857 22661 23891 22695
rect 23891 22661 23900 22695
rect 23848 22652 23900 22661
rect 11060 22627 11112 22636
rect 4620 22516 4672 22568
rect 6552 22516 6604 22568
rect 11060 22593 11069 22627
rect 11069 22593 11103 22627
rect 11103 22593 11112 22627
rect 11060 22584 11112 22593
rect 10968 22559 11020 22568
rect 10968 22525 10977 22559
rect 10977 22525 11011 22559
rect 11011 22525 11020 22559
rect 10968 22516 11020 22525
rect 13636 22516 13688 22568
rect 15568 22516 15620 22568
rect 22560 22559 22612 22568
rect 22560 22525 22569 22559
rect 22569 22525 22603 22559
rect 22603 22525 22612 22559
rect 22560 22516 22612 22525
rect 2320 22448 2372 22500
rect 7840 22448 7892 22500
rect 8116 22448 8168 22500
rect 9772 22448 9824 22500
rect 12440 22491 12492 22500
rect 12440 22457 12449 22491
rect 12449 22457 12483 22491
rect 12483 22457 12492 22491
rect 12440 22448 12492 22457
rect 13084 22491 13136 22500
rect 13084 22457 13093 22491
rect 13093 22457 13127 22491
rect 13127 22457 13136 22491
rect 13084 22448 13136 22457
rect 14372 22448 14424 22500
rect 16212 22448 16264 22500
rect 17868 22448 17920 22500
rect 1676 22423 1728 22432
rect 1676 22389 1685 22423
rect 1685 22389 1719 22423
rect 1719 22389 1728 22423
rect 1676 22380 1728 22389
rect 2596 22380 2648 22432
rect 5448 22380 5500 22432
rect 6276 22423 6328 22432
rect 6276 22389 6285 22423
rect 6285 22389 6319 22423
rect 6319 22389 6328 22423
rect 6276 22380 6328 22389
rect 8944 22380 8996 22432
rect 10692 22380 10744 22432
rect 12348 22380 12400 22432
rect 13912 22380 13964 22432
rect 15292 22380 15344 22432
rect 15936 22380 15988 22432
rect 17316 22380 17368 22432
rect 18880 22423 18932 22432
rect 18880 22389 18889 22423
rect 18889 22389 18923 22423
rect 18923 22389 18932 22423
rect 18880 22380 18932 22389
rect 20812 22380 20864 22432
rect 22192 22423 22244 22432
rect 22192 22389 22201 22423
rect 22201 22389 22235 22423
rect 22235 22389 22244 22423
rect 22192 22380 22244 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 1768 22176 1820 22228
rect 2044 22176 2096 22228
rect 2228 22219 2280 22228
rect 2228 22185 2237 22219
rect 2237 22185 2271 22219
rect 2271 22185 2280 22219
rect 2228 22176 2280 22185
rect 2504 22176 2556 22228
rect 4712 22219 4764 22228
rect 4712 22185 4721 22219
rect 4721 22185 4755 22219
rect 4755 22185 4764 22219
rect 4712 22176 4764 22185
rect 5080 22219 5132 22228
rect 5080 22185 5089 22219
rect 5089 22185 5123 22219
rect 5123 22185 5132 22219
rect 5080 22176 5132 22185
rect 6644 22176 6696 22228
rect 7748 22219 7800 22228
rect 7748 22185 7757 22219
rect 7757 22185 7791 22219
rect 7791 22185 7800 22219
rect 7748 22176 7800 22185
rect 9772 22219 9824 22228
rect 9772 22185 9781 22219
rect 9781 22185 9815 22219
rect 9815 22185 9824 22219
rect 9772 22176 9824 22185
rect 10968 22176 11020 22228
rect 12348 22176 12400 22228
rect 12808 22176 12860 22228
rect 2688 22108 2740 22160
rect 6368 22108 6420 22160
rect 7932 22108 7984 22160
rect 8116 22108 8168 22160
rect 3056 22040 3108 22092
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 2412 22015 2464 22024
rect 2412 21981 2421 22015
rect 2421 21981 2455 22015
rect 2455 21981 2464 22015
rect 2412 21972 2464 21981
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 6000 21972 6052 22024
rect 7104 22015 7156 22024
rect 7104 21981 7113 22015
rect 7113 21981 7147 22015
rect 7147 21981 7156 22015
rect 7104 21972 7156 21981
rect 2228 21904 2280 21956
rect 8944 21972 8996 22024
rect 10140 22108 10192 22160
rect 11060 22108 11112 22160
rect 11612 22108 11664 22160
rect 10876 22040 10928 22092
rect 11704 22040 11756 22092
rect 12532 22040 12584 22092
rect 11336 22015 11388 22024
rect 11336 21981 11345 22015
rect 11345 21981 11379 22015
rect 11379 21981 11388 22015
rect 11336 21972 11388 21981
rect 13912 21972 13964 22024
rect 8024 21904 8076 21956
rect 8668 21904 8720 21956
rect 2044 21836 2096 21888
rect 3332 21879 3384 21888
rect 3332 21845 3341 21879
rect 3341 21845 3375 21879
rect 3375 21845 3384 21879
rect 3332 21836 3384 21845
rect 3608 21836 3660 21888
rect 6184 21879 6236 21888
rect 6184 21845 6193 21879
rect 6193 21845 6227 21879
rect 6227 21845 6236 21879
rect 6184 21836 6236 21845
rect 6644 21879 6696 21888
rect 6644 21845 6653 21879
rect 6653 21845 6687 21879
rect 6687 21845 6696 21879
rect 6644 21836 6696 21845
rect 8484 21836 8536 21888
rect 9588 21836 9640 21888
rect 12716 21836 12768 21888
rect 13636 21879 13688 21888
rect 13636 21845 13645 21879
rect 13645 21845 13679 21879
rect 13679 21845 13688 21879
rect 13636 21836 13688 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2136 21632 2188 21684
rect 4528 21675 4580 21684
rect 4528 21641 4537 21675
rect 4537 21641 4571 21675
rect 4571 21641 4580 21675
rect 4528 21632 4580 21641
rect 6368 21632 6420 21684
rect 6552 21675 6604 21684
rect 6552 21641 6561 21675
rect 6561 21641 6595 21675
rect 6595 21641 6604 21675
rect 6552 21632 6604 21641
rect 6736 21632 6788 21684
rect 8668 21632 8720 21684
rect 10876 21675 10928 21684
rect 10876 21641 10885 21675
rect 10885 21641 10919 21675
rect 10919 21641 10928 21675
rect 10876 21632 10928 21641
rect 11612 21675 11664 21684
rect 11612 21641 11621 21675
rect 11621 21641 11655 21675
rect 11655 21641 11664 21675
rect 11612 21632 11664 21641
rect 12348 21632 12400 21684
rect 14372 21675 14424 21684
rect 14372 21641 14381 21675
rect 14381 21641 14415 21675
rect 14415 21641 14424 21675
rect 14372 21632 14424 21641
rect 3700 21539 3752 21548
rect 3700 21505 3709 21539
rect 3709 21505 3743 21539
rect 3743 21505 3752 21539
rect 3700 21496 3752 21505
rect 3976 21496 4028 21548
rect 5080 21496 5132 21548
rect 6184 21496 6236 21548
rect 7748 21496 7800 21548
rect 4068 21428 4120 21480
rect 4896 21471 4948 21480
rect 4896 21437 4905 21471
rect 4905 21437 4939 21471
rect 4939 21437 4948 21471
rect 4896 21428 4948 21437
rect 6920 21428 6972 21480
rect 8944 21471 8996 21480
rect 8944 21437 8978 21471
rect 8978 21437 8996 21471
rect 8944 21428 8996 21437
rect 11152 21471 11204 21480
rect 11152 21437 11161 21471
rect 11161 21437 11195 21471
rect 11195 21437 11204 21471
rect 11152 21428 11204 21437
rect 2412 21403 2464 21412
rect 2412 21369 2421 21403
rect 2421 21369 2455 21403
rect 2455 21369 2464 21403
rect 2412 21360 2464 21369
rect 3884 21360 3936 21412
rect 4344 21360 4396 21412
rect 4528 21360 4580 21412
rect 5356 21403 5408 21412
rect 5356 21369 5365 21403
rect 5365 21369 5399 21403
rect 5399 21369 5408 21403
rect 5356 21360 5408 21369
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 4988 21335 5040 21344
rect 4988 21301 4997 21335
rect 4997 21301 5031 21335
rect 5031 21301 5040 21335
rect 4988 21292 5040 21301
rect 9956 21292 10008 21344
rect 11244 21292 11296 21344
rect 12440 21292 12492 21344
rect 13636 21428 13688 21480
rect 26240 21360 26292 21412
rect 27620 21360 27672 21412
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 1768 21088 1820 21140
rect 2780 21088 2832 21140
rect 5540 21088 5592 21140
rect 7104 21088 7156 21140
rect 10140 21131 10192 21140
rect 10140 21097 10149 21131
rect 10149 21097 10183 21131
rect 10183 21097 10192 21131
rect 10140 21088 10192 21097
rect 11336 21088 11388 21140
rect 13636 21088 13688 21140
rect 6000 21063 6052 21072
rect 6000 21029 6009 21063
rect 6009 21029 6043 21063
rect 6043 21029 6052 21063
rect 6000 21020 6052 21029
rect 6276 21020 6328 21072
rect 8944 21020 8996 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 4344 20995 4396 21004
rect 4344 20961 4378 20995
rect 4378 20961 4396 20995
rect 4344 20952 4396 20961
rect 10416 20952 10468 21004
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 9496 20927 9548 20936
rect 9496 20893 9505 20927
rect 9505 20893 9539 20927
rect 9539 20893 9548 20927
rect 9496 20884 9548 20893
rect 9956 20884 10008 20936
rect 11428 20927 11480 20936
rect 11428 20893 11437 20927
rect 11437 20893 11471 20927
rect 11471 20893 11480 20927
rect 11428 20884 11480 20893
rect 2688 20859 2740 20868
rect 2688 20825 2697 20859
rect 2697 20825 2731 20859
rect 2731 20825 2740 20859
rect 2688 20816 2740 20825
rect 2780 20816 2832 20868
rect 13452 20952 13504 21004
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 2228 20748 2280 20800
rect 5080 20748 5132 20800
rect 6000 20748 6052 20800
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 11336 20748 11388 20800
rect 13636 20748 13688 20800
rect 14372 20791 14424 20800
rect 14372 20757 14381 20791
rect 14381 20757 14415 20791
rect 14415 20757 14424 20791
rect 14372 20748 14424 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20544 1452 20596
rect 3424 20544 3476 20596
rect 4068 20544 4120 20596
rect 4344 20544 4396 20596
rect 6276 20587 6328 20596
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 6276 20544 6328 20553
rect 6552 20544 6604 20596
rect 8024 20544 8076 20596
rect 10140 20544 10192 20596
rect 13820 20587 13872 20596
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 1768 20408 1820 20460
rect 10416 20519 10468 20528
rect 10416 20485 10425 20519
rect 10425 20485 10459 20519
rect 10459 20485 10468 20519
rect 10416 20476 10468 20485
rect 2228 20383 2280 20392
rect 2228 20349 2262 20383
rect 2262 20349 2280 20383
rect 2228 20340 2280 20349
rect 4528 20340 4580 20392
rect 4896 20383 4948 20392
rect 4896 20349 4905 20383
rect 4905 20349 4939 20383
rect 4939 20349 4948 20383
rect 4896 20340 4948 20349
rect 3976 20272 4028 20324
rect 11244 20451 11296 20460
rect 11244 20417 11253 20451
rect 11253 20417 11287 20451
rect 11287 20417 11296 20451
rect 11244 20408 11296 20417
rect 11336 20451 11388 20460
rect 11336 20417 11345 20451
rect 11345 20417 11379 20451
rect 11379 20417 11388 20451
rect 11336 20408 11388 20417
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 13452 20408 13504 20460
rect 14372 20408 14424 20460
rect 7932 20340 7984 20392
rect 8300 20383 8352 20392
rect 1676 20204 1728 20256
rect 2320 20204 2372 20256
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 7012 20204 7064 20256
rect 8300 20349 8334 20383
rect 8334 20349 8352 20383
rect 8300 20340 8352 20349
rect 11428 20340 11480 20392
rect 13820 20340 13872 20392
rect 9588 20272 9640 20324
rect 11888 20315 11940 20324
rect 11888 20281 11897 20315
rect 11897 20281 11931 20315
rect 11931 20281 11940 20315
rect 11888 20272 11940 20281
rect 13912 20272 13964 20324
rect 9404 20247 9456 20256
rect 9404 20213 9413 20247
rect 9413 20213 9447 20247
rect 9447 20213 9456 20247
rect 9404 20204 9456 20213
rect 10968 20204 11020 20256
rect 13728 20204 13780 20256
rect 14004 20247 14056 20256
rect 14004 20213 14013 20247
rect 14013 20213 14047 20247
rect 14047 20213 14056 20247
rect 14004 20204 14056 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1768 20000 1820 20052
rect 2228 20000 2280 20052
rect 2596 20000 2648 20052
rect 3240 20000 3292 20052
rect 4528 20043 4580 20052
rect 4528 20009 4537 20043
rect 4537 20009 4571 20043
rect 4571 20009 4580 20043
rect 4528 20000 4580 20009
rect 4988 20000 5040 20052
rect 8300 20000 8352 20052
rect 9404 20000 9456 20052
rect 10048 20043 10100 20052
rect 10048 20009 10057 20043
rect 10057 20009 10091 20043
rect 10091 20009 10100 20043
rect 10048 20000 10100 20009
rect 10784 20000 10836 20052
rect 11428 20000 11480 20052
rect 13452 20043 13504 20052
rect 13452 20009 13461 20043
rect 13461 20009 13495 20043
rect 13495 20009 13504 20043
rect 13452 20000 13504 20009
rect 13912 20000 13964 20052
rect 5264 19975 5316 19984
rect 5264 19941 5273 19975
rect 5273 19941 5307 19975
rect 5307 19941 5316 19975
rect 5264 19932 5316 19941
rect 6000 19932 6052 19984
rect 8852 19932 8904 19984
rect 11244 19975 11296 19984
rect 11244 19941 11253 19975
rect 11253 19941 11287 19975
rect 11287 19941 11296 19975
rect 11244 19932 11296 19941
rect 12348 19975 12400 19984
rect 12348 19941 12360 19975
rect 12360 19941 12400 19975
rect 12348 19932 12400 19941
rect 2320 19864 2372 19916
rect 4528 19864 4580 19916
rect 6552 19864 6604 19916
rect 5080 19796 5132 19848
rect 10140 19796 10192 19848
rect 8024 19728 8076 19780
rect 3148 19660 3200 19712
rect 5172 19660 5224 19712
rect 5448 19660 5500 19712
rect 6184 19703 6236 19712
rect 6184 19669 6193 19703
rect 6193 19669 6227 19703
rect 6227 19669 6236 19703
rect 6184 19660 6236 19669
rect 9680 19703 9732 19712
rect 9680 19669 9689 19703
rect 9689 19669 9723 19703
rect 9723 19669 9732 19703
rect 9680 19660 9732 19669
rect 15384 19796 15436 19848
rect 12440 19660 12492 19712
rect 13728 19660 13780 19712
rect 14464 19703 14516 19712
rect 14464 19669 14473 19703
rect 14473 19669 14507 19703
rect 14507 19669 14516 19703
rect 14464 19660 14516 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2596 19499 2648 19508
rect 2596 19465 2605 19499
rect 2605 19465 2639 19499
rect 2639 19465 2648 19499
rect 2596 19456 2648 19465
rect 3148 19499 3200 19508
rect 3148 19465 3157 19499
rect 3157 19465 3191 19499
rect 3191 19465 3200 19499
rect 3148 19456 3200 19465
rect 12072 19456 12124 19508
rect 1952 19388 2004 19440
rect 2412 19388 2464 19440
rect 3332 19388 3384 19440
rect 3240 19320 3292 19372
rect 6184 19388 6236 19440
rect 12624 19388 12676 19440
rect 3148 19252 3200 19304
rect 3516 19295 3568 19304
rect 3516 19261 3525 19295
rect 3525 19261 3559 19295
rect 3559 19261 3568 19295
rect 4436 19320 4488 19372
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 10784 19320 10836 19372
rect 3516 19252 3568 19261
rect 4988 19252 5040 19304
rect 6184 19252 6236 19304
rect 7196 19295 7248 19304
rect 7196 19261 7205 19295
rect 7205 19261 7239 19295
rect 7239 19261 7248 19295
rect 7196 19252 7248 19261
rect 8852 19252 8904 19304
rect 9220 19295 9272 19304
rect 9220 19261 9229 19295
rect 9229 19261 9263 19295
rect 9263 19261 9272 19295
rect 9220 19252 9272 19261
rect 14464 19320 14516 19372
rect 1768 19184 1820 19236
rect 2688 19184 2740 19236
rect 6000 19184 6052 19236
rect 9404 19184 9456 19236
rect 2136 19116 2188 19168
rect 4528 19116 4580 19168
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 4988 19116 5040 19168
rect 7288 19159 7340 19168
rect 7288 19125 7297 19159
rect 7297 19125 7331 19159
rect 7331 19125 7340 19159
rect 7288 19116 7340 19125
rect 10140 19116 10192 19168
rect 10876 19116 10928 19168
rect 13360 19252 13412 19304
rect 23664 19295 23716 19304
rect 23664 19261 23673 19295
rect 23673 19261 23707 19295
rect 23707 19261 23716 19295
rect 23664 19252 23716 19261
rect 14096 19227 14148 19236
rect 14096 19193 14105 19227
rect 14105 19193 14139 19227
rect 14139 19193 14148 19227
rect 14096 19184 14148 19193
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13452 19116 13504 19125
rect 13728 19116 13780 19168
rect 14188 19159 14240 19168
rect 14188 19125 14197 19159
rect 14197 19125 14231 19159
rect 14231 19125 14240 19159
rect 14188 19116 14240 19125
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 15752 19159 15804 19168
rect 15752 19125 15761 19159
rect 15761 19125 15795 19159
rect 15795 19125 15804 19159
rect 15752 19116 15804 19125
rect 24768 19116 24820 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 1860 18912 1912 18964
rect 2504 18912 2556 18964
rect 3516 18955 3568 18964
rect 3516 18921 3525 18955
rect 3525 18921 3559 18955
rect 3559 18921 3568 18955
rect 3516 18912 3568 18921
rect 4160 18912 4212 18964
rect 5264 18912 5316 18964
rect 7564 18912 7616 18964
rect 8116 18955 8168 18964
rect 8116 18921 8125 18955
rect 8125 18921 8159 18955
rect 8159 18921 8168 18955
rect 8116 18912 8168 18921
rect 9680 18912 9732 18964
rect 10140 18955 10192 18964
rect 10140 18921 10149 18955
rect 10149 18921 10183 18955
rect 10183 18921 10192 18955
rect 10140 18912 10192 18921
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 12440 18912 12492 18964
rect 2872 18887 2924 18896
rect 2872 18853 2881 18887
rect 2881 18853 2915 18887
rect 2915 18853 2924 18887
rect 2872 18844 2924 18853
rect 3976 18844 4028 18896
rect 5448 18887 5500 18896
rect 5448 18853 5482 18887
rect 5482 18853 5500 18887
rect 5448 18844 5500 18853
rect 10232 18844 10284 18896
rect 10692 18844 10744 18896
rect 11428 18844 11480 18896
rect 12348 18844 12400 18896
rect 14096 18912 14148 18964
rect 16580 18912 16632 18964
rect 14464 18844 14516 18896
rect 15292 18844 15344 18896
rect 4344 18776 4396 18828
rect 7748 18776 7800 18828
rect 12532 18776 12584 18828
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 4620 18708 4672 18760
rect 9404 18708 9456 18760
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 3332 18640 3384 18692
rect 6828 18640 6880 18692
rect 7656 18683 7708 18692
rect 1676 18615 1728 18624
rect 1676 18581 1685 18615
rect 1685 18581 1719 18615
rect 1719 18581 1728 18615
rect 1676 18572 1728 18581
rect 3976 18572 4028 18624
rect 6920 18572 6972 18624
rect 7656 18649 7665 18683
rect 7665 18649 7699 18683
rect 7699 18649 7708 18683
rect 7656 18640 7708 18649
rect 9772 18640 9824 18692
rect 9220 18615 9272 18624
rect 9220 18581 9229 18615
rect 9229 18581 9263 18615
rect 9263 18581 9272 18615
rect 9220 18572 9272 18581
rect 13452 18708 13504 18760
rect 11888 18572 11940 18624
rect 13820 18572 13872 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 15660 18572 15712 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1676 18368 1728 18420
rect 1860 18300 1912 18352
rect 3332 18368 3384 18420
rect 5448 18368 5500 18420
rect 6092 18411 6144 18420
rect 6092 18377 6101 18411
rect 6101 18377 6135 18411
rect 6135 18377 6144 18411
rect 6092 18368 6144 18377
rect 8208 18411 8260 18420
rect 8208 18377 8217 18411
rect 8217 18377 8251 18411
rect 8251 18377 8260 18411
rect 8208 18368 8260 18377
rect 9128 18411 9180 18420
rect 9128 18377 9137 18411
rect 9137 18377 9171 18411
rect 9171 18377 9180 18411
rect 9128 18368 9180 18377
rect 10232 18411 10284 18420
rect 10232 18377 10241 18411
rect 10241 18377 10275 18411
rect 10275 18377 10284 18411
rect 10232 18368 10284 18377
rect 12532 18368 12584 18420
rect 15292 18368 15344 18420
rect 4068 18232 4120 18284
rect 5172 18275 5224 18284
rect 5172 18241 5181 18275
rect 5181 18241 5215 18275
rect 5215 18241 5224 18275
rect 5172 18232 5224 18241
rect 9404 18300 9456 18352
rect 15660 18343 15712 18352
rect 15660 18309 15669 18343
rect 15669 18309 15703 18343
rect 15703 18309 15712 18343
rect 15660 18300 15712 18309
rect 11244 18275 11296 18284
rect 11244 18241 11253 18275
rect 11253 18241 11287 18275
rect 11287 18241 11296 18275
rect 11244 18232 11296 18241
rect 11428 18275 11480 18284
rect 11428 18241 11437 18275
rect 11437 18241 11471 18275
rect 11471 18241 11480 18275
rect 11428 18232 11480 18241
rect 2872 18164 2924 18216
rect 6828 18207 6880 18216
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 9128 18164 9180 18216
rect 10324 18164 10376 18216
rect 11060 18164 11112 18216
rect 13452 18164 13504 18216
rect 6920 18096 6972 18148
rect 8300 18028 8352 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11888 18071 11940 18080
rect 11888 18037 11897 18071
rect 11897 18037 11931 18071
rect 11931 18037 11940 18071
rect 15200 18164 15252 18216
rect 14004 18139 14056 18148
rect 14004 18105 14038 18139
rect 14038 18105 14056 18139
rect 14004 18096 14056 18105
rect 11888 18028 11940 18037
rect 16396 18071 16448 18080
rect 16396 18037 16405 18071
rect 16405 18037 16439 18071
rect 16439 18037 16448 18071
rect 16396 18028 16448 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2228 17867 2280 17876
rect 2228 17833 2237 17867
rect 2237 17833 2271 17867
rect 2271 17833 2280 17867
rect 2228 17824 2280 17833
rect 4068 17824 4120 17876
rect 6092 17867 6144 17876
rect 6092 17833 6101 17867
rect 6101 17833 6135 17867
rect 6135 17833 6144 17867
rect 6092 17824 6144 17833
rect 7564 17867 7616 17876
rect 7564 17833 7573 17867
rect 7573 17833 7607 17867
rect 7607 17833 7616 17867
rect 7564 17824 7616 17833
rect 7748 17867 7800 17876
rect 7748 17833 7757 17867
rect 7757 17833 7791 17867
rect 7791 17833 7800 17867
rect 7748 17824 7800 17833
rect 10140 17824 10192 17876
rect 15108 17824 15160 17876
rect 2412 17756 2464 17808
rect 3148 17756 3200 17808
rect 4160 17756 4212 17808
rect 7932 17756 7984 17808
rect 10876 17756 10928 17808
rect 2596 17731 2648 17740
rect 2596 17697 2605 17731
rect 2605 17697 2639 17731
rect 2639 17697 2648 17731
rect 2596 17688 2648 17697
rect 4988 17731 5040 17740
rect 4988 17697 5022 17731
rect 5022 17697 5040 17731
rect 4988 17688 5040 17697
rect 8116 17731 8168 17740
rect 8116 17697 8125 17731
rect 8125 17697 8159 17731
rect 8159 17697 8168 17731
rect 8116 17688 8168 17697
rect 9864 17688 9916 17740
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 2872 17620 2924 17629
rect 4620 17620 4672 17672
rect 7472 17620 7524 17672
rect 8392 17663 8444 17672
rect 8392 17629 8401 17663
rect 8401 17629 8435 17663
rect 8435 17629 8444 17663
rect 8392 17620 8444 17629
rect 9220 17620 9272 17672
rect 10692 17620 10744 17672
rect 11888 17688 11940 17740
rect 13912 17688 13964 17740
rect 14556 17620 14608 17672
rect 16488 17688 16540 17740
rect 16856 17731 16908 17740
rect 16856 17697 16865 17731
rect 16865 17697 16899 17731
rect 16899 17697 16908 17731
rect 16856 17688 16908 17697
rect 17868 17731 17920 17740
rect 17868 17697 17877 17731
rect 17877 17697 17911 17731
rect 17911 17697 17920 17731
rect 17868 17688 17920 17697
rect 1400 17552 1452 17604
rect 3056 17552 3108 17604
rect 14004 17552 14056 17604
rect 15292 17552 15344 17604
rect 4344 17527 4396 17536
rect 4344 17493 4353 17527
rect 4353 17493 4387 17527
rect 4387 17493 4396 17527
rect 4344 17484 4396 17493
rect 4896 17484 4948 17536
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 8760 17527 8812 17536
rect 8760 17493 8769 17527
rect 8769 17493 8803 17527
rect 8803 17493 8812 17527
rect 8760 17484 8812 17493
rect 9772 17484 9824 17536
rect 11060 17484 11112 17536
rect 12072 17484 12124 17536
rect 14740 17484 14792 17536
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 17040 17527 17092 17536
rect 17040 17493 17049 17527
rect 17049 17493 17083 17527
rect 17083 17493 17092 17527
rect 17040 17484 17092 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 3148 17323 3200 17332
rect 3148 17289 3157 17323
rect 3157 17289 3191 17323
rect 3191 17289 3200 17323
rect 3148 17280 3200 17289
rect 3884 17323 3936 17332
rect 3884 17289 3893 17323
rect 3893 17289 3927 17323
rect 3927 17289 3936 17323
rect 3884 17280 3936 17289
rect 4896 17280 4948 17332
rect 7472 17323 7524 17332
rect 7472 17289 7481 17323
rect 7481 17289 7515 17323
rect 7515 17289 7524 17323
rect 7472 17280 7524 17289
rect 8024 17280 8076 17332
rect 2596 17212 2648 17264
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 4896 17187 4948 17196
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 10968 17280 11020 17332
rect 13912 17323 13964 17332
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 14832 17280 14884 17332
rect 15292 17280 15344 17332
rect 16856 17280 16908 17332
rect 8392 17212 8444 17264
rect 9128 17255 9180 17264
rect 9128 17221 9137 17255
rect 9137 17221 9171 17255
rect 9171 17221 9180 17255
rect 9128 17212 9180 17221
rect 13820 17212 13872 17264
rect 14004 17212 14056 17264
rect 14556 17255 14608 17264
rect 14556 17221 14565 17255
rect 14565 17221 14599 17255
rect 14599 17221 14608 17255
rect 14556 17212 14608 17221
rect 18236 17255 18288 17264
rect 18236 17221 18245 17255
rect 18245 17221 18279 17255
rect 18279 17221 18288 17255
rect 18236 17212 18288 17221
rect 19340 17212 19392 17264
rect 20260 17212 20312 17264
rect 4896 17144 4948 17153
rect 12808 17144 12860 17196
rect 1952 17076 2004 17128
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 7932 17076 7984 17128
rect 9496 17119 9548 17128
rect 9496 17085 9530 17119
rect 9530 17085 9548 17119
rect 9496 17076 9548 17085
rect 8024 17051 8076 17060
rect 8024 17017 8033 17051
rect 8033 17017 8067 17051
rect 8067 17017 8076 17051
rect 8024 17008 8076 17017
rect 4344 16983 4396 16992
rect 4344 16949 4353 16983
rect 4353 16949 4387 16983
rect 4387 16949 4396 16983
rect 4344 16940 4396 16949
rect 4620 16940 4672 16992
rect 10692 16940 10744 16992
rect 11704 16940 11756 16992
rect 12164 17008 12216 17060
rect 13452 17051 13504 17060
rect 13452 17017 13461 17051
rect 13461 17017 13495 17051
rect 13495 17017 13504 17051
rect 13452 17008 13504 17017
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 15844 17008 15896 17060
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1492 16736 1544 16788
rect 2504 16736 2556 16788
rect 3056 16736 3108 16788
rect 3608 16779 3660 16788
rect 3608 16745 3617 16779
rect 3617 16745 3651 16779
rect 3651 16745 3660 16779
rect 3608 16736 3660 16745
rect 3884 16736 3936 16788
rect 4988 16736 5040 16788
rect 6552 16736 6604 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 9496 16736 9548 16788
rect 7104 16668 7156 16720
rect 8116 16668 8168 16720
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 4712 16600 4764 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7472 16600 7524 16652
rect 9772 16668 9824 16720
rect 10876 16736 10928 16788
rect 12532 16736 12584 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 14740 16736 14792 16788
rect 15476 16779 15528 16788
rect 15476 16745 15485 16779
rect 15485 16745 15519 16779
rect 15519 16745 15528 16779
rect 15476 16736 15528 16745
rect 15844 16779 15896 16788
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 17960 16779 18012 16788
rect 17960 16745 17969 16779
rect 17969 16745 18003 16779
rect 18003 16745 18012 16779
rect 17960 16736 18012 16745
rect 10968 16668 11020 16720
rect 8392 16643 8444 16652
rect 8392 16609 8401 16643
rect 8401 16609 8435 16643
rect 8435 16609 8444 16643
rect 8392 16600 8444 16609
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 9864 16600 9916 16652
rect 2872 16532 2924 16584
rect 3608 16532 3660 16584
rect 6552 16532 6604 16584
rect 9496 16532 9548 16584
rect 10692 16532 10744 16584
rect 13544 16532 13596 16584
rect 14556 16643 14608 16652
rect 14556 16609 14565 16643
rect 14565 16609 14599 16643
rect 14599 16609 14608 16643
rect 14556 16600 14608 16609
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 16856 16643 16908 16652
rect 16856 16609 16890 16643
rect 16890 16609 16908 16643
rect 16856 16600 16908 16609
rect 16304 16532 16356 16584
rect 4160 16396 4212 16448
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 13452 16396 13504 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 3240 16192 3292 16244
rect 4804 16192 4856 16244
rect 6920 16235 6972 16244
rect 20 16124 72 16176
rect 6920 16201 6929 16235
rect 6929 16201 6963 16235
rect 6963 16201 6972 16235
rect 6920 16192 6972 16201
rect 7472 16192 7524 16244
rect 9496 16192 9548 16244
rect 11244 16235 11296 16244
rect 11244 16201 11253 16235
rect 11253 16201 11287 16235
rect 11287 16201 11296 16235
rect 11244 16192 11296 16201
rect 15844 16192 15896 16244
rect 16856 16192 16908 16244
rect 2136 16056 2188 16108
rect 2596 15920 2648 15972
rect 11060 16124 11112 16176
rect 15292 16124 15344 16176
rect 3608 16056 3660 16108
rect 3056 15988 3108 16040
rect 3516 16031 3568 16040
rect 3516 15997 3525 16031
rect 3525 15997 3559 16031
rect 3559 15997 3568 16031
rect 3516 15988 3568 15997
rect 7748 16056 7800 16108
rect 8392 16056 8444 16108
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 12532 16056 12584 16108
rect 16580 16056 16632 16108
rect 6460 15988 6512 16040
rect 8760 15988 8812 16040
rect 9312 15988 9364 16040
rect 11520 15988 11572 16040
rect 12808 16031 12860 16040
rect 12808 15997 12817 16031
rect 12817 15997 12851 16031
rect 12851 15997 12860 16031
rect 12808 15988 12860 15997
rect 3240 15920 3292 15972
rect 5264 15920 5316 15972
rect 9772 15920 9824 15972
rect 2872 15852 2924 15904
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 3700 15852 3752 15904
rect 4436 15852 4488 15904
rect 4712 15852 4764 15904
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6000 15852 6052 15904
rect 6920 15852 6972 15904
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12900 15895 12952 15904
rect 12440 15852 12492 15861
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 13728 15852 13780 15904
rect 14832 15988 14884 16040
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 19064 16031 19116 16040
rect 19064 15997 19073 16031
rect 19073 15997 19107 16031
rect 19107 15997 19116 16031
rect 19064 15988 19116 15997
rect 14556 15920 14608 15972
rect 16304 15852 16356 15904
rect 19248 15895 19300 15904
rect 19248 15861 19257 15895
rect 19257 15861 19291 15895
rect 19291 15861 19300 15895
rect 19248 15852 19300 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 4160 15648 4212 15700
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 9680 15648 9732 15700
rect 12532 15691 12584 15700
rect 12532 15657 12541 15691
rect 12541 15657 12575 15691
rect 12575 15657 12584 15691
rect 12532 15648 12584 15657
rect 12900 15691 12952 15700
rect 12900 15657 12909 15691
rect 12909 15657 12943 15691
rect 12943 15657 12952 15691
rect 12900 15648 12952 15657
rect 14556 15648 14608 15700
rect 15936 15648 15988 15700
rect 16856 15648 16908 15700
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 1676 15580 1728 15632
rect 1952 15580 2004 15632
rect 2780 15580 2832 15632
rect 8852 15580 8904 15632
rect 10048 15580 10100 15632
rect 11060 15580 11112 15632
rect 11980 15580 12032 15632
rect 17040 15580 17092 15632
rect 2504 15512 2556 15564
rect 5264 15512 5316 15564
rect 8392 15512 8444 15564
rect 13360 15512 13412 15564
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 16580 15555 16632 15564
rect 16580 15521 16614 15555
rect 16614 15521 16632 15555
rect 20904 15555 20956 15564
rect 16580 15512 16632 15521
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 2872 15444 2924 15496
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 6920 15444 6972 15496
rect 7104 15444 7156 15496
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 13452 15444 13504 15496
rect 14096 15444 14148 15496
rect 16304 15487 16356 15496
rect 16304 15453 16313 15487
rect 16313 15453 16347 15487
rect 16347 15453 16356 15487
rect 16304 15444 16356 15453
rect 3608 15376 3660 15428
rect 11796 15419 11848 15428
rect 11796 15385 11805 15419
rect 11805 15385 11839 15419
rect 11839 15385 11848 15419
rect 11796 15376 11848 15385
rect 12348 15376 12400 15428
rect 12900 15376 12952 15428
rect 9312 15308 9364 15360
rect 9772 15308 9824 15360
rect 11520 15308 11572 15360
rect 13820 15308 13872 15360
rect 14188 15308 14240 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1400 15104 1452 15156
rect 1676 15104 1728 15156
rect 2504 15104 2556 15156
rect 4620 15104 4672 15156
rect 6552 15104 6604 15156
rect 11060 15104 11112 15156
rect 14096 15104 14148 15156
rect 2596 15036 2648 15088
rect 4528 15036 4580 15088
rect 6184 15036 6236 15088
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 20904 15079 20956 15088
rect 20904 15045 20913 15079
rect 20913 15045 20947 15079
rect 20947 15045 20956 15079
rect 20904 15036 20956 15045
rect 9128 14968 9180 15020
rect 2320 14900 2372 14952
rect 3608 14900 3660 14952
rect 5356 14943 5408 14952
rect 5356 14909 5365 14943
rect 5365 14909 5399 14943
rect 5399 14909 5408 14943
rect 5356 14900 5408 14909
rect 3516 14832 3568 14884
rect 5080 14832 5132 14884
rect 6736 14900 6788 14952
rect 16856 14968 16908 15020
rect 2320 14807 2372 14816
rect 2320 14773 2329 14807
rect 2329 14773 2363 14807
rect 2363 14773 2372 14807
rect 2320 14764 2372 14773
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 6092 14832 6144 14884
rect 7748 14832 7800 14884
rect 10140 14832 10192 14884
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 10416 14900 10468 14952
rect 12624 14832 12676 14884
rect 13360 14875 13412 14884
rect 13360 14841 13369 14875
rect 13369 14841 13403 14875
rect 13403 14841 13412 14875
rect 13360 14832 13412 14841
rect 16304 14900 16356 14952
rect 19432 14943 19484 14952
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 14188 14875 14240 14884
rect 14188 14841 14222 14875
rect 14222 14841 14240 14875
rect 14188 14832 14240 14841
rect 17500 14832 17552 14884
rect 10784 14764 10836 14816
rect 11796 14764 11848 14816
rect 13176 14764 13228 14816
rect 13728 14807 13780 14816
rect 13728 14773 13737 14807
rect 13737 14773 13771 14807
rect 13771 14773 13780 14807
rect 13728 14764 13780 14773
rect 15292 14807 15344 14816
rect 15292 14773 15301 14807
rect 15301 14773 15335 14807
rect 15335 14773 15344 14807
rect 15292 14764 15344 14773
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2136 14560 2188 14612
rect 2504 14560 2556 14612
rect 3516 14603 3568 14612
rect 2872 14492 2924 14544
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 4528 14603 4580 14612
rect 4528 14569 4537 14603
rect 4537 14569 4571 14603
rect 4571 14569 4580 14603
rect 4528 14560 4580 14569
rect 6092 14560 6144 14612
rect 7472 14603 7524 14612
rect 7472 14569 7481 14603
rect 7481 14569 7515 14603
rect 7515 14569 7524 14603
rect 7472 14560 7524 14569
rect 8392 14603 8444 14612
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 9036 14603 9088 14612
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 10784 14603 10836 14612
rect 10784 14569 10793 14603
rect 10793 14569 10827 14603
rect 10827 14569 10836 14603
rect 10784 14560 10836 14569
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 12348 14560 12400 14612
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 13820 14560 13872 14612
rect 14464 14560 14516 14612
rect 15384 14560 15436 14612
rect 16856 14560 16908 14612
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 6552 14492 6604 14544
rect 11704 14492 11756 14544
rect 14740 14492 14792 14544
rect 16396 14535 16448 14544
rect 16396 14501 16405 14535
rect 16405 14501 16439 14535
rect 16439 14501 16448 14535
rect 16396 14492 16448 14501
rect 3884 14467 3936 14476
rect 3884 14433 3893 14467
rect 3893 14433 3927 14467
rect 3927 14433 3936 14467
rect 3884 14424 3936 14433
rect 4160 14424 4212 14476
rect 6184 14424 6236 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 11152 14424 11204 14476
rect 11428 14424 11480 14476
rect 13176 14424 13228 14476
rect 15936 14424 15988 14476
rect 3792 14356 3844 14408
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 8024 14399 8076 14408
rect 8024 14365 8033 14399
rect 8033 14365 8067 14399
rect 8067 14365 8076 14399
rect 8024 14356 8076 14365
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 3148 14288 3200 14340
rect 5080 14288 5132 14340
rect 5356 14288 5408 14340
rect 9404 14288 9456 14340
rect 10692 14356 10744 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 14188 14399 14240 14408
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 16580 14399 16632 14408
rect 14188 14356 14240 14365
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 2504 14220 2556 14272
rect 3424 14220 3476 14272
rect 3976 14220 4028 14272
rect 5264 14263 5316 14272
rect 5264 14229 5273 14263
rect 5273 14229 5307 14263
rect 5307 14229 5316 14263
rect 5264 14220 5316 14229
rect 9680 14263 9732 14272
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2320 14016 2372 14068
rect 2780 14016 2832 14068
rect 3332 14016 3384 14068
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 7196 14016 7248 14068
rect 9128 14016 9180 14068
rect 10140 14016 10192 14068
rect 11704 14016 11756 14068
rect 13176 14059 13228 14068
rect 13176 14025 13185 14059
rect 13185 14025 13219 14059
rect 13219 14025 13228 14059
rect 13176 14016 13228 14025
rect 16396 14059 16448 14068
rect 16396 14025 16405 14059
rect 16405 14025 16439 14059
rect 16439 14025 16448 14059
rect 16396 14016 16448 14025
rect 16580 14016 16632 14068
rect 3608 13948 3660 14000
rect 1860 13880 1912 13932
rect 2320 13880 2372 13932
rect 8208 13948 8260 14000
rect 6920 13880 6972 13932
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 11152 13923 11204 13932
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3608 13855 3660 13864
rect 3056 13812 3108 13821
rect 3608 13821 3617 13855
rect 3617 13821 3651 13855
rect 3651 13821 3660 13855
rect 3608 13812 3660 13821
rect 3516 13787 3568 13796
rect 3516 13753 3525 13787
rect 3525 13753 3559 13787
rect 3559 13753 3568 13787
rect 3516 13744 3568 13753
rect 5264 13744 5316 13796
rect 6736 13744 6788 13796
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 9404 13855 9456 13864
rect 9404 13821 9438 13855
rect 9438 13821 9456 13855
rect 9404 13812 9456 13821
rect 11428 13812 11480 13864
rect 13728 13855 13780 13864
rect 7196 13744 7248 13796
rect 12808 13744 12860 13796
rect 2412 13676 2464 13728
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 6552 13676 6604 13685
rect 7380 13676 7432 13728
rect 13176 13676 13228 13728
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 15936 13855 15988 13864
rect 15936 13821 15945 13855
rect 15945 13821 15979 13855
rect 15979 13821 15988 13855
rect 15936 13812 15988 13821
rect 14096 13744 14148 13796
rect 14188 13676 14240 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3516 13472 3568 13524
rect 4436 13515 4488 13524
rect 4436 13481 4445 13515
rect 4445 13481 4479 13515
rect 4479 13481 4488 13515
rect 4436 13472 4488 13481
rect 4896 13472 4948 13524
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 8116 13515 8168 13524
rect 8116 13481 8125 13515
rect 8125 13481 8159 13515
rect 8159 13481 8168 13515
rect 8116 13472 8168 13481
rect 9680 13472 9732 13524
rect 12532 13472 12584 13524
rect 14188 13472 14240 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 16580 13472 16632 13524
rect 21180 13472 21232 13524
rect 1860 13404 1912 13456
rect 2228 13404 2280 13456
rect 2412 13404 2464 13456
rect 3148 13404 3200 13456
rect 4804 13404 4856 13456
rect 6276 13447 6328 13456
rect 6276 13413 6285 13447
rect 6285 13413 6319 13447
rect 6319 13413 6328 13447
rect 6276 13404 6328 13413
rect 9404 13447 9456 13456
rect 9404 13413 9413 13447
rect 9413 13413 9447 13447
rect 9447 13413 9456 13447
rect 9404 13404 9456 13413
rect 11244 13404 11296 13456
rect 12256 13404 12308 13456
rect 4068 13336 4120 13388
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 6552 13336 6604 13388
rect 7472 13379 7524 13388
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 8300 13336 8352 13388
rect 15844 13379 15896 13388
rect 15844 13345 15878 13379
rect 15878 13345 15896 13379
rect 15844 13336 15896 13345
rect 19156 13336 19208 13388
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 9128 13268 9180 13320
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 15476 13268 15528 13320
rect 17776 13268 17828 13320
rect 5264 13200 5316 13252
rect 6000 13200 6052 13252
rect 7656 13243 7708 13252
rect 7656 13209 7665 13243
rect 7665 13209 7699 13243
rect 7699 13209 7708 13243
rect 7656 13200 7708 13209
rect 9772 13200 9824 13252
rect 19432 13243 19484 13252
rect 19432 13209 19441 13243
rect 19441 13209 19475 13243
rect 19475 13209 19484 13243
rect 19432 13200 19484 13209
rect 2228 13132 2280 13184
rect 4068 13175 4120 13184
rect 4068 13141 4077 13175
rect 4077 13141 4111 13175
rect 4111 13141 4120 13175
rect 4068 13132 4120 13141
rect 5540 13132 5592 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 14832 13132 14884 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2596 12928 2648 12980
rect 3884 12928 3936 12980
rect 4620 12928 4672 12980
rect 5264 12928 5316 12980
rect 6184 12928 6236 12980
rect 6368 12928 6420 12980
rect 8300 12928 8352 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9312 12971 9364 12980
rect 9312 12937 9321 12971
rect 9321 12937 9355 12971
rect 9355 12937 9364 12971
rect 9312 12928 9364 12937
rect 10232 12928 10284 12980
rect 11244 12971 11296 12980
rect 11244 12937 11253 12971
rect 11253 12937 11287 12971
rect 11287 12937 11296 12971
rect 11244 12928 11296 12937
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 1952 12792 2004 12844
rect 9588 12860 9640 12912
rect 4804 12792 4856 12844
rect 5356 12792 5408 12844
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 6276 12792 6328 12844
rect 8484 12792 8536 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 11336 12860 11388 12912
rect 12716 12928 12768 12980
rect 16212 12928 16264 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 22284 12928 22336 12980
rect 13820 12903 13872 12912
rect 13820 12869 13829 12903
rect 13829 12869 13863 12903
rect 13863 12869 13872 12903
rect 13820 12860 13872 12869
rect 15108 12903 15160 12912
rect 15108 12869 15117 12903
rect 15117 12869 15151 12903
rect 15151 12869 15160 12903
rect 15108 12860 15160 12869
rect 2504 12724 2556 12776
rect 5632 12724 5684 12776
rect 2964 12656 3016 12708
rect 5448 12656 5500 12708
rect 6920 12724 6972 12776
rect 9128 12724 9180 12776
rect 11336 12767 11388 12776
rect 11336 12733 11337 12767
rect 11337 12733 11371 12767
rect 11371 12733 11388 12767
rect 11336 12724 11388 12733
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 6736 12588 6788 12640
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 11796 12588 11848 12640
rect 13820 12724 13872 12776
rect 14832 12724 14884 12776
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 12532 12656 12584 12708
rect 12716 12699 12768 12708
rect 12716 12665 12728 12699
rect 12728 12665 12768 12699
rect 12716 12656 12768 12665
rect 13176 12588 13228 12640
rect 15200 12656 15252 12708
rect 15476 12656 15528 12708
rect 17776 12656 17828 12708
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 17224 12588 17276 12640
rect 19156 12588 19208 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2320 12384 2372 12436
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 4896 12384 4948 12436
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 9588 12384 9640 12436
rect 9772 12384 9824 12436
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 11704 12384 11756 12436
rect 12716 12384 12768 12436
rect 19156 12427 19208 12436
rect 19156 12393 19165 12427
rect 19165 12393 19199 12427
rect 19199 12393 19208 12427
rect 19156 12384 19208 12393
rect 22008 12427 22060 12436
rect 22008 12393 22017 12427
rect 22017 12393 22051 12427
rect 22051 12393 22060 12427
rect 22008 12384 22060 12393
rect 2780 12359 2832 12368
rect 2780 12325 2789 12359
rect 2789 12325 2823 12359
rect 2823 12325 2832 12359
rect 2780 12316 2832 12325
rect 15292 12316 15344 12368
rect 1768 12155 1820 12164
rect 1768 12121 1777 12155
rect 1777 12121 1811 12155
rect 1811 12121 1820 12155
rect 1768 12112 1820 12121
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 2688 12248 2740 12300
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 5356 12248 5408 12300
rect 6000 12248 6052 12300
rect 8300 12291 8352 12300
rect 8300 12257 8309 12291
rect 8309 12257 8343 12291
rect 8343 12257 8352 12291
rect 8300 12248 8352 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10784 12248 10836 12300
rect 11520 12248 11572 12300
rect 14004 12291 14056 12300
rect 14004 12257 14013 12291
rect 14013 12257 14047 12291
rect 14047 12257 14056 12291
rect 14004 12248 14056 12257
rect 17776 12291 17828 12300
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8668 12180 8720 12232
rect 10692 12180 10744 12232
rect 10968 12180 11020 12232
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 2228 12112 2280 12164
rect 2596 12044 2648 12096
rect 4712 12044 4764 12096
rect 5264 12044 5316 12096
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 14464 12180 14516 12232
rect 14832 12180 14884 12232
rect 15200 12180 15252 12232
rect 17776 12257 17785 12291
rect 17785 12257 17819 12291
rect 17819 12257 17828 12291
rect 17776 12248 17828 12257
rect 18052 12291 18104 12300
rect 18052 12257 18086 12291
rect 18086 12257 18104 12291
rect 18052 12248 18104 12257
rect 22008 12180 22060 12232
rect 16580 12112 16632 12164
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2320 11840 2372 11892
rect 2780 11840 2832 11892
rect 3516 11883 3568 11892
rect 3516 11849 3525 11883
rect 3525 11849 3559 11883
rect 3559 11849 3568 11883
rect 3516 11840 3568 11849
rect 5540 11840 5592 11892
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 1952 11815 2004 11824
rect 1952 11781 1961 11815
rect 1961 11781 1995 11815
rect 1995 11781 2004 11815
rect 1952 11772 2004 11781
rect 6000 11704 6052 11756
rect 8300 11840 8352 11892
rect 10784 11883 10836 11892
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 11796 11840 11848 11892
rect 15476 11840 15528 11892
rect 17224 11840 17276 11892
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 22192 11840 22244 11892
rect 16396 11704 16448 11756
rect 17132 11704 17184 11756
rect 18052 11704 18104 11756
rect 2412 11679 2464 11688
rect 2412 11645 2446 11679
rect 2446 11645 2464 11679
rect 2412 11636 2464 11645
rect 8668 11679 8720 11688
rect 2504 11568 2556 11620
rect 4068 11611 4120 11620
rect 4068 11577 4077 11611
rect 4077 11577 4111 11611
rect 4111 11577 4120 11611
rect 4068 11568 4120 11577
rect 4160 11568 4212 11620
rect 8668 11645 8702 11679
rect 8702 11645 8720 11679
rect 8668 11636 8720 11645
rect 10876 11636 10928 11688
rect 11520 11636 11572 11688
rect 13176 11679 13228 11688
rect 13176 11645 13185 11679
rect 13185 11645 13219 11679
rect 13219 11645 13228 11679
rect 13176 11636 13228 11645
rect 13452 11636 13504 11688
rect 21180 11679 21232 11688
rect 21180 11645 21189 11679
rect 21189 11645 21223 11679
rect 21223 11645 21232 11679
rect 21180 11636 21232 11645
rect 13728 11568 13780 11620
rect 17960 11568 18012 11620
rect 2780 11500 2832 11552
rect 4712 11500 4764 11552
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 7840 11500 7892 11552
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10048 11500 10100 11552
rect 11796 11543 11848 11552
rect 11796 11509 11805 11543
rect 11805 11509 11839 11543
rect 11839 11509 11848 11543
rect 11796 11500 11848 11509
rect 14004 11500 14056 11552
rect 15108 11500 15160 11552
rect 15844 11543 15896 11552
rect 15844 11509 15853 11543
rect 15853 11509 15887 11543
rect 15887 11509 15896 11543
rect 15844 11500 15896 11509
rect 17132 11543 17184 11552
rect 17132 11509 17141 11543
rect 17141 11509 17175 11543
rect 17175 11509 17184 11543
rect 17132 11500 17184 11509
rect 22008 11543 22060 11552
rect 22008 11509 22017 11543
rect 22017 11509 22051 11543
rect 22051 11509 22060 11543
rect 22008 11500 22060 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 3240 11296 3292 11348
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 5540 11296 5592 11348
rect 6092 11339 6144 11348
rect 6092 11305 6101 11339
rect 6101 11305 6135 11339
rect 6135 11305 6144 11339
rect 6092 11296 6144 11305
rect 7104 11296 7156 11348
rect 8668 11296 8720 11348
rect 11796 11296 11848 11348
rect 13452 11296 13504 11348
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 14464 11339 14516 11348
rect 14464 11305 14473 11339
rect 14473 11305 14507 11339
rect 14507 11305 14516 11339
rect 14464 11296 14516 11305
rect 14740 11296 14792 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 7380 11271 7432 11280
rect 7380 11237 7414 11271
rect 7414 11237 7432 11271
rect 7380 11228 7432 11237
rect 8208 11228 8260 11280
rect 11244 11228 11296 11280
rect 2412 11160 2464 11212
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 3976 11160 4028 11212
rect 1768 11092 1820 11144
rect 3608 11092 3660 11144
rect 4344 11092 4396 11144
rect 4068 11067 4120 11076
rect 4068 11033 4077 11067
rect 4077 11033 4111 11067
rect 4111 11033 4120 11067
rect 4068 11024 4120 11033
rect 10968 11160 11020 11212
rect 15292 11160 15344 11212
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 6276 11092 6328 11144
rect 6920 11092 6972 11144
rect 10784 11092 10836 11144
rect 12256 11092 12308 11144
rect 13084 11092 13136 11144
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 13912 11092 13964 11101
rect 13360 11067 13412 11076
rect 13360 11033 13369 11067
rect 13369 11033 13403 11067
rect 13403 11033 13412 11067
rect 13360 11024 13412 11033
rect 11980 10956 12032 11008
rect 14004 10956 14056 11008
rect 15108 11067 15160 11076
rect 15108 11033 15117 11067
rect 15117 11033 15151 11067
rect 15151 11033 15160 11067
rect 16488 11092 16540 11144
rect 15108 11024 15160 11033
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1952 10752 2004 10804
rect 2320 10752 2372 10804
rect 4344 10752 4396 10804
rect 8392 10752 8444 10804
rect 11244 10752 11296 10804
rect 13912 10752 13964 10804
rect 15568 10752 15620 10804
rect 16580 10795 16632 10804
rect 16580 10761 16589 10795
rect 16589 10761 16623 10795
rect 16623 10761 16632 10795
rect 16580 10752 16632 10761
rect 17316 10752 17368 10804
rect 19248 10752 19300 10804
rect 3884 10548 3936 10600
rect 6736 10616 6788 10668
rect 7104 10616 7156 10668
rect 7380 10659 7432 10668
rect 7380 10625 7389 10659
rect 7389 10625 7423 10659
rect 7423 10625 7432 10659
rect 7380 10616 7432 10625
rect 14004 10616 14056 10668
rect 16028 10616 16080 10668
rect 4436 10591 4488 10600
rect 4436 10557 4459 10591
rect 4459 10557 4488 10591
rect 4436 10548 4488 10557
rect 6644 10548 6696 10600
rect 6920 10548 6972 10600
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 9496 10591 9548 10600
rect 7840 10548 7892 10557
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 9680 10591 9732 10600
rect 9680 10557 9689 10591
rect 9689 10557 9723 10591
rect 9723 10557 9732 10591
rect 9680 10548 9732 10557
rect 10784 10548 10836 10600
rect 13176 10548 13228 10600
rect 16764 10591 16816 10600
rect 16764 10557 16773 10591
rect 16773 10557 16807 10591
rect 16807 10557 16816 10591
rect 16764 10548 16816 10557
rect 18236 10548 18288 10600
rect 1952 10523 2004 10532
rect 1952 10489 1986 10523
rect 1986 10489 2004 10523
rect 1952 10480 2004 10489
rect 9772 10480 9824 10532
rect 10140 10480 10192 10532
rect 11980 10480 12032 10532
rect 15108 10480 15160 10532
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 14832 10412 14884 10464
rect 15292 10412 15344 10464
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 17592 10455 17644 10464
rect 17592 10421 17601 10455
rect 17601 10421 17635 10455
rect 17635 10421 17644 10455
rect 17592 10412 17644 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3148 10208 3200 10260
rect 4436 10208 4488 10260
rect 7380 10208 7432 10260
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 7840 10208 7892 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 10876 10208 10928 10260
rect 12256 10208 12308 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 17132 10251 17184 10260
rect 17132 10217 17141 10251
rect 17141 10217 17175 10251
rect 17175 10217 17184 10251
rect 17132 10208 17184 10217
rect 1768 10183 1820 10192
rect 1768 10149 1777 10183
rect 1777 10149 1811 10183
rect 1811 10149 1820 10183
rect 1768 10140 1820 10149
rect 3240 10140 3292 10192
rect 3516 10183 3568 10192
rect 3516 10149 3525 10183
rect 3525 10149 3559 10183
rect 3559 10149 3568 10183
rect 3516 10140 3568 10149
rect 4344 10140 4396 10192
rect 5356 10140 5408 10192
rect 8208 10140 8260 10192
rect 8852 10140 8904 10192
rect 11704 10183 11756 10192
rect 11704 10149 11713 10183
rect 11713 10149 11747 10183
rect 11747 10149 11756 10183
rect 11704 10140 11756 10149
rect 13728 10140 13780 10192
rect 14004 10183 14056 10192
rect 14004 10149 14013 10183
rect 14013 10149 14047 10183
rect 14047 10149 14056 10183
rect 14004 10140 14056 10149
rect 16028 10183 16080 10192
rect 16028 10149 16062 10183
rect 16062 10149 16080 10183
rect 16028 10140 16080 10149
rect 2964 10115 3016 10124
rect 2964 10081 2973 10115
rect 2973 10081 3007 10115
rect 3007 10081 3016 10115
rect 2964 10072 3016 10081
rect 3424 10072 3476 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 9680 10072 9732 10124
rect 11244 10072 11296 10124
rect 11520 10072 11572 10124
rect 13820 10072 13872 10124
rect 15476 10072 15528 10124
rect 15752 10115 15804 10124
rect 15752 10081 15761 10115
rect 15761 10081 15795 10115
rect 15795 10081 15804 10115
rect 15752 10072 15804 10081
rect 1952 10047 2004 10056
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 3148 10004 3200 10056
rect 4160 10004 4212 10056
rect 5172 10047 5224 10056
rect 5172 10013 5181 10047
rect 5181 10013 5215 10047
rect 5215 10013 5224 10047
rect 5172 10004 5224 10013
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 9404 10004 9456 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 11980 10004 12032 10056
rect 2228 9936 2280 9988
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 5080 9868 5132 9920
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 12808 9868 12860 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1860 9664 1912 9716
rect 3608 9664 3660 9716
rect 3884 9707 3936 9716
rect 3884 9673 3893 9707
rect 3893 9673 3927 9707
rect 3927 9673 3936 9707
rect 3884 9664 3936 9673
rect 4712 9664 4764 9716
rect 5172 9664 5224 9716
rect 5356 9707 5408 9716
rect 5356 9673 5365 9707
rect 5365 9673 5399 9707
rect 5399 9673 5408 9707
rect 5356 9664 5408 9673
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 10324 9664 10376 9716
rect 11704 9664 11756 9716
rect 14004 9707 14056 9716
rect 14004 9673 14013 9707
rect 14013 9673 14047 9707
rect 14047 9673 14056 9707
rect 14004 9664 14056 9673
rect 16028 9664 16080 9716
rect 17592 9664 17644 9716
rect 18236 9707 18288 9716
rect 18236 9673 18245 9707
rect 18245 9673 18279 9707
rect 18279 9673 18288 9707
rect 18236 9664 18288 9673
rect 1492 9596 1544 9648
rect 1768 9596 1820 9648
rect 2412 9596 2464 9648
rect 9680 9639 9732 9648
rect 9680 9605 9689 9639
rect 9689 9605 9723 9639
rect 9723 9605 9732 9639
rect 9680 9596 9732 9605
rect 11152 9596 11204 9648
rect 12348 9596 12400 9648
rect 12808 9596 12860 9648
rect 2320 9460 2372 9512
rect 3884 9460 3936 9512
rect 4620 9460 4672 9512
rect 5448 9460 5500 9512
rect 10692 9528 10744 9580
rect 15752 9596 15804 9648
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 7932 9460 7984 9512
rect 12900 9460 12952 9512
rect 7012 9392 7064 9444
rect 12716 9392 12768 9444
rect 14556 9460 14608 9512
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 15752 9392 15804 9444
rect 4252 9324 4304 9376
rect 8484 9324 8536 9376
rect 9404 9324 9456 9376
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 10140 9367 10192 9376
rect 9496 9324 9548 9333
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11520 9324 11572 9376
rect 12440 9367 12492 9376
rect 12440 9333 12449 9367
rect 12449 9333 12483 9367
rect 12483 9333 12492 9367
rect 12440 9324 12492 9333
rect 12992 9324 13044 9376
rect 13452 9324 13504 9376
rect 13820 9324 13872 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1860 9163 1912 9172
rect 1860 9129 1869 9163
rect 1869 9129 1903 9163
rect 1903 9129 1912 9163
rect 1860 9120 1912 9129
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 2596 9163 2648 9172
rect 2596 9129 2605 9163
rect 2605 9129 2639 9163
rect 2639 9129 2648 9163
rect 2596 9120 2648 9129
rect 2688 9120 2740 9172
rect 3976 9120 4028 9172
rect 4160 9120 4212 9172
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 5356 9120 5408 9172
rect 6920 9120 6972 9172
rect 8024 9120 8076 9172
rect 2964 9095 3016 9104
rect 2964 9061 2973 9095
rect 2973 9061 3007 9095
rect 3007 9061 3016 9095
rect 2964 9052 3016 9061
rect 6368 9095 6420 9104
rect 6368 9061 6377 9095
rect 6377 9061 6411 9095
rect 6411 9061 6420 9095
rect 6368 9052 6420 9061
rect 6736 9052 6788 9104
rect 7472 9052 7524 9104
rect 8484 9095 8536 9104
rect 8484 9061 8493 9095
rect 8493 9061 8527 9095
rect 8527 9061 8536 9095
rect 8484 9052 8536 9061
rect 10140 9120 10192 9172
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 12992 9120 13044 9172
rect 15568 9120 15620 9172
rect 16028 9120 16080 9172
rect 16672 9120 16724 9172
rect 1952 8984 2004 9036
rect 2136 8984 2188 9036
rect 7748 8984 7800 9036
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 7012 8959 7064 8968
rect 6552 8916 6604 8925
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 2504 8848 2556 8900
rect 7840 8848 7892 8900
rect 9956 9027 10008 9036
rect 9956 8993 9990 9027
rect 9990 8993 10008 9027
rect 9956 8984 10008 8993
rect 12440 8984 12492 9036
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 12808 8984 12860 9036
rect 16396 9027 16448 9036
rect 16396 8993 16405 9027
rect 16405 8993 16439 9027
rect 16439 8993 16448 9027
rect 16396 8984 16448 8993
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 14556 8848 14608 8900
rect 10692 8780 10744 8832
rect 11612 8823 11664 8832
rect 11612 8789 11621 8823
rect 11621 8789 11655 8823
rect 11655 8789 11664 8823
rect 11612 8780 11664 8789
rect 12900 8780 12952 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 2136 8576 2188 8628
rect 4160 8576 4212 8628
rect 4620 8576 4672 8628
rect 6552 8576 6604 8628
rect 7472 8619 7524 8628
rect 7472 8585 7481 8619
rect 7481 8585 7515 8619
rect 7515 8585 7524 8619
rect 7472 8576 7524 8585
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 10784 8576 10836 8585
rect 12808 8576 12860 8628
rect 16396 8619 16448 8628
rect 16396 8585 16405 8619
rect 16405 8585 16439 8619
rect 16439 8585 16448 8619
rect 16396 8576 16448 8585
rect 1676 8551 1728 8560
rect 1676 8517 1685 8551
rect 1685 8517 1719 8551
rect 1719 8517 1728 8551
rect 1676 8508 1728 8517
rect 6368 8508 6420 8560
rect 6736 8508 6788 8560
rect 9956 8508 10008 8560
rect 4528 8440 4580 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 11704 8508 11756 8560
rect 11612 8440 11664 8492
rect 2044 8372 2096 8424
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8208 8415 8260 8424
rect 8208 8381 8242 8415
rect 8242 8381 8260 8415
rect 8208 8372 8260 8381
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 10600 8347 10652 8356
rect 10600 8313 10609 8347
rect 10609 8313 10643 8347
rect 10643 8313 10652 8347
rect 10600 8304 10652 8313
rect 9680 8236 9732 8288
rect 10140 8236 10192 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1952 8032 2004 8084
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 11612 8032 11664 8084
rect 12440 8032 12492 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 10140 7964 10192 8016
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 10692 7939 10744 7948
rect 10692 7905 10726 7939
rect 10726 7905 10744 7939
rect 10692 7896 10744 7905
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 10416 7531 10468 7540
rect 10416 7497 10425 7531
rect 10425 7497 10459 7531
rect 10459 7497 10468 7531
rect 10416 7488 10468 7497
rect 10692 7488 10744 7540
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 4804 6400 4856 6452
rect 9496 6400 9548 6452
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 10968 5856 11020 5908
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9956 5763 10008 5772
rect 9680 5720 9732 5729
rect 9956 5729 9990 5763
rect 9990 5729 10008 5763
rect 9956 5720 10008 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 9680 5312 9732 5364
rect 9956 4972 10008 5024
rect 13912 4972 13964 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3146 27520 3202 28000
rect 3698 27520 3754 28000
rect 3790 27704 3846 27713
rect 3790 27639 3846 27648
rect 308 24834 336 27520
rect 32 24806 336 24834
rect 32 16182 60 24806
rect 20 16176 72 16182
rect 20 16118 72 16124
rect 860 14793 888 27520
rect 1306 23624 1362 23633
rect 1306 23559 1362 23568
rect 1320 23066 1348 23559
rect 1412 23202 1440 27520
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 23225 1624 25094
rect 1872 24886 1900 25298
rect 1860 24880 1912 24886
rect 1860 24822 1912 24828
rect 1676 24744 1728 24750
rect 1676 24686 1728 24692
rect 1688 24070 1716 24686
rect 1768 24608 1820 24614
rect 1820 24568 1900 24596
rect 1768 24550 1820 24556
rect 1676 24064 1728 24070
rect 1676 24006 1728 24012
rect 1688 23361 1716 24006
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1674 23352 1730 23361
rect 1674 23287 1730 23296
rect 1582 23216 1638 23225
rect 1412 23174 1532 23202
rect 1320 23038 1440 23066
rect 1412 21010 1440 23038
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 20602 1440 20946
rect 1400 20596 1452 20602
rect 1400 20538 1452 20544
rect 1504 19802 1532 23174
rect 1582 23151 1638 23160
rect 1780 23118 1808 23462
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 1596 21690 1624 22471
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 1688 22114 1716 22374
rect 1780 22234 1808 23054
rect 1768 22228 1820 22234
rect 1768 22170 1820 22176
rect 1688 22086 1808 22114
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1582 21448 1638 21457
rect 1582 21383 1638 21392
rect 1596 21146 1624 21383
rect 1780 21146 1808 22086
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1780 20466 1808 21082
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1676 20256 1728 20262
rect 1676 20198 1728 20204
rect 1412 19774 1532 19802
rect 1412 17610 1440 19774
rect 1582 19680 1638 19689
rect 1582 19615 1638 19624
rect 1490 19136 1546 19145
rect 1490 19071 1546 19080
rect 1400 17604 1452 17610
rect 1400 17546 1452 17552
rect 1398 17504 1454 17513
rect 1398 17439 1454 17448
rect 1412 15162 1440 17439
rect 1504 16794 1532 19071
rect 1596 17338 1624 19615
rect 1688 18850 1716 20198
rect 1780 20058 1808 20402
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1768 19236 1820 19242
rect 1768 19178 1820 19184
rect 1780 18970 1808 19178
rect 1872 19122 1900 24568
rect 1964 19446 1992 27520
rect 2320 25356 2372 25362
rect 2320 25298 2372 25304
rect 2332 24886 2360 25298
rect 2320 24880 2372 24886
rect 2318 24848 2320 24857
rect 2372 24848 2374 24857
rect 2318 24783 2374 24792
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 24410 2452 24550
rect 2412 24404 2464 24410
rect 2412 24346 2464 24352
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 2134 23080 2190 23089
rect 2134 23015 2190 23024
rect 2044 22976 2096 22982
rect 2044 22918 2096 22924
rect 2056 22234 2084 22918
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 2044 21888 2096 21894
rect 2044 21830 2096 21836
rect 1952 19440 2004 19446
rect 1952 19382 2004 19388
rect 1872 19094 1992 19122
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 1688 18822 1808 18850
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 18426 1716 18566
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1582 17096 1638 17105
rect 1582 17031 1638 17040
rect 1492 16788 1544 16794
rect 1492 16730 1544 16736
rect 1596 16250 1624 17031
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1688 15638 1716 18362
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 1688 15162 1716 15574
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 846 14784 902 14793
rect 846 14719 902 14728
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1504 9654 1532 14583
rect 1780 14113 1808 18822
rect 1872 18358 1900 18906
rect 1860 18352 1912 18358
rect 1860 18294 1912 18300
rect 1964 17134 1992 19094
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1952 15632 2004 15638
rect 1952 15574 2004 15580
rect 1858 14784 1914 14793
rect 1858 14719 1914 14728
rect 1766 14104 1822 14113
rect 1766 14039 1822 14048
rect 1872 13938 1900 14719
rect 1964 14618 1992 15574
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 13462 1900 13874
rect 1964 13870 1992 14554
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12345 1624 12582
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1766 12200 1822 12209
rect 1766 12135 1768 12144
rect 1820 12135 1822 12144
rect 1768 12106 1820 12112
rect 1964 11830 1992 12786
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 1964 11354 1992 11766
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10198 1808 11086
rect 1964 10810 1992 11290
rect 1952 10804 2004 10810
rect 1952 10746 2004 10752
rect 1858 10568 1914 10577
rect 1858 10503 1914 10512
rect 1952 10532 2004 10538
rect 1872 10266 1900 10503
rect 1952 10474 2004 10480
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 1780 9654 1808 10134
rect 1872 9722 1900 10202
rect 1964 10062 1992 10474
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1768 9648 1820 9654
rect 1964 9602 1992 9998
rect 1768 9590 1820 9596
rect 1872 9574 1992 9602
rect 1872 9178 1900 9574
rect 2056 9330 2084 21830
rect 2148 21690 2176 23015
rect 2240 22234 2268 24006
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2424 23526 2452 23598
rect 2412 23520 2464 23526
rect 2412 23462 2464 23468
rect 2320 23180 2372 23186
rect 2320 23122 2372 23128
rect 2332 22506 2360 23122
rect 2424 22778 2452 23462
rect 2412 22772 2464 22778
rect 2412 22714 2464 22720
rect 2320 22500 2372 22506
rect 2320 22442 2372 22448
rect 2516 22386 2544 27520
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2792 24750 2820 26551
rect 3054 25392 3110 25401
rect 3054 25327 3056 25336
rect 3108 25327 3110 25336
rect 3056 25298 3108 25304
rect 2964 25220 3016 25226
rect 2964 25162 3016 25168
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 2608 24256 2636 24346
rect 2608 24228 2820 24256
rect 2688 24132 2740 24138
rect 2688 24074 2740 24080
rect 2700 23594 2728 24074
rect 2688 23588 2740 23594
rect 2688 23530 2740 23536
rect 2792 23322 2820 24228
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2608 23225 2636 23258
rect 2594 23216 2650 23225
rect 2594 23151 2650 23160
rect 2778 23216 2834 23225
rect 2778 23151 2834 23160
rect 2608 22438 2636 23151
rect 2792 22953 2820 23151
rect 2778 22944 2834 22953
rect 2778 22879 2834 22888
rect 2332 22358 2544 22386
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2228 22228 2280 22234
rect 2228 22170 2280 22176
rect 2240 21962 2268 22170
rect 2228 21956 2280 21962
rect 2228 21898 2280 21904
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2228 20800 2280 20806
rect 2228 20742 2280 20748
rect 2240 20398 2268 20742
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2240 20058 2268 20334
rect 2332 20262 2360 22358
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2424 21418 2452 21966
rect 2412 21412 2464 21418
rect 2412 21354 2464 21360
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2148 16674 2176 19110
rect 2228 18760 2280 18766
rect 2332 18748 2360 19858
rect 2412 19440 2464 19446
rect 2412 19382 2464 19388
rect 2424 18850 2452 19382
rect 2516 18970 2544 22170
rect 2688 22160 2740 22166
rect 2740 22108 2820 22114
rect 2688 22102 2820 22108
rect 2700 22086 2820 22102
rect 2792 21146 2820 22086
rect 2884 22001 2912 25094
rect 2976 24818 3004 25162
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2976 23304 3004 24754
rect 3068 24682 3096 25298
rect 3056 24676 3108 24682
rect 3056 24618 3108 24624
rect 3068 24449 3096 24618
rect 3054 24440 3110 24449
rect 3054 24375 3110 24384
rect 2976 23276 3096 23304
rect 2962 23216 3018 23225
rect 3068 23186 3096 23276
rect 2962 23151 3018 23160
rect 3056 23180 3108 23186
rect 2870 21992 2926 22001
rect 2870 21927 2926 21936
rect 2780 21140 2832 21146
rect 2780 21082 2832 21088
rect 2686 20904 2742 20913
rect 2686 20839 2688 20848
rect 2740 20839 2742 20848
rect 2780 20868 2832 20874
rect 2688 20810 2740 20816
rect 2780 20810 2832 20816
rect 2792 20754 2820 20810
rect 2700 20726 2820 20754
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2608 19514 2636 19994
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2700 19242 2728 20726
rect 2976 20369 3004 23151
rect 3056 23122 3108 23128
rect 3056 23044 3108 23050
rect 3056 22986 3108 22992
rect 3068 22098 3096 22986
rect 3056 22092 3108 22098
rect 3056 22034 3108 22040
rect 3160 21298 3188 27520
rect 3332 25424 3384 25430
rect 3332 25366 3384 25372
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3252 24342 3280 24686
rect 3240 24336 3292 24342
rect 3240 24278 3292 24284
rect 3252 24177 3280 24278
rect 3238 24168 3294 24177
rect 3238 24103 3294 24112
rect 3344 23882 3372 25366
rect 3712 24834 3740 27520
rect 3528 24806 3740 24834
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 3436 24313 3464 24686
rect 3422 24304 3478 24313
rect 3422 24239 3478 24248
rect 3252 23854 3372 23882
rect 3252 23254 3280 23854
rect 3330 23760 3386 23769
rect 3330 23695 3386 23704
rect 3240 23248 3292 23254
rect 3240 23190 3292 23196
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 3252 22778 3280 22918
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3344 21894 3372 23695
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3068 21270 3188 21298
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 2962 20360 3018 20369
rect 2962 20295 3018 20304
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2872 18896 2924 18902
rect 2424 18822 2636 18850
rect 2872 18838 2924 18844
rect 2412 18760 2464 18766
rect 2332 18720 2412 18748
rect 2228 18702 2280 18708
rect 2412 18702 2464 18708
rect 2240 17882 2268 18702
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2424 17814 2452 18702
rect 2608 18680 2636 18822
rect 2608 18652 2820 18680
rect 2686 18592 2742 18601
rect 2686 18527 2742 18536
rect 2502 18048 2558 18057
rect 2502 17983 2558 17992
rect 2412 17808 2464 17814
rect 2412 17750 2464 17756
rect 2516 16794 2544 17983
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2608 17513 2636 17682
rect 2594 17504 2650 17513
rect 2594 17439 2650 17448
rect 2608 17270 2636 17439
rect 2700 17338 2728 18527
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2148 16646 2268 16674
rect 2134 16552 2190 16561
rect 2134 16487 2190 16496
rect 2148 16114 2176 16487
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2148 14618 2176 16050
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2240 14498 2268 16646
rect 2596 15972 2648 15978
rect 2596 15914 2648 15920
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2516 15162 2544 15506
rect 2608 15178 2636 15914
rect 2792 15638 2820 18652
rect 2884 18222 2912 18838
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2884 17678 2912 18158
rect 3068 17898 3096 21270
rect 3146 21176 3202 21185
rect 3146 21111 3202 21120
rect 3160 21010 3188 21111
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3252 20058 3280 21286
rect 3436 20602 3464 23122
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19514 3188 19654
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3160 19310 3188 19450
rect 3252 19378 3280 19994
rect 3332 19440 3384 19446
rect 3528 19394 3556 24806
rect 3698 24712 3754 24721
rect 3698 24647 3754 24656
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3620 21350 3648 21830
rect 3712 21554 3740 24647
rect 3804 22953 3832 27639
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 4158 27160 4214 27169
rect 4158 27095 4214 27104
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 4066 24576 4122 24585
rect 3988 24410 4016 24550
rect 4066 24511 4122 24520
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3790 22944 3846 22953
rect 3790 22879 3846 22888
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3896 21418 3924 23462
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3884 21412 3936 21418
rect 3884 21354 3936 21360
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3620 20505 3648 21286
rect 3606 20496 3662 20505
rect 3606 20431 3662 20440
rect 3988 20330 4016 21490
rect 4080 21486 4108 24511
rect 4172 23866 4200 27095
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4160 23656 4212 23662
rect 4160 23598 4212 23604
rect 4172 23186 4200 23598
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 4172 22778 4200 23122
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 4172 21026 4200 22714
rect 4080 21010 4200 21026
rect 4068 21004 4200 21010
rect 4120 20998 4200 21004
rect 4068 20946 4120 20952
rect 4080 20602 4108 20946
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 3332 19382 3384 19388
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3344 18698 3372 19382
rect 3436 19366 3556 19394
rect 3332 18692 3384 18698
rect 3332 18634 3384 18640
rect 3344 18426 3372 18634
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3068 17870 3280 17898
rect 3148 17808 3200 17814
rect 3148 17750 3200 17756
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2884 16590 2912 17614
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2962 17504 3018 17513
rect 2962 17439 3018 17448
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2872 15904 2924 15910
rect 2976 15892 3004 17439
rect 3068 16794 3096 17546
rect 3160 17338 3188 17750
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3068 16046 3096 16730
rect 3252 16250 3280 17870
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 3148 15904 3200 15910
rect 2976 15864 3096 15892
rect 2872 15846 2924 15852
rect 2884 15706 2912 15846
rect 2872 15700 2924 15706
rect 2924 15660 3004 15688
rect 2872 15642 2924 15648
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2504 15156 2556 15162
rect 2608 15150 2820 15178
rect 2504 15098 2556 15104
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2332 14822 2360 14894
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 1964 9302 2084 9330
rect 2148 14470 2268 14498
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1964 9042 1992 9302
rect 2042 9208 2098 9217
rect 2042 9143 2098 9152
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1676 8560 1728 8566
rect 1674 8528 1676 8537
rect 1728 8528 1730 8537
rect 1674 8463 1730 8472
rect 1964 8090 1992 8978
rect 2056 8634 2084 9143
rect 2148 9042 2176 14470
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 13462 2268 14214
rect 2332 14074 2360 14758
rect 2516 14618 2544 15098
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2516 14278 2544 14554
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12306 2268 13126
rect 2332 12442 2360 13874
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2424 13462 2452 13670
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2608 12986 2636 15030
rect 2792 14657 2820 15150
rect 2884 15026 2912 15438
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2778 14648 2834 14657
rect 2778 14583 2834 14592
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 14074 2820 14418
rect 2884 14249 2912 14486
rect 2870 14240 2926 14249
rect 2870 14175 2926 14184
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2516 12594 2544 12718
rect 2516 12566 2636 12594
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2332 12322 2360 12378
rect 2228 12300 2280 12306
rect 2332 12294 2452 12322
rect 2228 12242 2280 12248
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2240 9994 2268 12106
rect 2332 11898 2360 12174
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2332 10810 2360 11834
rect 2424 11694 2452 12294
rect 2608 12102 2636 12566
rect 2700 12458 2728 13262
rect 2976 12714 3004 15660
rect 3068 14226 3096 15864
rect 3148 15846 3200 15852
rect 3160 14346 3188 15846
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3068 14198 3188 14226
rect 3054 14104 3110 14113
rect 3054 14039 3110 14048
rect 3068 13870 3096 14039
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3160 13682 3188 14198
rect 3068 13654 3188 13682
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2700 12430 2820 12458
rect 2792 12374 2820 12430
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2424 11218 2452 11630
rect 2504 11620 2556 11626
rect 2504 11562 2556 11568
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2410 11112 2466 11121
rect 2410 11047 2466 11056
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2424 9654 2452 11047
rect 2412 9648 2464 9654
rect 2318 9616 2374 9625
rect 2412 9590 2464 9596
rect 2318 9551 2374 9560
rect 2332 9518 2360 9551
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 9178 2360 9454
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2148 8634 2176 8978
rect 2516 8906 2544 11562
rect 2608 9178 2636 12038
rect 2700 9178 2728 12242
rect 2792 11898 2820 12310
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 11218 2820 11494
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10266 2820 11154
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2976 9110 3004 10066
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2504 8900 2556 8906
rect 2504 8842 2556 8848
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2056 8430 2084 8570
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 3068 2802 3096 13654
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3160 10266 3188 13398
rect 3252 12617 3280 15914
rect 3436 15688 3464 19366
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18970 3556 19246
rect 3516 18964 3568 18970
rect 3516 18906 3568 18912
rect 3988 18902 4016 20266
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 3976 18896 4028 18902
rect 3976 18838 4028 18844
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3606 18048 3662 18057
rect 3606 17983 3662 17992
rect 3620 16794 3648 17983
rect 3882 17912 3938 17921
rect 3882 17847 3938 17856
rect 3896 17338 3924 17847
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3620 16114 3648 16526
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3344 15660 3464 15688
rect 3344 14498 3372 15660
rect 3528 15473 3556 15982
rect 3514 15464 3570 15473
rect 3620 15434 3648 16050
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3514 15399 3570 15408
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3514 15056 3570 15065
rect 3514 14991 3570 15000
rect 3528 14890 3556 14991
rect 3620 14958 3648 15370
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3528 14618 3556 14826
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3344 14470 3556 14498
rect 3330 14376 3386 14385
rect 3330 14311 3386 14320
rect 3344 14074 3372 14311
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3238 12608 3294 12617
rect 3238 12543 3294 12552
rect 3252 11354 3280 12543
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3252 10198 3280 11290
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3436 10130 3464 14214
rect 3528 13802 3556 14470
rect 3620 14006 3648 14894
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3608 13864 3660 13870
rect 3606 13832 3608 13841
rect 3660 13832 3662 13841
rect 3516 13796 3568 13802
rect 3606 13767 3662 13776
rect 3516 13738 3568 13744
rect 3528 13569 3556 13738
rect 3514 13560 3570 13569
rect 3514 13495 3516 13504
rect 3568 13495 3570 13504
rect 3516 13466 3568 13472
rect 3528 13435 3556 13466
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3528 10198 3556 11834
rect 3608 11144 3660 11150
rect 3712 11121 3740 15846
rect 3896 14929 3924 16730
rect 3988 15201 4016 18566
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4080 17882 4108 18226
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4172 17814 4200 18906
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4264 17082 4292 27520
rect 4526 26072 4582 26081
rect 4526 26007 4582 26016
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4448 24313 4476 24550
rect 4434 24304 4490 24313
rect 4434 24239 4490 24248
rect 4540 21690 4568 26007
rect 4816 25514 4844 27520
rect 4632 25486 4844 25514
rect 4632 24721 4660 25486
rect 4712 25356 4764 25362
rect 4712 25298 4764 25304
rect 4724 24818 4752 25298
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4618 24712 4674 24721
rect 4618 24647 4674 24656
rect 4816 24342 4844 25230
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4632 23526 4660 24142
rect 4712 24064 4764 24070
rect 4712 24006 4764 24012
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 4632 23186 4660 23462
rect 4724 23186 4752 24006
rect 4816 23866 4844 24278
rect 5000 24070 5028 25230
rect 5368 24886 5396 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5356 24880 5408 24886
rect 5356 24822 5408 24828
rect 5540 24608 5592 24614
rect 5540 24550 5592 24556
rect 5080 24268 5132 24274
rect 5080 24210 5132 24216
rect 4988 24064 5040 24070
rect 4988 24006 5040 24012
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 5092 23730 5120 24210
rect 5446 23760 5502 23769
rect 5080 23724 5132 23730
rect 5446 23695 5502 23704
rect 5080 23666 5132 23672
rect 5092 23474 5120 23666
rect 5460 23662 5488 23695
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5000 23446 5120 23474
rect 5000 23322 5028 23446
rect 5078 23352 5134 23361
rect 4988 23316 5040 23322
rect 5078 23287 5134 23296
rect 4988 23258 5040 23264
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4618 22944 4674 22953
rect 4618 22879 4674 22888
rect 4632 22778 4660 22879
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4632 22574 4660 22714
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4724 22234 4752 23122
rect 5092 22234 5120 23287
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 5080 22228 5132 22234
rect 5080 22170 5132 22176
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4540 21418 4568 21626
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4344 21412 4396 21418
rect 4344 21354 4396 21360
rect 4528 21412 4580 21418
rect 4528 21354 4580 21360
rect 4356 21010 4384 21354
rect 4344 21004 4396 21010
rect 4344 20946 4396 20952
rect 4356 20602 4384 20946
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4540 20398 4568 21354
rect 4908 20398 4936 21422
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4528 20392 4580 20398
rect 4896 20392 4948 20398
rect 4528 20334 4580 20340
rect 4894 20360 4896 20369
rect 4948 20360 4950 20369
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4448 19378 4476 20198
rect 4540 20058 4568 20334
rect 4894 20295 4950 20304
rect 5000 20058 5028 21286
rect 5092 20806 5120 21490
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4540 19174 4568 19858
rect 5000 19310 5028 19994
rect 5092 19854 5120 20742
rect 5276 19990 5304 23530
rect 5552 23225 5580 24550
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5538 23216 5594 23225
rect 5538 23151 5594 23160
rect 6012 23089 6040 27520
rect 6564 24857 6592 27520
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6550 24848 6606 24857
rect 6550 24783 6606 24792
rect 6184 24744 6236 24750
rect 6182 24712 6184 24721
rect 6236 24712 6238 24721
rect 6182 24647 6238 24656
rect 6458 23896 6514 23905
rect 6458 23831 6460 23840
rect 6512 23831 6514 23840
rect 6460 23802 6512 23808
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6840 23118 6868 23462
rect 6828 23112 6880 23118
rect 5998 23080 6054 23089
rect 6828 23054 6880 23060
rect 5998 23015 6054 23024
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5630 22672 5686 22681
rect 6288 22642 6316 22918
rect 5630 22607 5632 22616
rect 5684 22607 5686 22616
rect 6276 22636 6328 22642
rect 5632 22578 5684 22584
rect 6276 22578 6328 22584
rect 6288 22438 6316 22578
rect 6552 22568 6604 22574
rect 6366 22536 6422 22545
rect 6552 22510 6604 22516
rect 6366 22471 6422 22480
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 5460 22114 5488 22374
rect 5460 22086 5580 22114
rect 5552 22030 5580 22086
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 5354 21448 5410 21457
rect 5354 21383 5356 21392
rect 5408 21383 5410 21392
rect 5356 21354 5408 21360
rect 5552 21146 5580 21966
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 6012 21078 6040 21966
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 21554 6224 21830
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 6288 21078 6316 22374
rect 6380 22166 6408 22471
rect 6368 22160 6420 22166
rect 6368 22102 6420 22108
rect 6380 21690 6408 22102
rect 6564 21690 6592 22510
rect 6656 22234 6684 22918
rect 6644 22228 6696 22234
rect 6696 22188 6776 22216
rect 6644 22170 6696 22176
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6000 21072 6052 21078
rect 6000 21014 6052 21020
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6012 20806 6040 21014
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 19990 6040 20742
rect 6288 20602 6316 21014
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6564 20602 6592 20878
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 6000 19984 6052 19990
rect 6000 19926 6052 19932
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5092 19417 5120 19790
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5078 19408 5134 19417
rect 5078 19343 5134 19352
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4988 19168 5040 19174
rect 5092 19122 5120 19343
rect 5040 19116 5120 19122
rect 4988 19110 5120 19116
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4356 17542 4384 18770
rect 4344 17536 4396 17542
rect 4540 17513 4568 19110
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4632 17678 4660 18702
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4344 17478 4396 17484
rect 4526 17504 4582 17513
rect 4356 17241 4384 17478
rect 4526 17439 4582 17448
rect 4342 17232 4398 17241
rect 4342 17167 4398 17176
rect 4264 17054 4568 17082
rect 4344 16992 4396 16998
rect 4158 16960 4214 16969
rect 4344 16934 4396 16940
rect 4158 16895 4214 16904
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 4080 15745 4108 16623
rect 4172 16454 4200 16895
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4066 15736 4122 15745
rect 4172 15706 4200 16390
rect 4066 15671 4122 15680
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4066 15600 4122 15609
rect 4066 15535 4122 15544
rect 3974 15192 4030 15201
rect 3974 15127 4030 15136
rect 3882 14920 3938 14929
rect 3882 14855 3938 14864
rect 4080 14770 4108 15535
rect 3988 14742 4108 14770
rect 3882 14512 3938 14521
rect 3882 14447 3884 14456
rect 3936 14447 3938 14456
rect 3884 14418 3936 14424
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 11354 3832 14350
rect 3988 14278 4016 14742
rect 4066 14648 4122 14657
rect 4066 14583 4068 14592
rect 4120 14583 4122 14592
rect 4068 14554 4120 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 3976 14272 4028 14278
rect 4172 14249 4200 14418
rect 3976 14214 4028 14220
rect 4158 14240 4214 14249
rect 4158 14175 4214 14184
rect 4172 14074 4200 14175
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 13190 4108 13330
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3896 12442 3924 12922
rect 4080 12753 4108 13126
rect 4250 12880 4306 12889
rect 4250 12815 4306 12824
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4264 12442 4292 12815
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4080 11626 4108 12242
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3608 11086 3660 11092
rect 3698 11112 3754 11121
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3148 10056 3200 10062
rect 3528 10010 3556 10134
rect 3200 10004 3556 10010
rect 3148 9998 3556 10004
rect 3160 9982 3556 9998
rect 3620 9722 3648 11086
rect 3698 11047 3754 11056
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3790 10432 3846 10441
rect 3790 10367 3846 10376
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3804 4865 3832 10367
rect 3896 9722 3924 10542
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3896 9518 3924 9658
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3988 9178 4016 11154
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4080 10713 4108 11018
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 4172 10554 4200 11562
rect 4356 11234 4384 16934
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4448 15910 4476 16594
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4540 15745 4568 17054
rect 4632 16998 4660 17614
rect 4724 17134 4752 18022
rect 4816 17202 4844 19110
rect 5000 19094 5120 19110
rect 5000 17746 5028 19094
rect 5184 18290 5212 19654
rect 5276 18970 5304 19926
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5460 19378 5488 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5460 18902 5488 19314
rect 6012 19242 6040 19926
rect 6564 19922 6592 20538
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 19446 6224 19654
rect 6184 19440 6236 19446
rect 6184 19382 6236 19388
rect 6196 19310 6224 19382
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6000 19236 6052 19242
rect 6000 19178 6052 19184
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 5460 18426 5488 18838
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5092 17785 5120 18022
rect 6104 17882 6132 18362
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 5078 17776 5134 17785
rect 4988 17740 5040 17746
rect 5078 17711 5134 17720
rect 4988 17682 5040 17688
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 17338 4936 17478
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4908 17202 4936 17274
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4526 15736 4582 15745
rect 4448 15694 4526 15722
rect 4448 13530 4476 15694
rect 4526 15671 4582 15680
rect 4540 15611 4568 15671
rect 4632 15502 4660 16934
rect 5000 16794 5028 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4724 15910 4752 16594
rect 6564 16590 6592 16730
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6460 16448 6512 16454
rect 6458 16416 6460 16425
rect 6512 16416 6514 16425
rect 5622 16348 5918 16368
rect 6458 16351 6514 16360
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4620 15496 4672 15502
rect 4540 15456 4620 15484
rect 4540 15094 4568 15456
rect 4620 15438 4672 15444
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4526 14920 4582 14929
rect 4526 14855 4582 14864
rect 4540 14618 4568 14855
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4632 14414 4660 15098
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 14074 4660 14350
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4632 12986 4660 13262
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12102 4752 15846
rect 4816 13462 4844 16186
rect 6472 16046 6500 16351
rect 6460 16040 6512 16046
rect 5170 16008 5226 16017
rect 6460 15982 6512 15988
rect 5170 15943 5226 15952
rect 5264 15972 5316 15978
rect 5184 15910 5212 15943
rect 5264 15914 5316 15920
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5276 15570 5304 15914
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5092 14793 5120 14826
rect 5276 14822 5304 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5264 14816 5316 14822
rect 5078 14784 5134 14793
rect 5078 14719 5134 14728
rect 5262 14784 5264 14793
rect 5316 14784 5318 14793
rect 5262 14719 5318 14728
rect 5368 14346 5396 14894
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4816 12850 4844 13398
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4908 12442 4936 13466
rect 4988 12640 5040 12646
rect 4986 12608 4988 12617
rect 5040 12608 5042 12617
rect 4986 12543 5042 12552
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11558 4752 12038
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4080 10526 4200 10554
rect 4264 11206 4384 11234
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4080 9058 4108 10526
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9178 4200 9998
rect 4264 9382 4292 11206
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10810 4384 11086
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4356 10198 4384 10746
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10266 4476 10542
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4526 10024 4582 10033
rect 4526 9959 4582 9968
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4540 9178 4568 9959
rect 5092 9926 5120 14282
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 13920 5304 14214
rect 5552 13977 5580 14758
rect 6012 14521 6040 15846
rect 6564 15162 6592 16526
rect 6656 15609 6684 21830
rect 6748 21690 6776 22188
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6932 21486 6960 25230
rect 7012 24268 7064 24274
rect 7012 24210 7064 24216
rect 7024 24177 7052 24210
rect 7010 24168 7066 24177
rect 7010 24103 7066 24112
rect 7024 23866 7052 24103
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7116 23633 7144 27520
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7576 23662 7604 24074
rect 7564 23656 7616 23662
rect 7102 23624 7158 23633
rect 7564 23598 7616 23604
rect 7102 23559 7158 23568
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 7024 22710 7052 23054
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 7116 22030 7144 23462
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7208 22778 7236 23122
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 7116 21146 7144 21966
rect 7668 21185 7696 27520
rect 8220 25106 8248 27520
rect 8128 25078 8248 25106
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8128 24721 8156 25078
rect 8206 24848 8262 24857
rect 8404 24818 8432 25094
rect 8206 24783 8208 24792
rect 8260 24783 8262 24792
rect 8392 24812 8444 24818
rect 8208 24754 8260 24760
rect 8392 24754 8444 24760
rect 8114 24712 8170 24721
rect 8114 24647 8170 24656
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7760 23730 7788 24006
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7760 23254 7788 23666
rect 7852 23662 7880 24550
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7852 23322 7880 23598
rect 7840 23316 7892 23322
rect 7840 23258 7892 23264
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 7760 22488 7788 23190
rect 7840 22500 7892 22506
rect 7760 22460 7840 22488
rect 7760 22234 7788 22460
rect 7840 22442 7892 22448
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7760 21554 7788 22170
rect 7944 22166 7972 24550
rect 8022 24440 8078 24449
rect 8022 24375 8024 24384
rect 8076 24375 8078 24384
rect 8024 24346 8076 24352
rect 8036 23798 8064 24346
rect 8404 24206 8432 24754
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8024 23792 8076 23798
rect 8024 23734 8076 23740
rect 8220 23662 8248 24142
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 8116 22772 8168 22778
rect 8220 22760 8248 23598
rect 8168 22732 8248 22760
rect 8116 22714 8168 22720
rect 8116 22500 8168 22506
rect 8036 22460 8116 22488
rect 7932 22160 7984 22166
rect 7932 22102 7984 22108
rect 8036 21962 8064 22460
rect 8116 22442 8168 22448
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7654 21176 7710 21185
rect 7104 21140 7156 21146
rect 7654 21111 7710 21120
rect 7104 21082 7156 21088
rect 7654 21040 7710 21049
rect 7654 20975 7710 20984
rect 7194 20496 7250 20505
rect 7194 20431 7250 20440
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6840 18222 6868 18634
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6932 18154 6960 18566
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17542 6960 18090
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6840 16658 6960 16674
rect 6828 16652 6960 16658
rect 6880 16646 6960 16652
rect 6828 16594 6880 16600
rect 6932 16250 6960 16646
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6932 15745 6960 15846
rect 6918 15736 6974 15745
rect 6918 15671 6920 15680
rect 6972 15671 6974 15680
rect 6920 15642 6972 15648
rect 6642 15600 6698 15609
rect 6642 15535 6698 15544
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6104 14618 6132 14826
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5998 14512 6054 14521
rect 6196 14482 6224 15030
rect 6564 14550 6592 15098
rect 6736 14952 6788 14958
rect 6932 14940 6960 15438
rect 6788 14912 6960 14940
rect 6736 14894 6788 14900
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 5998 14447 6054 14456
rect 6184 14476 6236 14482
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5538 13968 5594 13977
rect 5276 13892 5396 13920
rect 5538 13903 5594 13912
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13433 5212 13670
rect 5170 13424 5226 13433
rect 5170 13359 5226 13368
rect 5276 13258 5304 13738
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5276 12986 5304 13194
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5368 12850 5396 13892
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5552 13190 5580 13670
rect 6012 13258 6040 14447
rect 6184 14418 6236 14424
rect 6196 14074 6224 14418
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 6196 13138 6224 14010
rect 6274 13832 6330 13841
rect 6274 13767 6330 13776
rect 6288 13462 6316 13767
rect 6564 13734 6592 14486
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6564 13394 6592 13670
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5276 12102 5304 12543
rect 5368 12306 5396 12786
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5460 12238 5488 12650
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5552 11898 5580 13126
rect 6196 13110 6316 13138
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5814 12880 5870 12889
rect 5814 12815 5816 12824
rect 5868 12815 5870 12824
rect 5816 12786 5868 12792
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 6090 12744 6146 12753
rect 5644 12617 5672 12718
rect 6090 12679 6146 12688
rect 5630 12608 5686 12617
rect 5630 12543 5686 12552
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 6012 11762 6040 12242
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11354 5580 11494
rect 6104 11354 6132 12679
rect 6196 11801 6224 12922
rect 6288 12850 6316 13110
rect 6380 12986 6408 13262
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6288 11898 6316 12786
rect 6748 12646 6776 13738
rect 6932 13530 6960 13874
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6932 12782 6960 13466
rect 6920 12776 6972 12782
rect 6840 12736 6920 12764
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6840 12442 6868 12736
rect 6920 12718 6972 12724
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6182 11792 6238 11801
rect 6182 11727 6238 11736
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6288 11150 6316 11834
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 5540 10464 5592 10470
rect 6552 10464 6604 10470
rect 5540 10406 5592 10412
rect 6550 10432 6552 10441
rect 6604 10432 6606 10441
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5184 9722 5212 9998
rect 5368 9722 5396 10134
rect 5552 9738 5580 10406
rect 6550 10367 6606 10376
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5460 9710 5580 9738
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 3988 9030 4108 9058
rect 3882 6760 3938 6769
rect 3882 6695 3938 6704
rect 3790 4856 3846 4865
rect 3790 4791 3846 4800
rect 3896 3777 3924 6695
rect 3988 5409 4016 9030
rect 4172 8634 4200 9114
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4540 8498 4568 9114
rect 4632 8974 4660 9454
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8634 4660 8910
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4080 7177 4108 7919
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 3974 5400 4030 5409
rect 3974 5335 4030 5344
rect 4080 4321 4108 6831
rect 4724 4842 4752 9658
rect 5368 9178 5396 9658
rect 5460 9518 5488 9710
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 6366 9480 6422 9489
rect 6366 9415 6422 9424
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 6380 9110 6408 9415
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6380 8566 6408 9046
rect 6564 8974 6592 9862
rect 6656 9518 6684 10542
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6748 9110 6776 10610
rect 6932 10606 6960 11086
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 7024 9625 7052 20198
rect 7208 19310 7236 20431
rect 7378 19408 7434 19417
rect 7378 19343 7380 19352
rect 7432 19343 7434 19352
rect 7380 19314 7432 19320
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7300 18873 7328 19110
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7286 18864 7342 18873
rect 7286 18799 7342 18808
rect 7576 17882 7604 18906
rect 7668 18698 7696 20975
rect 8036 20602 8064 21898
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 7932 20392 7984 20398
rect 7984 20340 8064 20346
rect 7932 20334 8064 20340
rect 7944 20318 8064 20334
rect 7930 19816 7986 19825
rect 8036 19786 8064 20318
rect 8128 20097 8156 22102
rect 8114 20088 8170 20097
rect 8114 20023 8170 20032
rect 7930 19751 7986 19760
rect 8024 19780 8076 19786
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7760 17882 7788 18770
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7944 17814 7972 19751
rect 8024 19722 8076 19728
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7484 17678 7512 17709
rect 7472 17672 7524 17678
rect 7470 17640 7472 17649
rect 7524 17640 7526 17649
rect 7470 17575 7526 17584
rect 7484 17338 7512 17575
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7116 15706 7144 16662
rect 7484 16658 7512 17274
rect 7944 17134 7972 17750
rect 8036 17338 8064 19722
rect 8114 19272 8170 19281
rect 8114 19207 8170 19216
rect 8128 18970 8156 19207
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8220 18426 8248 22732
rect 8680 21962 8708 23666
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8298 20632 8354 20641
rect 8298 20567 8354 20576
rect 8312 20398 8340 20567
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8312 20058 8340 20334
rect 8300 20052 8352 20058
rect 8352 20012 8432 20040
rect 8300 19994 8352 20000
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8300 18080 8352 18086
rect 8298 18048 8300 18057
rect 8352 18048 8354 18057
rect 8298 17983 8354 17992
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8128 17649 8156 17682
rect 8404 17678 8432 20012
rect 8496 17921 8524 21830
rect 8680 21690 8708 21898
rect 8668 21684 8720 21690
rect 8668 21626 8720 21632
rect 8864 19990 8892 27520
rect 9128 25220 9180 25226
rect 9128 25162 9180 25168
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8956 22030 8984 22374
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8956 21486 8984 21966
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8956 21078 8984 21422
rect 8944 21072 8996 21078
rect 8944 21014 8996 21020
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8864 19310 8892 19926
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 9140 18426 9168 25162
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 9324 24614 9352 24686
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9324 23730 9352 24550
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 9416 20777 9444 27520
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9508 23118 9536 24618
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9600 23866 9628 24210
rect 9692 23905 9720 24550
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9678 23896 9734 23905
rect 9588 23860 9640 23866
rect 9784 23866 9812 24346
rect 9678 23831 9734 23840
rect 9772 23860 9824 23866
rect 9588 23802 9640 23808
rect 9772 23802 9824 23808
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9600 23322 9628 23530
rect 9692 23322 9720 23598
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9508 22098 9536 23054
rect 9692 22778 9720 23258
rect 9876 23254 9904 23666
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9968 22681 9996 27520
rect 10520 25786 10548 27520
rect 10520 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10140 24064 10192 24070
rect 10140 24006 10192 24012
rect 10152 23322 10180 24006
rect 10336 23594 10364 24142
rect 10704 23769 10732 25758
rect 10968 24404 11020 24410
rect 11072 24392 11100 27520
rect 11020 24364 11100 24392
rect 10968 24346 11020 24352
rect 11612 24336 11664 24342
rect 11612 24278 11664 24284
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 10690 23760 10746 23769
rect 10690 23695 10746 23704
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 9954 22672 10010 22681
rect 9954 22607 10010 22616
rect 9772 22500 9824 22506
rect 9772 22442 9824 22448
rect 9784 22234 9812 22442
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 10060 22137 10088 22918
rect 10152 22166 10180 23258
rect 10980 23118 11008 23462
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 10980 22574 11008 22918
rect 11072 22642 11100 23530
rect 11440 23526 11468 24142
rect 11624 23594 11652 24278
rect 11612 23588 11664 23594
rect 11612 23530 11664 23536
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11440 23254 11468 23462
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22160 10192 22166
rect 10046 22128 10102 22137
rect 9496 22092 9548 22098
rect 10140 22102 10192 22108
rect 10046 22063 10102 22072
rect 9496 22034 9548 22040
rect 9588 21888 9640 21894
rect 9640 21848 9812 21876
rect 9588 21830 9640 21836
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9402 20768 9458 20777
rect 9402 20703 9458 20712
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 20058 9444 20198
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9232 18630 9260 19246
rect 9416 19242 9444 19994
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9416 18766 9444 19178
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9140 18222 9168 18362
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 8482 17912 8538 17921
rect 8482 17847 8538 17856
rect 9232 17678 9260 18566
rect 9416 18358 9444 18702
rect 9404 18352 9456 18358
rect 9404 18294 9456 18300
rect 8392 17672 8444 17678
rect 8114 17640 8170 17649
rect 9220 17672 9272 17678
rect 8392 17614 8444 17620
rect 9140 17632 9220 17660
rect 8114 17575 8170 17584
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 8036 16794 8064 17002
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8128 16726 8156 17575
rect 8404 17270 8432 17614
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 7484 16250 7512 16594
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 8404 16114 8432 16594
rect 8772 16561 8800 17478
rect 9140 17270 9168 17632
rect 9220 17614 9272 17620
rect 9232 17549 9260 17614
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9508 17134 9536 20878
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9600 19451 9628 20266
rect 9692 19825 9720 20742
rect 9678 19816 9734 19825
rect 9678 19751 9734 19760
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9586 19442 9642 19451
rect 9586 19377 9642 19386
rect 9692 18970 9720 19654
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9784 18698 9812 21848
rect 10138 21584 10194 21593
rect 10138 21519 10194 21528
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 20942 9996 21286
rect 10152 21146 10180 21519
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 10152 20602 10180 21082
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10428 20534 10456 20946
rect 10416 20528 10468 20534
rect 10414 20496 10416 20505
rect 10468 20496 10470 20505
rect 10414 20431 10470 20440
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10046 20088 10102 20097
rect 10289 20080 10585 20100
rect 10046 20023 10048 20032
rect 10100 20023 10102 20032
rect 10048 19994 10100 20000
rect 10704 19938 10732 22374
rect 10980 22234 11008 22510
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11072 22166 11100 22578
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 10888 21690 10916 22034
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 11164 21486 11192 22918
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11348 22030 11376 22714
rect 11612 22160 11664 22166
rect 11612 22102 11664 22108
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11164 21049 11192 21422
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11150 21040 11206 21049
rect 11150 20975 11206 20984
rect 11256 20618 11284 21286
rect 11348 21146 11376 21966
rect 11624 21690 11652 22102
rect 11716 22098 11744 27520
rect 12268 24818 12296 27520
rect 12820 27418 12848 27520
rect 12820 27390 12940 27418
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 11794 24712 11850 24721
rect 11794 24647 11796 24656
rect 11848 24647 11850 24656
rect 11796 24618 11848 24624
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12254 23352 12310 23361
rect 12254 23287 12310 23296
rect 12360 23304 12388 23530
rect 12440 23316 12492 23322
rect 12268 23254 12296 23287
rect 12360 23276 12440 23304
rect 12440 23258 12492 23264
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 11992 22710 12020 23122
rect 12268 22778 12296 23190
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 12360 22438 12388 22646
rect 12438 22536 12494 22545
rect 12438 22471 12440 22480
rect 12492 22471 12494 22480
rect 12440 22442 12492 22448
rect 12348 22432 12400 22438
rect 12400 22380 12480 22386
rect 12348 22374 12480 22380
rect 12360 22358 12480 22374
rect 12360 22309 12388 22358
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 12360 21690 12388 22170
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 11624 21457 11652 21626
rect 11610 21448 11666 21457
rect 11610 21383 11666 21392
rect 12452 21350 12480 22358
rect 12544 22098 12572 24550
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12820 22234 12848 23462
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 12452 20942 12480 21286
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11164 20590 11284 20618
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 9968 19910 10732 19938
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9678 17232 9734 17241
rect 9678 17167 9734 17176
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9508 16794 9536 17070
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9508 16590 9536 16730
rect 9692 16658 9720 17167
rect 9784 16833 9812 17478
rect 9770 16824 9826 16833
rect 9770 16759 9826 16768
rect 9772 16720 9824 16726
rect 9770 16688 9772 16697
rect 9824 16688 9826 16697
rect 9680 16652 9732 16658
rect 9876 16658 9904 17682
rect 9770 16623 9826 16632
rect 9864 16652 9916 16658
rect 9680 16594 9732 16600
rect 9864 16594 9916 16600
rect 9496 16584 9548 16590
rect 8758 16552 8814 16561
rect 9496 16526 9548 16532
rect 8758 16487 8814 16496
rect 8482 16416 8538 16425
rect 8482 16351 8538 16360
rect 8758 16416 8814 16425
rect 8758 16351 8814 16360
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7194 15464 7250 15473
rect 7116 11354 7144 15438
rect 7194 15399 7250 15408
rect 7208 14074 7236 15399
rect 7300 15337 7328 15846
rect 7760 15502 7788 16050
rect 8404 15570 8432 16050
rect 8496 15706 8524 16351
rect 8772 16046 8800 16351
rect 9508 16250 9536 16526
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 7748 15496 7800 15502
rect 7746 15464 7748 15473
rect 7800 15464 7802 15473
rect 7746 15399 7802 15408
rect 7286 15328 7342 15337
rect 7286 15263 7342 15272
rect 7760 14890 7788 15399
rect 8390 14920 8446 14929
rect 7748 14884 7800 14890
rect 8390 14855 8446 14864
rect 7748 14826 7800 14832
rect 7470 14784 7526 14793
rect 7470 14719 7526 14728
rect 7484 14618 7512 14719
rect 8404 14618 8432 14855
rect 8864 14822 8892 15574
rect 9324 15366 9352 15982
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9508 15609 9536 15846
rect 9692 15706 9720 16594
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9494 15600 9550 15609
rect 9494 15535 9550 15544
rect 9784 15366 9812 15914
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8024 14408 8076 14414
rect 8022 14376 8024 14385
rect 8576 14408 8628 14414
rect 8076 14376 8078 14385
rect 8576 14350 8628 14356
rect 8022 14311 8078 14320
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7208 13802 7236 14010
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7392 11370 7420 13670
rect 8128 13530 8156 13874
rect 8116 13524 8168 13530
rect 8116 13466 8168 13472
rect 8220 13410 8248 13942
rect 8588 13841 8616 14350
rect 8574 13832 8630 13841
rect 8574 13767 8630 13776
rect 8220 13394 8340 13410
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 8220 13388 8352 13394
rect 8220 13382 8300 13388
rect 7484 12102 7512 13330
rect 7654 13288 7710 13297
rect 7654 13223 7656 13232
rect 7708 13223 7710 13232
rect 7656 13194 7708 13200
rect 8220 13002 8248 13382
rect 8300 13330 8352 13336
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8220 12986 8340 13002
rect 8220 12980 8352 12986
rect 8220 12974 8300 12980
rect 8300 12922 8352 12928
rect 8496 12850 8524 13126
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7484 11665 7512 12038
rect 7944 11665 7972 12038
rect 7470 11656 7526 11665
rect 7470 11591 7526 11600
rect 7930 11656 7986 11665
rect 7930 11591 7986 11600
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7104 11348 7156 11354
rect 7392 11342 7512 11370
rect 7104 11290 7156 11296
rect 7116 10674 7144 11290
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7392 10674 7420 11222
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7392 10266 7420 10610
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7010 9616 7066 9625
rect 7010 9551 7066 9560
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8634 6592 8910
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6748 8566 6776 9046
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6932 8498 6960 9114
rect 7024 8974 7052 9386
rect 7484 9110 7512 11342
rect 7852 10606 7880 11494
rect 8220 11286 8248 12582
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8312 11898 8340 12242
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8404 10810 8432 12174
rect 8680 11694 8708 12174
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11354 8708 11630
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7668 10169 7696 10202
rect 7654 10160 7710 10169
rect 7654 10095 7710 10104
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7484 8634 7512 9046
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7760 8945 7788 8978
rect 7746 8936 7802 8945
rect 7852 8906 7880 10202
rect 8128 10146 8156 10202
rect 8864 10198 8892 14758
rect 9034 14648 9090 14657
rect 9034 14583 9036 14592
rect 9088 14583 9090 14592
rect 9036 14554 9088 14560
rect 9140 14074 9168 14962
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9140 13870 9168 14010
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9140 12986 9168 13262
rect 9324 12986 9352 15302
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9416 13870 9444 14282
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9402 13560 9458 13569
rect 9692 13530 9720 14214
rect 9402 13495 9458 13504
rect 9680 13524 9732 13530
rect 9416 13462 9444 13495
rect 9680 13466 9732 13472
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9784 13258 9812 15302
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9140 12782 9168 12922
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9600 12442 9628 12854
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9784 12442 9812 12786
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9496 10600 9548 10606
rect 9680 10600 9732 10606
rect 9548 10560 9680 10588
rect 9496 10542 9548 10548
rect 9680 10542 9732 10548
rect 9784 10538 9812 11494
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 8208 10192 8260 10198
rect 8128 10140 8208 10146
rect 8128 10134 8260 10140
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8024 10124 8076 10130
rect 8128 10118 8239 10134
rect 9680 10124 9732 10130
rect 8024 10066 8076 10072
rect 9680 10066 9732 10072
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7746 8871 7802 8880
rect 7840 8900 7892 8906
rect 7760 8634 7788 8871
rect 7840 8842 7892 8848
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7944 8430 7972 9454
rect 8036 9178 8064 10066
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 9404 10056 9456 10062
rect 9692 10010 9720 10066
rect 9404 9998 9456 10004
rect 8220 9722 8248 9998
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8220 8430 8248 9658
rect 9416 9382 9444 9998
rect 9600 9982 9720 10010
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9496 9376 9548 9382
rect 9600 9364 9628 9982
rect 9680 9648 9732 9654
rect 9678 9616 9680 9625
rect 9732 9616 9734 9625
rect 9678 9551 9734 9560
rect 9548 9336 9628 9364
rect 9496 9318 9548 9324
rect 8496 9110 8524 9318
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8208 8424 8260 8430
rect 8260 8372 8340 8378
rect 8208 8366 8340 8372
rect 7944 8090 7972 8366
rect 8220 8350 8340 8366
rect 8220 8301 8248 8350
rect 8312 8090 8340 8350
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 9508 6905 9536 9318
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8294 9720 8910
rect 9876 8537 9904 16594
rect 9968 9217 9996 19910
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10152 19174 10180 19790
rect 10796 19378 10824 19994
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10690 19000 10746 19009
rect 10140 18964 10192 18970
rect 10690 18935 10746 18944
rect 10140 18906 10192 18912
rect 10152 17882 10180 18906
rect 10704 18902 10732 18935
rect 10232 18896 10284 18902
rect 10232 18838 10284 18844
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10244 18426 10272 18838
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10336 18222 10364 18702
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10704 16998 10732 17614
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16590 10732 16934
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10060 15638 10088 16050
rect 10704 16028 10732 16526
rect 10796 16153 10824 18022
rect 10888 17814 10916 19110
rect 10980 17921 11008 20198
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10966 17912 11022 17921
rect 10966 17847 11022 17856
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10888 16794 10916 17750
rect 11072 17542 11100 18158
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10980 16726 11008 17274
rect 10968 16720 11020 16726
rect 11164 16697 11192 20590
rect 11348 20466 11376 20742
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11256 19990 11284 20402
rect 11440 20398 11468 20878
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11886 20360 11942 20369
rect 11440 20058 11468 20334
rect 11886 20295 11888 20304
rect 11940 20295 11942 20304
rect 11888 20266 11940 20272
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 12348 19984 12400 19990
rect 12348 19926 12400 19932
rect 12070 19680 12126 19689
rect 12070 19615 12126 19624
rect 12084 19514 12112 19615
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11256 18290 11284 18906
rect 12360 18902 12388 19926
rect 12452 19718 12480 20878
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12530 19680 12586 19689
rect 12530 19615 12586 19624
rect 12544 19530 12572 19615
rect 12452 19502 12572 19530
rect 12452 18970 12480 19502
rect 12624 19440 12676 19446
rect 12544 19400 12624 19428
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 11440 18290 11468 18838
rect 12544 18834 12572 19400
rect 12624 19382 12676 19388
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11900 18086 11928 18566
rect 12544 18426 12572 18770
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17746 11928 18022
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11150 16688 11206 16697
rect 11020 16668 11100 16674
rect 10968 16662 11100 16668
rect 10980 16646 11100 16662
rect 11072 16182 11100 16646
rect 11150 16623 11206 16632
rect 11242 16280 11298 16289
rect 11242 16215 11244 16224
rect 11296 16215 11298 16224
rect 11244 16186 11296 16192
rect 11060 16176 11112 16182
rect 10782 16144 10838 16153
rect 11060 16118 11112 16124
rect 10782 16079 10838 16088
rect 11520 16040 11572 16046
rect 10704 16000 10824 16028
rect 10796 15910 10824 16000
rect 11520 15982 11572 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14958 10456 15438
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 14385 10088 14418
rect 10046 14376 10102 14385
rect 10046 14311 10102 14320
rect 10060 13569 10088 14311
rect 10152 14074 10180 14826
rect 10796 14822 10824 15846
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 11072 15162 11100 15574
rect 11532 15366 11560 15982
rect 11520 15360 11572 15366
rect 11716 15337 11744 16934
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11794 15464 11850 15473
rect 11794 15399 11796 15408
rect 11848 15399 11850 15408
rect 11796 15370 11848 15376
rect 11520 15302 11572 15308
rect 11702 15328 11758 15337
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10796 14618 10824 14758
rect 11072 14618 11100 15098
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10046 13560 10102 13569
rect 10046 13495 10102 13504
rect 10152 13308 10180 14010
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10232 13320 10284 13326
rect 10152 13280 10232 13308
rect 10232 13262 10284 13268
rect 10244 12986 10272 13262
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11558 10088 12242
rect 10704 12238 10732 14350
rect 11164 13977 11192 14418
rect 11150 13968 11206 13977
rect 11150 13903 11152 13912
rect 11204 13903 11206 13912
rect 11152 13874 11204 13880
rect 11440 13870 11468 14418
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11244 13456 11296 13462
rect 11244 13398 11296 13404
rect 11256 12986 11284 13398
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11348 12782 11376 12854
rect 11336 12776 11388 12782
rect 10782 12744 10838 12753
rect 11336 12718 11388 12724
rect 10782 12679 10838 12688
rect 10796 12306 10824 12679
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11256 12345 11284 12378
rect 11242 12336 11298 12345
rect 10784 12300 10836 12306
rect 11242 12271 11298 12280
rect 10784 12242 10836 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10796 11898 10824 12242
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9954 9208 10010 9217
rect 9954 9143 10010 9152
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9968 8566 9996 8978
rect 9956 8560 10008 8566
rect 9862 8528 9918 8537
rect 9956 8502 10008 8508
rect 9862 8463 9918 8472
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9494 6896 9550 6905
rect 9494 6831 9550 6840
rect 4802 6624 4858 6633
rect 4802 6559 4858 6568
rect 4816 6458 4844 6559
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9508 6361 9536 6394
rect 9494 6352 9550 6361
rect 9494 6287 9550 6296
rect 9692 5778 9720 8230
rect 9968 8090 9996 8502
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 9692 5370 9720 5714
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9968 5030 9996 5714
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 4540 4814 4752 4842
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 3882 3768 3938 3777
rect 3882 3703 3938 3712
rect 2976 2774 3096 2802
rect 2976 377 3004 2774
rect 4540 2666 4568 4814
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 4540 2638 4660 2666
rect 4632 480 4660 2638
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 10060 921 10088 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10606 10824 11086
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10152 10146 10180 10474
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10888 10266 10916 11630
rect 10980 11218 11008 12174
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11256 11286 11284 11834
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10152 10118 10364 10146
rect 10336 10062 10364 10118
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10336 9722 10364 9998
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 9382 10732 9522
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10152 9178 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10704 8838 10732 9318
rect 10782 9208 10838 9217
rect 10782 9143 10838 9152
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10598 8392 10654 8401
rect 10598 8327 10600 8336
rect 10652 8327 10654 8336
rect 10600 8298 10652 8304
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 8022 10180 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10704 7954 10732 8774
rect 10796 8634 10824 9143
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10428 7546 10456 7890
rect 10704 7546 10732 7890
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10980 5914 11008 11154
rect 11256 10810 11284 11222
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 11256 10130 11284 10746
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11164 1465 11192 9590
rect 11440 6225 11468 13806
rect 11532 12986 11560 15302
rect 11702 15263 11758 15272
rect 11716 14550 11744 15263
rect 11992 15065 12020 15574
rect 11978 15056 12034 15065
rect 11978 14991 12034 15000
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11716 14074 11744 14486
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11808 13326 11836 14758
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11808 12646 11836 13262
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 11694 11560 12242
rect 11716 11778 11744 12378
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11898 11836 12174
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11716 11750 11836 11778
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11808 11558 11836 11750
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 11354 11836 11494
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10538 12020 10950
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9382 11560 10066
rect 11716 9722 11744 10134
rect 11992 10062 12020 10474
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11532 6769 11560 9318
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11624 8498 11652 8774
rect 11716 8566 11744 9658
rect 11992 9178 12020 9998
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11624 8090 11652 8434
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11518 6760 11574 6769
rect 11518 6695 11574 6704
rect 11426 6216 11482 6225
rect 11426 6151 11482 6160
rect 12084 3505 12112 17478
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12176 13308 12204 17002
rect 12544 16794 12572 18362
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12532 16108 12584 16114
rect 12532 16050 12584 16056
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15473 12480 15846
rect 12544 15706 12572 16050
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12438 15464 12494 15473
rect 12348 15428 12400 15434
rect 12438 15399 12494 15408
rect 12348 15370 12400 15376
rect 12360 14618 12388 15370
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12254 14512 12310 14521
rect 12254 14447 12310 14456
rect 12268 14414 12296 14447
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12268 13462 12296 14350
rect 12544 13530 12572 15642
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12176 13280 12388 13308
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12268 10266 12296 11086
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12360 9654 12388 13280
rect 12544 12714 12572 13466
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12636 12594 12664 14826
rect 12728 12986 12756 21830
rect 12912 20466 12940 27390
rect 13084 25152 13136 25158
rect 13084 25094 13136 25100
rect 13096 24818 13124 25094
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13096 22506 13124 24754
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 13372 19310 13400 27520
rect 13924 27418 13952 27520
rect 13832 27390 13952 27418
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13648 22574 13676 23462
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13648 21486 13676 21830
rect 13832 21593 13860 27390
rect 14568 24857 14596 27520
rect 15120 27418 15148 27520
rect 15672 27418 15700 27520
rect 14752 27390 15148 27418
rect 15580 27390 15700 27418
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13924 23594 13952 24006
rect 13912 23588 13964 23594
rect 13912 23530 13964 23536
rect 13924 22438 13952 23530
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13924 22030 13952 22374
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 14384 21690 14412 22442
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 13818 21584 13874 21593
rect 13818 21519 13874 21528
rect 13636 21480 13688 21486
rect 13636 21422 13688 21428
rect 13648 21146 13676 21422
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13464 20466 13492 20946
rect 13648 20806 13676 21082
rect 13636 20800 13688 20806
rect 14372 20800 14424 20806
rect 13636 20742 13688 20748
rect 13818 20768 13874 20777
rect 14372 20742 14424 20748
rect 13818 20703 13874 20712
rect 13832 20602 13860 20703
rect 14384 20641 14412 20742
rect 14370 20632 14426 20641
rect 13820 20596 13872 20602
rect 14370 20567 14426 20576
rect 13820 20538 13872 20544
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13464 20058 13492 20402
rect 13832 20398 13860 20538
rect 13910 20496 13966 20505
rect 14384 20466 14412 20567
rect 13910 20431 13966 20440
rect 14372 20460 14424 20466
rect 13820 20392 13872 20398
rect 13820 20334 13872 20340
rect 13924 20330 13952 20431
rect 14372 20402 14424 20408
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13740 19718 13768 20198
rect 13924 20058 13952 20266
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13740 19174 13768 19654
rect 14016 19281 14044 20198
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 19378 14504 19654
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14002 19272 14058 19281
rect 14186 19272 14242 19281
rect 14002 19207 14058 19216
rect 14096 19236 14148 19242
rect 14186 19207 14242 19216
rect 14096 19178 14148 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13464 18766 13492 19110
rect 14108 18970 14136 19178
rect 14200 19174 14228 19207
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14476 18902 14504 19314
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14464 18896 14516 18902
rect 14464 18838 14516 18844
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13464 18222 13492 18702
rect 14660 18630 14688 19110
rect 14752 18873 14780 27390
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15580 24313 15608 27390
rect 15658 24576 15714 24585
rect 15658 24511 15714 24520
rect 15672 24410 15700 24511
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15566 24304 15622 24313
rect 15384 24268 15436 24274
rect 15566 24239 15622 24248
rect 15384 24210 15436 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15396 23594 15424 24210
rect 16224 23730 16252 27520
rect 16776 24857 16804 27520
rect 16578 24848 16634 24857
rect 16578 24783 16634 24792
rect 16762 24848 16818 24857
rect 16762 24783 16818 24792
rect 16486 23896 16542 23905
rect 16486 23831 16488 23840
rect 16540 23831 16542 23840
rect 16488 23802 16540 23808
rect 15476 23724 15528 23730
rect 15476 23666 15528 23672
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 14832 23588 14884 23594
rect 14832 23530 14884 23536
rect 15384 23588 15436 23594
rect 15384 23530 15436 23536
rect 14738 18864 14794 18873
rect 14738 18799 14794 18808
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13832 17270 13860 18566
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13924 17338 13952 17682
rect 14016 17610 14044 18090
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 17270 14044 17546
rect 14568 17270 14596 17614
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16794 12848 17138
rect 13450 17096 13506 17105
rect 13450 17031 13452 17040
rect 13504 17031 13506 17040
rect 13452 17002 13504 17008
rect 14752 16794 14780 17478
rect 14844 17338 14872 23530
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23361 15240 23462
rect 15198 23352 15254 23361
rect 15198 23287 15254 23296
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22438 15332 23122
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18426 15332 18838
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15200 18216 15252 18222
rect 15120 18164 15200 18170
rect 15120 18158 15252 18164
rect 15120 18142 15240 18158
rect 15120 17882 15148 18142
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15396 17649 15424 19790
rect 15382 17640 15438 17649
rect 15292 17604 15344 17610
rect 15382 17575 15438 17584
rect 15292 17546 15344 17552
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17338 15332 17546
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14554 16688 14610 16697
rect 14554 16623 14556 16632
rect 14608 16623 14610 16632
rect 14556 16594 14608 16600
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 13802 12848 15982
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15706 12940 15846
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12912 15434 12940 15642
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 13372 14890 13400 15506
rect 13464 15502 13492 16390
rect 13556 15910 13584 16526
rect 14568 15978 14596 16594
rect 14738 16416 14794 16425
rect 14738 16351 14794 16360
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13188 14482 13216 14758
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13188 14074 13216 14418
rect 13360 14408 13412 14414
rect 13358 14376 13360 14385
rect 13464 14396 13492 15438
rect 13412 14376 13492 14396
rect 13414 14368 13492 14376
rect 13358 14311 13414 14320
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12544 12566 12664 12594
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12452 9382 12480 9415
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 8430 12480 8978
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12544 7857 12572 12566
rect 12728 12442 12756 12650
rect 13188 12646 13216 13670
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13096 11150 13124 12038
rect 13188 11694 13216 12582
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13464 11694 13492 12038
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13188 10606 13216 11630
rect 13464 11354 13492 11630
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13358 11112 13414 11121
rect 13358 11047 13360 11056
rect 13412 11047 13414 11056
rect 13360 11018 13412 11024
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9654 12848 9862
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12728 9042 12756 9386
rect 12820 9042 12848 9590
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8634 12848 8978
rect 12912 8838 12940 9454
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13004 9217 13032 9318
rect 12990 9208 13046 9217
rect 12990 9143 12992 9152
rect 13044 9143 13046 9152
rect 12992 9114 13044 9120
rect 13004 9083 13032 9114
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12912 8090 12940 8774
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12530 7848 12586 7857
rect 12530 7783 12586 7792
rect 13464 7449 13492 9318
rect 13450 7440 13506 7449
rect 13450 7375 13506 7384
rect 12070 3496 12126 3505
rect 12070 3431 12126 3440
rect 13556 1737 13584 15846
rect 13740 14822 13768 15846
rect 14568 15706 14596 15914
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13634 14648 13690 14657
rect 13634 14583 13636 14592
rect 13688 14583 13690 14592
rect 13636 14554 13688 14560
rect 13740 13870 13768 14758
rect 13832 14618 13860 15302
rect 14108 15162 14136 15438
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13910 13968 13966 13977
rect 13910 13903 13966 13912
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13820 12912 13872 12918
rect 13818 12880 13820 12889
rect 13872 12880 13874 12889
rect 13818 12815 13874 12824
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12209 13860 12718
rect 13818 12200 13874 12209
rect 13818 12135 13874 12144
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11801 13676 12038
rect 13634 11792 13690 11801
rect 13634 11727 13690 11736
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11354 13768 11562
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 10198 13768 11290
rect 13924 11234 13952 13903
rect 14108 13802 14136 15098
rect 14200 14890 14228 15302
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14200 14414 14228 14826
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14108 13410 14136 13738
rect 14200 13734 14228 14350
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14200 13530 14228 13670
rect 14476 13530 14504 14554
rect 14752 14550 14780 16351
rect 14844 16046 14872 16934
rect 15488 16794 15516 23666
rect 16394 23624 16450 23633
rect 16592 23610 16620 24783
rect 17420 24585 17448 27520
rect 17406 24576 17462 24585
rect 17406 24511 17462 24520
rect 17314 24440 17370 24449
rect 17314 24375 17316 24384
rect 17368 24375 17370 24384
rect 17316 24346 17368 24352
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 16394 23559 16450 23568
rect 16500 23582 16620 23610
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16182 15332 16594
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 15290 16008 15346 16017
rect 15290 15943 15346 15952
rect 15304 15570 15332 15943
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 14906 15332 15506
rect 15304 14878 15424 14906
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 14740 14544 14792 14550
rect 15304 14521 15332 14758
rect 15396 14618 15424 14878
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 14740 14486 14792 14492
rect 15290 14512 15346 14521
rect 15290 14447 15346 14456
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14108 13382 14228 13410
rect 14200 13326 14228 13382
rect 14188 13320 14240 13326
rect 14186 13288 14188 13297
rect 15476 13320 15528 13326
rect 14240 13288 14242 13297
rect 15476 13262 15528 13268
rect 14186 13223 14242 13232
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14844 12782 14872 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15108 12912 15160 12918
rect 15106 12880 15108 12889
rect 15160 12880 15162 12889
rect 15106 12815 15162 12824
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15488 12714 15516 13262
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14844 12481 14872 12582
rect 14830 12472 14886 12481
rect 14830 12407 14886 12416
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14016 12209 14044 12242
rect 14844 12238 14872 12407
rect 15212 12238 15240 12650
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 14464 12232 14516 12238
rect 14002 12200 14058 12209
rect 14464 12174 14516 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 14002 12135 14058 12144
rect 14016 11558 14044 12135
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14476 11354 14504 12174
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11354 14780 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11880 15332 12310
rect 15488 11898 15516 12650
rect 15120 11852 15332 11880
rect 15476 11892 15528 11898
rect 15120 11558 15148 11852
rect 15476 11834 15528 11840
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 13924 11206 14044 11234
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10810 13952 11086
rect 14016 11014 14044 11206
rect 15120 11082 15148 11494
rect 15292 11212 15344 11218
rect 15292 11154 15344 11160
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 14016 10674 14044 10950
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10198 14044 10610
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13832 9382 13860 10066
rect 14016 9722 14044 10134
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14568 9518 14596 9930
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 14568 8906 14596 9454
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13542 1728 13598 1737
rect 13542 1663 13598 1672
rect 11150 1456 11206 1465
rect 11150 1391 11206 1400
rect 10046 912 10102 921
rect 10046 847 10102 856
rect 13924 480 13952 4966
rect 14844 2961 14872 10406
rect 15120 10266 15148 10474
rect 15304 10470 15332 11154
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15488 10130 15516 11834
rect 15580 10810 15608 22510
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 19009 15792 19110
rect 15750 19000 15806 19009
rect 15750 18935 15806 18944
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15672 18358 15700 18566
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17066 15884 17614
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15856 16794 15884 17002
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15856 16250 15884 16730
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15948 15706 15976 22374
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15948 13870 15976 14418
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15856 12481 15884 13330
rect 15842 12472 15898 12481
rect 15842 12407 15898 12416
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10266 15608 10406
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15580 9178 15608 10202
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15764 9654 15792 10066
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15764 9450 15792 9590
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15856 7993 15884 11494
rect 15842 7984 15898 7993
rect 15842 7919 15898 7928
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 14830 2952 14886 2961
rect 14830 2887 14886 2896
rect 15948 2553 15976 13806
rect 16040 12889 16068 23462
rect 16408 22778 16436 23559
rect 16500 23322 16528 23582
rect 17144 23526 17172 24210
rect 17972 23905 18000 27520
rect 18418 24168 18474 24177
rect 18418 24103 18474 24112
rect 17958 23896 18014 23905
rect 18432 23866 18460 24103
rect 17958 23831 18014 23840
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18236 23656 18288 23662
rect 18234 23624 18236 23633
rect 18288 23624 18290 23633
rect 18234 23559 18290 23568
rect 16580 23520 16632 23526
rect 17132 23520 17184 23526
rect 16580 23462 16632 23468
rect 16762 23488 16818 23497
rect 16488 23316 16540 23322
rect 16488 23258 16540 23264
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16212 22500 16264 22506
rect 16212 22442 16264 22448
rect 16224 12986 16252 22442
rect 16592 19530 16620 23462
rect 18524 23497 18552 27520
rect 19076 24449 19104 27520
rect 19628 25786 19656 27520
rect 19444 25758 19656 25786
rect 19062 24440 19118 24449
rect 19062 24375 19118 24384
rect 19444 23746 19472 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19522 23896 19578 23905
rect 19522 23831 19524 23840
rect 19576 23831 19578 23840
rect 19524 23802 19576 23808
rect 19444 23718 19564 23746
rect 19432 23656 19484 23662
rect 19260 23604 19432 23610
rect 19260 23598 19484 23604
rect 19260 23582 19472 23598
rect 17132 23462 17184 23468
rect 18510 23488 18566 23497
rect 16762 23423 16818 23432
rect 18510 23423 18566 23432
rect 16776 23322 16804 23423
rect 19260 23322 19288 23582
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 17316 23180 17368 23186
rect 17316 23122 17368 23128
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 17328 22438 17356 23122
rect 17880 22506 17908 23122
rect 17868 22500 17920 22506
rect 17868 22442 17920 22448
rect 18892 22438 18920 23122
rect 19352 23050 19380 23462
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 16854 22128 16910 22137
rect 16854 22063 16910 22072
rect 16592 19502 16712 19530
rect 16578 19408 16634 19417
rect 16578 19343 16634 19352
rect 16592 18970 16620 19343
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16394 18184 16450 18193
rect 16394 18119 16450 18128
rect 16408 18086 16436 18119
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16500 17626 16528 17682
rect 16500 17598 16620 17626
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16316 15910 16344 16526
rect 16592 16114 16620 17598
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15502 16344 15846
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16316 14958 16344 15438
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16394 14920 16450 14929
rect 16394 14855 16450 14864
rect 16408 14822 16436 14855
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16408 14074 16436 14486
rect 16592 14414 16620 15506
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16592 14074 16620 14350
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16026 12880 16082 12889
rect 16026 12815 16082 12824
rect 16408 11762 16436 14010
rect 16592 13530 16620 14010
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16578 12472 16634 12481
rect 16578 12407 16634 12416
rect 16592 12170 16620 12407
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16408 11354 16436 11698
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16488 11144 16540 11150
rect 16540 11104 16620 11132
rect 16488 11086 16540 11092
rect 16592 10810 16620 11104
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16040 10198 16068 10610
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16394 10160 16450 10169
rect 16040 9722 16068 10134
rect 16394 10095 16450 10104
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16040 9178 16068 9658
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16408 9042 16436 10095
rect 16684 9178 16712 19502
rect 16868 17746 16896 22063
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16868 17338 16896 17682
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16868 16250 16896 16594
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16868 15706 16896 16186
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16868 15026 16896 15642
rect 17052 15638 17080 17478
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16868 14618 16896 14758
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 12102 17264 12582
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11898 17264 12038
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17144 11558 17172 11698
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 16762 10704 16818 10713
rect 16762 10639 16818 10648
rect 16776 10606 16804 10639
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 17144 10266 17172 11494
rect 17328 10810 17356 22374
rect 18050 17912 18106 17921
rect 18050 17847 18106 17856
rect 17866 17776 17922 17785
rect 17866 17711 17868 17720
rect 17920 17711 17922 17720
rect 17868 17682 17920 17688
rect 18064 17134 18092 17847
rect 18236 17264 18288 17270
rect 18234 17232 18236 17241
rect 18288 17232 18290 17241
rect 18234 17167 18290 17176
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17972 16697 18000 16730
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18064 15609 18092 15982
rect 18050 15600 18106 15609
rect 18050 15535 18106 15544
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17512 14618 17540 14826
rect 18892 14657 18920 22374
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19062 16144 19118 16153
rect 19062 16079 19118 16088
rect 19076 16046 19104 16079
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19246 16008 19302 16017
rect 19246 15943 19302 15952
rect 19260 15910 19288 15943
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 18878 14648 18934 14657
rect 17500 14612 17552 14618
rect 18878 14583 18934 14592
rect 17500 14554 17552 14560
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17788 12714 17816 13262
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17788 12306 17816 12650
rect 19168 12646 19196 13330
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12442 19196 12582
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17788 11898 17816 12242
rect 17958 12200 18014 12209
rect 17958 12135 18014 12144
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17774 11656 17830 11665
rect 17972 11626 18000 12135
rect 18064 11762 18092 12242
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17774 11591 17830 11600
rect 17960 11620 18012 11626
rect 17788 11354 17816 11591
rect 17960 11562 18012 11568
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17604 10470 17632 11154
rect 19352 10826 19380 17206
rect 19430 15464 19486 15473
rect 19430 15399 19486 15408
rect 19444 14958 19472 15399
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19430 13288 19486 13297
rect 19430 13223 19432 13232
rect 19484 13223 19486 13232
rect 19432 13194 19484 13200
rect 19536 11665 19564 23718
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20272 17270 20300 27520
rect 20824 24177 20852 27520
rect 20810 24168 20866 24177
rect 20810 24103 20866 24112
rect 20626 24032 20682 24041
rect 20626 23967 20682 23976
rect 20640 23866 20668 23967
rect 21376 23905 21404 27520
rect 21822 24440 21878 24449
rect 21822 24375 21824 24384
rect 21876 24375 21878 24384
rect 21824 24346 21876 24352
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21362 23896 21418 23905
rect 20628 23860 20680 23866
rect 21362 23831 21418 23840
rect 20628 23802 20680 23808
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20824 22438 20852 23122
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20260 17264 20312 17270
rect 20260 17206 20312 17212
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19522 11656 19578 11665
rect 19522 11591 19578 11600
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20824 11257 20852 22374
rect 21086 21448 21142 21457
rect 21086 21383 21142 21392
rect 21100 15706 21128 21383
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20916 15094 20944 15506
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 21192 13530 21220 23598
rect 21652 23594 21680 24210
rect 21928 24041 21956 27520
rect 21914 24032 21970 24041
rect 21914 23967 21970 23976
rect 21730 23896 21786 23905
rect 21730 23831 21732 23840
rect 21784 23831 21786 23840
rect 21732 23802 21784 23808
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21652 23322 21680 23530
rect 22284 23520 22336 23526
rect 22284 23462 22336 23468
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22204 22438 22232 23122
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20902 13424 20958 13433
rect 20902 13359 20904 13368
rect 20956 13359 20958 13368
rect 20904 13330 20956 13336
rect 20916 12986 20944 13330
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 22020 12345 22048 12378
rect 21178 12336 21234 12345
rect 21178 12271 21234 12280
rect 22006 12336 22062 12345
rect 22006 12271 22062 12280
rect 21192 11694 21220 12271
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 22020 11558 22048 12174
rect 22204 11898 22232 22374
rect 22296 12986 22324 23462
rect 22374 23352 22430 23361
rect 22374 23287 22376 23296
rect 22428 23287 22430 23296
rect 22376 23258 22428 23264
rect 22480 21457 22508 27520
rect 23124 23905 23152 27520
rect 23676 24449 23704 27520
rect 23662 24440 23718 24449
rect 23662 24375 23718 24384
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 23110 23896 23166 23905
rect 23110 23831 23166 23840
rect 23308 23526 23336 24210
rect 24228 23610 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 27520
rect 25332 24410 25360 27520
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 24950 23896 25006 23905
rect 24768 23860 24820 23866
rect 24950 23831 24952 23840
rect 24768 23802 24820 23808
rect 25004 23831 25006 23840
rect 24952 23802 25004 23808
rect 24768 23656 24820 23662
rect 24228 23582 24348 23610
rect 24768 23598 24820 23604
rect 23296 23520 23348 23526
rect 24216 23520 24268 23526
rect 23296 23462 23348 23468
rect 24030 23488 24086 23497
rect 24216 23462 24268 23468
rect 24030 23423 24086 23432
rect 24044 23322 24072 23423
rect 24032 23316 24084 23322
rect 24032 23258 24084 23264
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23860 22710 23888 23122
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 22560 22568 22612 22574
rect 22560 22510 22612 22516
rect 22466 21448 22522 21457
rect 22466 21383 22522 21392
rect 22572 14929 22600 22510
rect 23664 19304 23716 19310
rect 23662 19272 23664 19281
rect 23716 19272 23718 19281
rect 23662 19207 23718 19216
rect 22558 14920 22614 14929
rect 22558 14855 22614 14864
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 11937 22324 12718
rect 24228 12345 24256 23462
rect 24320 23361 24348 23582
rect 24306 23352 24362 23361
rect 24306 23287 24362 23296
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24780 19174 24808 23598
rect 25976 23497 26004 27520
rect 25962 23488 26018 23497
rect 25962 23423 26018 23432
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 26252 12753 26280 21354
rect 26528 18193 26556 27520
rect 27080 23905 27108 27520
rect 27066 23896 27122 23905
rect 27066 23831 27122 23840
rect 27632 21418 27660 27520
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 26514 18184 26570 18193
rect 26514 18119 26570 18128
rect 26238 12744 26294 12753
rect 26238 12679 26294 12688
rect 24214 12336 24270 12345
rect 24214 12271 24270 12280
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 22282 11928 22338 11937
rect 22192 11892 22244 11898
rect 24289 11920 24585 11940
rect 22282 11863 22338 11872
rect 22192 11834 22244 11840
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 20810 11248 20866 11257
rect 20810 11183 20866 11192
rect 22020 11121 22048 11494
rect 22006 11112 22062 11121
rect 22006 11047 22062 11056
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19260 10810 19380 10826
rect 19248 10804 19380 10810
rect 19300 10798 19380 10804
rect 19248 10746 19300 10752
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17604 9722 17632 10406
rect 18248 9722 18276 10542
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 16946 9616 17002 9625
rect 16946 9551 17002 9560
rect 16960 9518 16988 9551
rect 16948 9512 17000 9518
rect 18052 9512 18104 9518
rect 16948 9454 17000 9460
rect 18050 9480 18052 9489
rect 18104 9480 18106 9489
rect 18050 9415 18106 9424
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16408 8634 16436 8978
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 23202 3496 23258 3505
rect 23202 3431 23258 3440
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 15934 2544 15990 2553
rect 15934 2479 15990 2488
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 23216 480 23244 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 2962 368 3018 377
rect 2962 303 3018 312
rect 4618 0 4674 480
rect 13910 0 13966 480
rect 23202 0 23258 480
<< via2 >>
rect 3790 27648 3846 27704
rect 1306 23568 1362 23624
rect 1674 23296 1730 23352
rect 1582 23160 1638 23216
rect 1582 22480 1638 22536
rect 1582 21392 1638 21448
rect 1582 19624 1638 19680
rect 1490 19080 1546 19136
rect 1398 17448 1454 17504
rect 2318 24828 2320 24848
rect 2320 24828 2372 24848
rect 2372 24828 2374 24848
rect 2318 24792 2374 24828
rect 2134 23024 2190 23080
rect 1582 17040 1638 17096
rect 846 14728 902 14784
rect 1490 14592 1546 14648
rect 1858 14728 1914 14784
rect 1766 14048 1822 14104
rect 1582 12280 1638 12336
rect 1766 12164 1822 12200
rect 1766 12144 1768 12164
rect 1768 12144 1820 12164
rect 1820 12144 1822 12164
rect 1858 10512 1914 10568
rect 2778 26560 2834 26616
rect 3054 25356 3110 25392
rect 3054 25336 3056 25356
rect 3056 25336 3108 25356
rect 3108 25336 3110 25356
rect 2594 23160 2650 23216
rect 2778 23160 2834 23216
rect 2778 22888 2834 22944
rect 3054 24384 3110 24440
rect 2962 23160 3018 23216
rect 2870 21936 2926 21992
rect 2686 20868 2742 20904
rect 2686 20848 2688 20868
rect 2688 20848 2740 20868
rect 2740 20848 2742 20868
rect 3238 24112 3294 24168
rect 3422 24248 3478 24304
rect 3330 23704 3386 23760
rect 2962 20304 3018 20360
rect 2686 18536 2742 18592
rect 2502 17992 2558 18048
rect 2594 17448 2650 17504
rect 2134 16496 2190 16552
rect 3146 21120 3202 21176
rect 3698 24656 3754 24712
rect 4158 27104 4214 27160
rect 4066 24520 4122 24576
rect 3790 22888 3846 22944
rect 3606 20440 3662 20496
rect 2962 17448 3018 17504
rect 2042 9152 2098 9208
rect 1674 8508 1676 8528
rect 1676 8508 1728 8528
rect 1728 8508 1730 8528
rect 1674 8472 1730 8508
rect 2778 14592 2834 14648
rect 2870 14184 2926 14240
rect 3054 14048 3110 14104
rect 2410 11056 2466 11112
rect 2318 9560 2374 9616
rect 3606 17992 3662 18048
rect 3882 17856 3938 17912
rect 3514 15408 3570 15464
rect 3514 15000 3570 15056
rect 3330 14320 3386 14376
rect 3238 12552 3294 12608
rect 3606 13812 3608 13832
rect 3608 13812 3660 13832
rect 3660 13812 3662 13832
rect 3606 13776 3662 13812
rect 3514 13524 3570 13560
rect 3514 13504 3516 13524
rect 3516 13504 3568 13524
rect 3568 13504 3570 13524
rect 4526 26016 4582 26072
rect 4434 24248 4490 24304
rect 4618 24656 4674 24712
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5446 23704 5502 23760
rect 5078 23296 5134 23352
rect 4618 22888 4674 22944
rect 4894 20340 4896 20360
rect 4896 20340 4948 20360
rect 4948 20340 4950 20360
rect 4894 20304 4950 20340
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5538 23160 5594 23216
rect 6550 24792 6606 24848
rect 6182 24692 6184 24712
rect 6184 24692 6236 24712
rect 6236 24692 6238 24712
rect 6182 24656 6238 24692
rect 6458 23860 6514 23896
rect 6458 23840 6460 23860
rect 6460 23840 6512 23860
rect 6512 23840 6514 23860
rect 5998 23024 6054 23080
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5630 22636 5686 22672
rect 5630 22616 5632 22636
rect 5632 22616 5684 22636
rect 5684 22616 5686 22636
rect 6366 22480 6422 22536
rect 5354 21412 5410 21448
rect 5354 21392 5356 21412
rect 5356 21392 5408 21412
rect 5408 21392 5410 21412
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5078 19352 5134 19408
rect 4526 17448 4582 17504
rect 4342 17176 4398 17232
rect 4158 16904 4214 16960
rect 4066 16632 4122 16688
rect 4066 15680 4122 15736
rect 4066 15544 4122 15600
rect 3974 15136 4030 15192
rect 3882 14864 3938 14920
rect 3882 14476 3938 14512
rect 3882 14456 3884 14476
rect 3884 14456 3936 14476
rect 3936 14456 3938 14476
rect 4066 14612 4122 14648
rect 4066 14592 4068 14612
rect 4068 14592 4120 14612
rect 4120 14592 4122 14612
rect 4158 14184 4214 14240
rect 4250 12824 4306 12880
rect 4066 12688 4122 12744
rect 3698 11056 3754 11112
rect 3790 10376 3846 10432
rect 4066 10648 4122 10704
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5078 17720 5134 17776
rect 4526 15680 4582 15736
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6458 16396 6460 16416
rect 6460 16396 6512 16416
rect 6512 16396 6514 16416
rect 6458 16360 6514 16396
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4526 14864 4582 14920
rect 5170 15952 5226 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5078 14728 5134 14784
rect 5262 14764 5264 14784
rect 5264 14764 5316 14784
rect 5316 14764 5318 14784
rect 5262 14728 5318 14764
rect 4986 12588 4988 12608
rect 4988 12588 5040 12608
rect 5040 12588 5042 12608
rect 4986 12552 5042 12588
rect 4526 9968 4582 10024
rect 7010 24112 7066 24168
rect 7102 23568 7158 23624
rect 8206 24812 8262 24848
rect 8206 24792 8208 24812
rect 8208 24792 8260 24812
rect 8260 24792 8262 24812
rect 8114 24656 8170 24712
rect 8022 24404 8078 24440
rect 8022 24384 8024 24404
rect 8024 24384 8076 24404
rect 8076 24384 8078 24404
rect 7654 21120 7710 21176
rect 7654 20984 7710 21040
rect 7194 20440 7250 20496
rect 6918 15700 6974 15736
rect 6918 15680 6920 15700
rect 6920 15680 6972 15700
rect 6972 15680 6974 15700
rect 6642 15544 6698 15600
rect 5998 14456 6054 14512
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5538 13912 5594 13968
rect 5170 13368 5226 13424
rect 6274 13776 6330 13832
rect 5262 12552 5318 12608
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5814 12844 5870 12880
rect 5814 12824 5816 12844
rect 5816 12824 5868 12844
rect 5868 12824 5870 12844
rect 6090 12688 6146 12744
rect 5630 12552 5686 12608
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6182 11736 6238 11792
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6550 10412 6552 10432
rect 6552 10412 6604 10432
rect 6604 10412 6606 10432
rect 6550 10376 6606 10412
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 3882 6704 3938 6760
rect 3790 4800 3846 4856
rect 4066 7928 4122 7984
rect 4066 7112 4122 7168
rect 4066 6840 4122 6896
rect 3974 5344 4030 5400
rect 6366 9424 6422 9480
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 7378 19372 7434 19408
rect 7378 19352 7380 19372
rect 7380 19352 7432 19372
rect 7432 19352 7434 19372
rect 7286 18808 7342 18864
rect 7930 19760 7986 19816
rect 8114 20032 8170 20088
rect 7470 17620 7472 17640
rect 7472 17620 7524 17640
rect 7524 17620 7526 17640
rect 7470 17584 7526 17620
rect 8114 19216 8170 19272
rect 8298 20576 8354 20632
rect 8298 18028 8300 18048
rect 8300 18028 8352 18048
rect 8352 18028 8354 18048
rect 8298 17992 8354 18028
rect 9678 23840 9734 23896
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10690 23704 10746 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9954 22616 10010 22672
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10046 22072 10102 22128
rect 9402 20712 9458 20768
rect 8482 17856 8538 17912
rect 8114 17584 8170 17640
rect 9678 19760 9734 19816
rect 9586 19386 9642 19442
rect 10138 21528 10194 21584
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10414 20476 10416 20496
rect 10416 20476 10468 20496
rect 10468 20476 10470 20496
rect 10414 20440 10470 20476
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10046 20052 10102 20088
rect 10046 20032 10048 20052
rect 10048 20032 10100 20052
rect 10100 20032 10102 20052
rect 11150 20984 11206 21040
rect 11794 24676 11850 24712
rect 11794 24656 11796 24676
rect 11796 24656 11848 24676
rect 11848 24656 11850 24676
rect 12254 23296 12310 23352
rect 12438 22500 12494 22536
rect 12438 22480 12440 22500
rect 12440 22480 12492 22500
rect 12492 22480 12494 22500
rect 11610 21392 11666 21448
rect 9678 17176 9734 17232
rect 9770 16768 9826 16824
rect 9770 16668 9772 16688
rect 9772 16668 9824 16688
rect 9824 16668 9826 16688
rect 9770 16632 9826 16668
rect 8758 16496 8814 16552
rect 8482 16360 8538 16416
rect 8758 16360 8814 16416
rect 7194 15408 7250 15464
rect 7746 15444 7748 15464
rect 7748 15444 7800 15464
rect 7800 15444 7802 15464
rect 7746 15408 7802 15444
rect 7286 15272 7342 15328
rect 8390 14864 8446 14920
rect 7470 14728 7526 14784
rect 9494 15544 9550 15600
rect 8022 14356 8024 14376
rect 8024 14356 8076 14376
rect 8076 14356 8078 14376
rect 8022 14320 8078 14356
rect 8574 13776 8630 13832
rect 7654 13252 7710 13288
rect 7654 13232 7656 13252
rect 7656 13232 7708 13252
rect 7708 13232 7710 13252
rect 7470 11600 7526 11656
rect 7930 11600 7986 11656
rect 7010 9560 7066 9616
rect 7654 10104 7710 10160
rect 7746 8880 7802 8936
rect 9034 14612 9090 14648
rect 9034 14592 9036 14612
rect 9036 14592 9088 14612
rect 9088 14592 9090 14612
rect 9402 13504 9458 13560
rect 9678 9596 9680 9616
rect 9680 9596 9732 9616
rect 9732 9596 9734 9616
rect 9678 9560 9734 9596
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10690 18944 10746 19000
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10966 17856 11022 17912
rect 11886 20324 11942 20360
rect 11886 20304 11888 20324
rect 11888 20304 11940 20324
rect 11940 20304 11942 20324
rect 12070 19624 12126 19680
rect 12530 19624 12586 19680
rect 11150 16632 11206 16688
rect 11242 16244 11298 16280
rect 11242 16224 11244 16244
rect 11244 16224 11296 16244
rect 11296 16224 11298 16244
rect 10782 16088 10838 16144
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10046 14320 10102 14376
rect 11794 15428 11850 15464
rect 11794 15408 11796 15428
rect 11796 15408 11848 15428
rect 11848 15408 11850 15428
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10046 13504 10102 13560
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11150 13932 11206 13968
rect 11150 13912 11152 13932
rect 11152 13912 11204 13932
rect 11204 13912 11206 13932
rect 10782 12688 10838 12744
rect 11242 12280 11298 12336
rect 9954 9152 10010 9208
rect 9862 8472 9918 8528
rect 9494 6840 9550 6896
rect 4802 6568 4858 6624
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 9494 6296 9550 6352
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 4066 4256 4122 4312
rect 3882 3712 3938 3768
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10782 9152 10838 9208
rect 10598 8356 10654 8392
rect 10598 8336 10600 8356
rect 10600 8336 10652 8356
rect 10652 8336 10654 8356
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 11702 15272 11758 15328
rect 11978 15000 12034 15056
rect 11518 6704 11574 6760
rect 11426 6160 11482 6216
rect 12438 15408 12494 15464
rect 12254 14456 12310 14512
rect 14554 24792 14610 24848
rect 13818 21528 13874 21584
rect 13818 20712 13874 20768
rect 14370 20576 14426 20632
rect 13910 20440 13966 20496
rect 14002 19216 14058 19272
rect 14186 19216 14242 19272
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15658 24520 15714 24576
rect 15566 24248 15622 24304
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 16578 24792 16634 24848
rect 16762 24792 16818 24848
rect 16486 23860 16542 23896
rect 16486 23840 16488 23860
rect 16488 23840 16540 23860
rect 16540 23840 16542 23860
rect 14738 18808 14794 18864
rect 13450 17060 13506 17096
rect 13450 17040 13452 17060
rect 13452 17040 13504 17060
rect 13504 17040 13506 17060
rect 15198 23296 15254 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15382 17584 15438 17640
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14554 16652 14610 16688
rect 14554 16632 14556 16652
rect 14556 16632 14608 16652
rect 14608 16632 14610 16652
rect 14738 16360 14794 16416
rect 13358 14356 13360 14376
rect 13360 14356 13412 14376
rect 13412 14356 13414 14376
rect 13358 14320 13414 14356
rect 12438 9424 12494 9480
rect 13358 11076 13414 11112
rect 13358 11056 13360 11076
rect 13360 11056 13412 11076
rect 13412 11056 13414 11076
rect 12990 9172 13046 9208
rect 12990 9152 12992 9172
rect 12992 9152 13044 9172
rect 13044 9152 13046 9172
rect 12530 7792 12586 7848
rect 13450 7384 13506 7440
rect 12070 3440 12126 3496
rect 13634 14612 13690 14648
rect 13634 14592 13636 14612
rect 13636 14592 13688 14612
rect 13688 14592 13690 14612
rect 13910 13912 13966 13968
rect 13818 12860 13820 12880
rect 13820 12860 13872 12880
rect 13872 12860 13874 12880
rect 13818 12824 13874 12860
rect 13818 12144 13874 12200
rect 13634 11736 13690 11792
rect 16394 23568 16450 23624
rect 17406 24520 17462 24576
rect 17314 24404 17370 24440
rect 17314 24384 17316 24404
rect 17316 24384 17368 24404
rect 17368 24384 17370 24404
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15290 15952 15346 16008
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15290 14456 15346 14512
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14186 13268 14188 13288
rect 14188 13268 14240 13288
rect 14240 13268 14242 13288
rect 14186 13232 14242 13268
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15106 12860 15108 12880
rect 15108 12860 15160 12880
rect 15160 12860 15162 12880
rect 15106 12824 15162 12860
rect 14830 12416 14886 12472
rect 14002 12144 14058 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 13542 1672 13598 1728
rect 11150 1400 11206 1456
rect 10046 856 10102 912
rect 15750 18944 15806 19000
rect 15842 12416 15898 12472
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15842 7928 15898 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14830 2896 14886 2952
rect 18418 24112 18474 24168
rect 17958 23840 18014 23896
rect 18234 23604 18236 23624
rect 18236 23604 18288 23624
rect 18288 23604 18290 23624
rect 18234 23568 18290 23604
rect 16762 23432 16818 23488
rect 19062 24384 19118 24440
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19522 23860 19578 23896
rect 19522 23840 19524 23860
rect 19524 23840 19576 23860
rect 19576 23840 19578 23860
rect 18510 23432 18566 23488
rect 16854 22072 16910 22128
rect 16578 19352 16634 19408
rect 16394 18128 16450 18184
rect 16394 14864 16450 14920
rect 16026 12824 16082 12880
rect 16578 12416 16634 12472
rect 16394 10104 16450 10160
rect 16762 10648 16818 10704
rect 18050 17856 18106 17912
rect 17866 17740 17922 17776
rect 17866 17720 17868 17740
rect 17868 17720 17920 17740
rect 17920 17720 17922 17740
rect 18234 17212 18236 17232
rect 18236 17212 18288 17232
rect 18288 17212 18290 17232
rect 18234 17176 18290 17212
rect 17958 16632 18014 16688
rect 18050 15544 18106 15600
rect 19062 16088 19118 16144
rect 19246 15952 19302 16008
rect 18878 14592 18934 14648
rect 17958 12144 18014 12200
rect 17774 11600 17830 11656
rect 19430 15408 19486 15464
rect 19430 13252 19486 13288
rect 19430 13232 19432 13252
rect 19432 13232 19484 13252
rect 19484 13232 19486 13252
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20810 24112 20866 24168
rect 20626 23976 20682 24032
rect 21822 24404 21878 24440
rect 21822 24384 21824 24404
rect 21824 24384 21876 24404
rect 21876 24384 21878 24404
rect 21362 23840 21418 23896
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19522 11600 19578 11656
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 21086 21392 21142 21448
rect 21914 23976 21970 24032
rect 21730 23860 21786 23896
rect 21730 23840 21732 23860
rect 21732 23840 21784 23860
rect 21784 23840 21786 23860
rect 20902 13388 20958 13424
rect 20902 13368 20904 13388
rect 20904 13368 20956 13388
rect 20956 13368 20958 13388
rect 21178 12280 21234 12336
rect 22006 12280 22062 12336
rect 22374 23316 22430 23352
rect 22374 23296 22376 23316
rect 22376 23296 22428 23316
rect 22428 23296 22430 23316
rect 23662 24384 23718 24440
rect 23110 23840 23166 23896
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24950 23860 25006 23896
rect 24950 23840 24952 23860
rect 24952 23840 25004 23860
rect 25004 23840 25006 23860
rect 24030 23432 24086 23488
rect 22466 21392 22522 21448
rect 23662 19252 23664 19272
rect 23664 19252 23716 19272
rect 23716 19252 23718 19272
rect 23662 19216 23718 19252
rect 22558 14864 22614 14920
rect 24306 23296 24362 23352
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 25962 23432 26018 23488
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 27066 23840 27122 23896
rect 26514 18128 26570 18184
rect 26238 12688 26294 12744
rect 24214 12280 24270 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 22282 11872 22338 11928
rect 20810 11192 20866 11248
rect 22006 11056 22062 11112
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 16946 9560 17002 9616
rect 18050 9460 18052 9480
rect 18052 9460 18104 9480
rect 18104 9460 18106 9480
rect 18050 9424 18106 9460
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 23202 3440 23258 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 15934 2488 15990 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 2962 312 3018 368
<< metal3 >>
rect 0 27706 480 27736
rect 3785 27706 3851 27709
rect 0 27704 3851 27706
rect 0 27648 3790 27704
rect 3846 27648 3851 27704
rect 0 27646 3851 27648
rect 0 27616 480 27646
rect 3785 27643 3851 27646
rect 0 27162 480 27192
rect 4153 27162 4219 27165
rect 0 27160 4219 27162
rect 0 27104 4158 27160
rect 4214 27104 4219 27160
rect 0 27102 4219 27104
rect 0 27072 480 27102
rect 4153 27099 4219 27102
rect 0 26618 480 26648
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 480 26558
rect 2773 26555 2839 26558
rect 0 26074 480 26104
rect 4521 26074 4587 26077
rect 0 26072 4587 26074
rect 0 26016 4526 26072
rect 4582 26016 4587 26072
rect 0 26014 4587 26016
rect 0 25984 480 26014
rect 4521 26011 4587 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 3049 25394 3115 25397
rect 0 25392 3115 25394
rect 0 25336 3054 25392
rect 3110 25336 3115 25392
rect 0 25334 3115 25336
rect 0 25304 480 25334
rect 3049 25331 3115 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 2313 24850 2379 24853
rect 6545 24850 6611 24853
rect 0 24790 1410 24850
rect 0 24760 480 24790
rect 1350 24714 1410 24790
rect 2313 24848 6611 24850
rect 2313 24792 2318 24848
rect 2374 24792 6550 24848
rect 6606 24792 6611 24848
rect 2313 24790 6611 24792
rect 2313 24787 2379 24790
rect 6545 24787 6611 24790
rect 8201 24850 8267 24853
rect 14549 24850 14615 24853
rect 8201 24848 14615 24850
rect 8201 24792 8206 24848
rect 8262 24792 14554 24848
rect 14610 24792 14615 24848
rect 8201 24790 14615 24792
rect 8201 24787 8267 24790
rect 14549 24787 14615 24790
rect 16573 24850 16639 24853
rect 16757 24850 16823 24853
rect 16573 24848 16823 24850
rect 16573 24792 16578 24848
rect 16634 24792 16762 24848
rect 16818 24792 16823 24848
rect 16573 24790 16823 24792
rect 16573 24787 16639 24790
rect 16757 24787 16823 24790
rect 3693 24714 3759 24717
rect 4613 24714 4679 24717
rect 1350 24654 3434 24714
rect 3374 24578 3434 24654
rect 3693 24712 4679 24714
rect 3693 24656 3698 24712
rect 3754 24656 4618 24712
rect 4674 24656 4679 24712
rect 3693 24654 4679 24656
rect 3693 24651 3759 24654
rect 4613 24651 4679 24654
rect 6177 24714 6243 24717
rect 8109 24714 8175 24717
rect 11789 24714 11855 24717
rect 6177 24712 8175 24714
rect 6177 24656 6182 24712
rect 6238 24656 8114 24712
rect 8170 24656 8175 24712
rect 6177 24654 8175 24656
rect 6177 24651 6243 24654
rect 8109 24651 8175 24654
rect 8342 24712 11855 24714
rect 8342 24656 11794 24712
rect 11850 24656 11855 24712
rect 8342 24654 11855 24656
rect 4061 24578 4127 24581
rect 3374 24576 4127 24578
rect 3374 24520 4066 24576
rect 4122 24520 4127 24576
rect 3374 24518 4127 24520
rect 4061 24515 4127 24518
rect 3049 24442 3115 24445
rect 8017 24442 8083 24445
rect 8342 24442 8402 24654
rect 11789 24651 11855 24654
rect 15653 24578 15719 24581
rect 17401 24578 17467 24581
rect 15653 24576 17467 24578
rect 15653 24520 15658 24576
rect 15714 24520 17406 24576
rect 17462 24520 17467 24576
rect 15653 24518 17467 24520
rect 15653 24515 15719 24518
rect 17401 24515 17467 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 3049 24440 8402 24442
rect 3049 24384 3054 24440
rect 3110 24384 8022 24440
rect 8078 24384 8402 24440
rect 3049 24382 8402 24384
rect 17309 24442 17375 24445
rect 19057 24442 19123 24445
rect 17309 24440 19123 24442
rect 17309 24384 17314 24440
rect 17370 24384 19062 24440
rect 19118 24384 19123 24440
rect 17309 24382 19123 24384
rect 3049 24379 3115 24382
rect 8017 24379 8083 24382
rect 17309 24379 17375 24382
rect 19057 24379 19123 24382
rect 21817 24442 21883 24445
rect 23657 24442 23723 24445
rect 21817 24440 23723 24442
rect 21817 24384 21822 24440
rect 21878 24384 23662 24440
rect 23718 24384 23723 24440
rect 21817 24382 23723 24384
rect 21817 24379 21883 24382
rect 23657 24379 23723 24382
rect 0 24306 480 24336
rect 3417 24306 3483 24309
rect 0 24304 3483 24306
rect 0 24248 3422 24304
rect 3478 24248 3483 24304
rect 0 24246 3483 24248
rect 0 24216 480 24246
rect 3417 24243 3483 24246
rect 4429 24306 4495 24309
rect 15561 24306 15627 24309
rect 4429 24304 15627 24306
rect 4429 24248 4434 24304
rect 4490 24248 15566 24304
rect 15622 24248 15627 24304
rect 4429 24246 15627 24248
rect 4429 24243 4495 24246
rect 15561 24243 15627 24246
rect 3233 24170 3299 24173
rect 7005 24170 7071 24173
rect 3233 24168 7071 24170
rect 3233 24112 3238 24168
rect 3294 24112 7010 24168
rect 7066 24112 7071 24168
rect 3233 24110 7071 24112
rect 3233 24107 3299 24110
rect 7005 24107 7071 24110
rect 18413 24170 18479 24173
rect 20805 24170 20871 24173
rect 18413 24168 20871 24170
rect 18413 24112 18418 24168
rect 18474 24112 20810 24168
rect 20866 24112 20871 24168
rect 18413 24110 20871 24112
rect 18413 24107 18479 24110
rect 20805 24107 20871 24110
rect 20621 24034 20687 24037
rect 21909 24034 21975 24037
rect 20621 24032 21975 24034
rect 20621 23976 20626 24032
rect 20682 23976 21914 24032
rect 21970 23976 21975 24032
rect 20621 23974 21975 23976
rect 20621 23971 20687 23974
rect 21909 23971 21975 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 6453 23898 6519 23901
rect 9673 23898 9739 23901
rect 6453 23896 9739 23898
rect 6453 23840 6458 23896
rect 6514 23840 9678 23896
rect 9734 23840 9739 23896
rect 6453 23838 9739 23840
rect 6453 23835 6519 23838
rect 9673 23835 9739 23838
rect 16481 23898 16547 23901
rect 17953 23898 18019 23901
rect 16481 23896 18019 23898
rect 16481 23840 16486 23896
rect 16542 23840 17958 23896
rect 18014 23840 18019 23896
rect 16481 23838 18019 23840
rect 16481 23835 16547 23838
rect 17953 23835 18019 23838
rect 19517 23898 19583 23901
rect 21357 23898 21423 23901
rect 19517 23896 21423 23898
rect 19517 23840 19522 23896
rect 19578 23840 21362 23896
rect 21418 23840 21423 23896
rect 19517 23838 21423 23840
rect 19517 23835 19583 23838
rect 21357 23835 21423 23838
rect 21725 23898 21791 23901
rect 23105 23898 23171 23901
rect 21725 23896 23171 23898
rect 21725 23840 21730 23896
rect 21786 23840 23110 23896
rect 23166 23840 23171 23896
rect 21725 23838 23171 23840
rect 21725 23835 21791 23838
rect 23105 23835 23171 23838
rect 24945 23898 25011 23901
rect 27061 23898 27127 23901
rect 24945 23896 27127 23898
rect 24945 23840 24950 23896
rect 25006 23840 27066 23896
rect 27122 23840 27127 23896
rect 24945 23838 27127 23840
rect 24945 23835 25011 23838
rect 27061 23835 27127 23838
rect 0 23762 480 23792
rect 3325 23762 3391 23765
rect 0 23760 3391 23762
rect 0 23704 3330 23760
rect 3386 23704 3391 23760
rect 0 23702 3391 23704
rect 0 23672 480 23702
rect 3325 23699 3391 23702
rect 5441 23762 5507 23765
rect 10685 23762 10751 23765
rect 5441 23760 10751 23762
rect 5441 23704 5446 23760
rect 5502 23704 10690 23760
rect 10746 23704 10751 23760
rect 5441 23702 10751 23704
rect 5441 23699 5507 23702
rect 10685 23699 10751 23702
rect 1301 23626 1367 23629
rect 7097 23626 7163 23629
rect 1301 23624 7163 23626
rect 1301 23568 1306 23624
rect 1362 23568 7102 23624
rect 7158 23568 7163 23624
rect 1301 23566 7163 23568
rect 1301 23563 1367 23566
rect 7097 23563 7163 23566
rect 16389 23626 16455 23629
rect 18229 23626 18295 23629
rect 16389 23624 18295 23626
rect 16389 23568 16394 23624
rect 16450 23568 18234 23624
rect 18290 23568 18295 23624
rect 16389 23566 18295 23568
rect 16389 23563 16455 23566
rect 18229 23563 18295 23566
rect 16757 23490 16823 23493
rect 18505 23490 18571 23493
rect 16757 23488 18571 23490
rect 16757 23432 16762 23488
rect 16818 23432 18510 23488
rect 18566 23432 18571 23488
rect 16757 23430 18571 23432
rect 16757 23427 16823 23430
rect 18505 23427 18571 23430
rect 24025 23490 24091 23493
rect 25957 23490 26023 23493
rect 24025 23488 26023 23490
rect 24025 23432 24030 23488
rect 24086 23432 25962 23488
rect 26018 23432 26023 23488
rect 24025 23430 26023 23432
rect 24025 23427 24091 23430
rect 25957 23427 26023 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 1669 23354 1735 23357
rect 5073 23354 5139 23357
rect 1669 23352 5139 23354
rect 1669 23296 1674 23352
rect 1730 23296 5078 23352
rect 5134 23296 5139 23352
rect 1669 23294 5139 23296
rect 1669 23291 1735 23294
rect 5073 23291 5139 23294
rect 12249 23354 12315 23357
rect 15193 23354 15259 23357
rect 12249 23352 15259 23354
rect 12249 23296 12254 23352
rect 12310 23296 15198 23352
rect 15254 23296 15259 23352
rect 12249 23294 15259 23296
rect 12249 23291 12315 23294
rect 15193 23291 15259 23294
rect 22369 23354 22435 23357
rect 24301 23354 24367 23357
rect 22369 23352 24367 23354
rect 22369 23296 22374 23352
rect 22430 23296 24306 23352
rect 24362 23296 24367 23352
rect 22369 23294 24367 23296
rect 22369 23291 22435 23294
rect 24301 23291 24367 23294
rect 0 23218 480 23248
rect 1577 23218 1643 23221
rect 0 23216 1643 23218
rect 0 23160 1582 23216
rect 1638 23160 1643 23216
rect 0 23158 1643 23160
rect 0 23128 480 23158
rect 1577 23155 1643 23158
rect 2589 23218 2655 23221
rect 2773 23218 2839 23221
rect 2589 23216 2839 23218
rect 2589 23160 2594 23216
rect 2650 23160 2778 23216
rect 2834 23160 2839 23216
rect 2589 23158 2839 23160
rect 2589 23155 2655 23158
rect 2773 23155 2839 23158
rect 2957 23218 3023 23221
rect 5533 23218 5599 23221
rect 2957 23216 5599 23218
rect 2957 23160 2962 23216
rect 3018 23160 5538 23216
rect 5594 23160 5599 23216
rect 2957 23158 5599 23160
rect 2957 23155 3023 23158
rect 5533 23155 5599 23158
rect 2129 23082 2195 23085
rect 5993 23082 6059 23085
rect 2129 23080 6059 23082
rect 2129 23024 2134 23080
rect 2190 23024 5998 23080
rect 6054 23024 6059 23080
rect 2129 23022 6059 23024
rect 2129 23019 2195 23022
rect 5993 23019 6059 23022
rect 2773 22946 2839 22949
rect 3785 22946 3851 22949
rect 4613 22946 4679 22949
rect 2773 22944 4679 22946
rect 2773 22888 2778 22944
rect 2834 22888 3790 22944
rect 3846 22888 4618 22944
rect 4674 22888 4679 22944
rect 2773 22886 4679 22888
rect 2773 22883 2839 22886
rect 3785 22883 3851 22886
rect 4613 22883 4679 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 5625 22674 5691 22677
rect 9949 22674 10015 22677
rect 5625 22672 10015 22674
rect 5625 22616 5630 22672
rect 5686 22616 9954 22672
rect 10010 22616 10015 22672
rect 5625 22614 10015 22616
rect 5625 22611 5691 22614
rect 9949 22611 10015 22614
rect 0 22538 480 22568
rect 1577 22538 1643 22541
rect 0 22536 1643 22538
rect 0 22480 1582 22536
rect 1638 22480 1643 22536
rect 0 22478 1643 22480
rect 0 22448 480 22478
rect 1577 22475 1643 22478
rect 6361 22538 6427 22541
rect 12433 22538 12499 22541
rect 6361 22536 12499 22538
rect 6361 22480 6366 22536
rect 6422 22480 12438 22536
rect 12494 22480 12499 22536
rect 6361 22478 12499 22480
rect 6361 22475 6427 22478
rect 12433 22475 12499 22478
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 10041 22130 10107 22133
rect 16849 22130 16915 22133
rect 10041 22128 16915 22130
rect 10041 22072 10046 22128
rect 10102 22072 16854 22128
rect 16910 22072 16915 22128
rect 10041 22070 16915 22072
rect 10041 22067 10107 22070
rect 16849 22067 16915 22070
rect 0 21994 480 22024
rect 2865 21994 2931 21997
rect 0 21992 2931 21994
rect 0 21936 2870 21992
rect 2926 21936 2931 21992
rect 0 21934 2931 21936
rect 0 21904 480 21934
rect 2865 21931 2931 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 10133 21586 10199 21589
rect 13813 21586 13879 21589
rect 10133 21584 13879 21586
rect 10133 21528 10138 21584
rect 10194 21528 13818 21584
rect 13874 21528 13879 21584
rect 10133 21526 13879 21528
rect 10133 21523 10199 21526
rect 13813 21523 13879 21526
rect 0 21450 480 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 480 21390
rect 1577 21387 1643 21390
rect 5349 21450 5415 21453
rect 11605 21450 11671 21453
rect 5349 21448 11671 21450
rect 5349 21392 5354 21448
rect 5410 21392 11610 21448
rect 11666 21392 11671 21448
rect 5349 21390 11671 21392
rect 5349 21387 5415 21390
rect 11605 21387 11671 21390
rect 21081 21450 21147 21453
rect 22461 21450 22527 21453
rect 21081 21448 22527 21450
rect 21081 21392 21086 21448
rect 21142 21392 22466 21448
rect 22522 21392 22527 21448
rect 21081 21390 22527 21392
rect 21081 21387 21147 21390
rect 22461 21387 22527 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 3141 21178 3207 21181
rect 7649 21178 7715 21181
rect 3141 21176 7715 21178
rect 3141 21120 3146 21176
rect 3202 21120 7654 21176
rect 7710 21120 7715 21176
rect 3141 21118 7715 21120
rect 3141 21115 3207 21118
rect 7649 21115 7715 21118
rect 7649 21042 7715 21045
rect 11145 21042 11211 21045
rect 7649 21040 11211 21042
rect 7649 20984 7654 21040
rect 7710 20984 11150 21040
rect 11206 20984 11211 21040
rect 7649 20982 11211 20984
rect 7649 20979 7715 20982
rect 11145 20979 11211 20982
rect 0 20906 480 20936
rect 2681 20906 2747 20909
rect 0 20904 2747 20906
rect 0 20848 2686 20904
rect 2742 20848 2747 20904
rect 0 20846 2747 20848
rect 0 20816 480 20846
rect 2681 20843 2747 20846
rect 9397 20770 9463 20773
rect 13813 20770 13879 20773
rect 9397 20768 13879 20770
rect 9397 20712 9402 20768
rect 9458 20712 13818 20768
rect 13874 20712 13879 20768
rect 9397 20710 13879 20712
rect 9397 20707 9463 20710
rect 13813 20707 13879 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 8293 20634 8359 20637
rect 14365 20634 14431 20637
rect 8293 20632 14431 20634
rect 8293 20576 8298 20632
rect 8354 20576 14370 20632
rect 14426 20576 14431 20632
rect 8293 20574 14431 20576
rect 8293 20571 8359 20574
rect 14365 20571 14431 20574
rect 3601 20498 3667 20501
rect 7189 20498 7255 20501
rect 10409 20498 10475 20501
rect 13905 20498 13971 20501
rect 3601 20496 13971 20498
rect 3601 20440 3606 20496
rect 3662 20440 7194 20496
rect 7250 20440 10414 20496
rect 10470 20440 13910 20496
rect 13966 20440 13971 20496
rect 3601 20438 13971 20440
rect 3601 20435 3667 20438
rect 7189 20435 7255 20438
rect 10409 20435 10475 20438
rect 13905 20435 13971 20438
rect 0 20362 480 20392
rect 2957 20362 3023 20365
rect 0 20360 3023 20362
rect 0 20304 2962 20360
rect 3018 20304 3023 20360
rect 0 20302 3023 20304
rect 0 20272 480 20302
rect 2957 20299 3023 20302
rect 4889 20362 4955 20365
rect 11881 20362 11947 20365
rect 4889 20360 11947 20362
rect 4889 20304 4894 20360
rect 4950 20304 11886 20360
rect 11942 20304 11947 20360
rect 4889 20302 11947 20304
rect 4889 20299 4955 20302
rect 11881 20299 11947 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 8109 20090 8175 20093
rect 10041 20090 10107 20093
rect 8109 20088 10107 20090
rect 8109 20032 8114 20088
rect 8170 20032 10046 20088
rect 10102 20032 10107 20088
rect 8109 20030 10107 20032
rect 8109 20027 8175 20030
rect 10041 20027 10107 20030
rect 7925 19818 7991 19821
rect 9673 19818 9739 19821
rect 7925 19816 9739 19818
rect 7925 19760 7930 19816
rect 7986 19760 9678 19816
rect 9734 19760 9739 19816
rect 7925 19758 9739 19760
rect 7925 19755 7991 19758
rect 9673 19755 9739 19758
rect 0 19682 480 19712
rect 1577 19682 1643 19685
rect 0 19680 1643 19682
rect 0 19624 1582 19680
rect 1638 19624 1643 19680
rect 0 19622 1643 19624
rect 0 19592 480 19622
rect 1577 19619 1643 19622
rect 12065 19682 12131 19685
rect 12525 19682 12591 19685
rect 12065 19680 12591 19682
rect 12065 19624 12070 19680
rect 12126 19624 12530 19680
rect 12586 19624 12591 19680
rect 12065 19622 12591 19624
rect 12065 19619 12131 19622
rect 12525 19619 12591 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 9630 19486 13370 19546
rect 9630 19447 9690 19486
rect 9581 19442 9690 19447
rect 5073 19410 5139 19413
rect 7373 19410 7439 19413
rect 5073 19408 7439 19410
rect 5073 19352 5078 19408
rect 5134 19352 7378 19408
rect 7434 19352 7439 19408
rect 9581 19386 9586 19442
rect 9642 19386 9690 19442
rect 9581 19384 9690 19386
rect 13310 19410 13370 19486
rect 16573 19410 16639 19413
rect 13310 19408 16639 19410
rect 9581 19381 9647 19384
rect 5073 19350 7439 19352
rect 13310 19352 16578 19408
rect 16634 19352 16639 19408
rect 13310 19350 16639 19352
rect 5073 19347 5139 19350
rect 7373 19347 7439 19350
rect 16573 19347 16639 19350
rect 8109 19274 8175 19277
rect 13997 19274 14063 19277
rect 8109 19272 14063 19274
rect 8109 19216 8114 19272
rect 8170 19216 14002 19272
rect 14058 19216 14063 19272
rect 8109 19214 14063 19216
rect 8109 19211 8175 19214
rect 13997 19211 14063 19214
rect 14181 19274 14247 19277
rect 23657 19274 23723 19277
rect 14181 19272 23723 19274
rect 14181 19216 14186 19272
rect 14242 19216 23662 19272
rect 23718 19216 23723 19272
rect 14181 19214 23723 19216
rect 14181 19211 14247 19214
rect 23657 19211 23723 19214
rect 0 19138 480 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 480 19078
rect 1485 19075 1551 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 10685 19002 10751 19005
rect 15745 19002 15811 19005
rect 10685 19000 15811 19002
rect 10685 18944 10690 19000
rect 10746 18944 15750 19000
rect 15806 18944 15811 19000
rect 10685 18942 15811 18944
rect 10685 18939 10751 18942
rect 15745 18939 15811 18942
rect 7281 18866 7347 18869
rect 14733 18866 14799 18869
rect 7281 18864 14799 18866
rect 7281 18808 7286 18864
rect 7342 18808 14738 18864
rect 14794 18808 14799 18864
rect 7281 18806 14799 18808
rect 7281 18803 7347 18806
rect 14733 18803 14799 18806
rect 0 18594 480 18624
rect 2681 18594 2747 18597
rect 0 18592 2747 18594
rect 0 18536 2686 18592
rect 2742 18536 2747 18592
rect 0 18534 2747 18536
rect 0 18504 480 18534
rect 2681 18531 2747 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 16389 18186 16455 18189
rect 26509 18186 26575 18189
rect 16389 18184 26575 18186
rect 16389 18128 16394 18184
rect 16450 18128 26514 18184
rect 26570 18128 26575 18184
rect 16389 18126 26575 18128
rect 16389 18123 16455 18126
rect 26509 18123 26575 18126
rect 0 18050 480 18080
rect 2497 18050 2563 18053
rect 0 18048 2563 18050
rect 0 17992 2502 18048
rect 2558 17992 2563 18048
rect 0 17990 2563 17992
rect 0 17960 480 17990
rect 2497 17987 2563 17990
rect 3601 18050 3667 18053
rect 8293 18050 8359 18053
rect 3601 18048 8359 18050
rect 3601 17992 3606 18048
rect 3662 17992 8298 18048
rect 8354 17992 8359 18048
rect 3601 17990 8359 17992
rect 3601 17987 3667 17990
rect 8293 17987 8359 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3877 17914 3943 17917
rect 8477 17914 8543 17917
rect 3877 17912 8543 17914
rect 3877 17856 3882 17912
rect 3938 17856 8482 17912
rect 8538 17856 8543 17912
rect 3877 17854 8543 17856
rect 3877 17851 3943 17854
rect 8477 17851 8543 17854
rect 10961 17914 11027 17917
rect 18045 17914 18111 17917
rect 10961 17912 18111 17914
rect 10961 17856 10966 17912
rect 11022 17856 18050 17912
rect 18106 17856 18111 17912
rect 10961 17854 18111 17856
rect 10961 17851 11027 17854
rect 18045 17851 18111 17854
rect 5073 17778 5139 17781
rect 17861 17778 17927 17781
rect 5073 17776 17927 17778
rect 5073 17720 5078 17776
rect 5134 17720 17866 17776
rect 17922 17720 17927 17776
rect 5073 17718 17927 17720
rect 5073 17715 5139 17718
rect 17861 17715 17927 17718
rect 7465 17642 7531 17645
rect 5398 17640 7531 17642
rect 5398 17584 7470 17640
rect 7526 17584 7531 17640
rect 5398 17582 7531 17584
rect 0 17506 480 17536
rect 1393 17506 1459 17509
rect 0 17504 1459 17506
rect 0 17448 1398 17504
rect 1454 17448 1459 17504
rect 0 17446 1459 17448
rect 0 17416 480 17446
rect 1393 17443 1459 17446
rect 2589 17506 2655 17509
rect 2957 17506 3023 17509
rect 4521 17506 4587 17509
rect 5398 17506 5458 17582
rect 7465 17579 7531 17582
rect 8109 17642 8175 17645
rect 15377 17642 15443 17645
rect 8109 17640 15443 17642
rect 8109 17584 8114 17640
rect 8170 17584 15382 17640
rect 15438 17584 15443 17640
rect 8109 17582 15443 17584
rect 8109 17579 8175 17582
rect 15377 17579 15443 17582
rect 2589 17504 5458 17506
rect 2589 17448 2594 17504
rect 2650 17448 2962 17504
rect 3018 17448 4526 17504
rect 4582 17448 5458 17504
rect 2589 17446 5458 17448
rect 2589 17443 2655 17446
rect 2957 17443 3023 17446
rect 4521 17443 4587 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 4337 17234 4403 17237
rect 6126 17234 6132 17236
rect 4337 17232 6132 17234
rect 4337 17176 4342 17232
rect 4398 17176 6132 17232
rect 4337 17174 6132 17176
rect 4337 17171 4403 17174
rect 6126 17172 6132 17174
rect 6196 17172 6202 17236
rect 9673 17234 9739 17237
rect 18229 17234 18295 17237
rect 9673 17232 18295 17234
rect 9673 17176 9678 17232
rect 9734 17176 18234 17232
rect 18290 17176 18295 17232
rect 9673 17174 18295 17176
rect 9673 17171 9739 17174
rect 18229 17171 18295 17174
rect 1577 17098 1643 17101
rect 13445 17098 13511 17101
rect 1577 17096 13511 17098
rect 1577 17040 1582 17096
rect 1638 17040 13450 17096
rect 13506 17040 13511 17096
rect 1577 17038 13511 17040
rect 1577 17035 1643 17038
rect 13445 17035 13511 17038
rect 4153 16962 4219 16965
rect 4153 16960 10058 16962
rect 4153 16904 4158 16960
rect 4214 16904 10058 16960
rect 4153 16902 10058 16904
rect 4153 16899 4219 16902
rect 0 16826 480 16856
rect 9765 16826 9831 16829
rect 0 16824 9831 16826
rect 0 16768 9770 16824
rect 9826 16768 9831 16824
rect 0 16766 9831 16768
rect 0 16736 480 16766
rect 9765 16763 9831 16766
rect 4061 16690 4127 16693
rect 9765 16690 9831 16693
rect 4061 16688 9831 16690
rect 4061 16632 4066 16688
rect 4122 16632 9770 16688
rect 9826 16632 9831 16688
rect 4061 16630 9831 16632
rect 9998 16690 10058 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 11145 16690 11211 16693
rect 9998 16688 11211 16690
rect 9998 16632 11150 16688
rect 11206 16632 11211 16688
rect 9998 16630 11211 16632
rect 4061 16627 4127 16630
rect 9765 16627 9831 16630
rect 11145 16627 11211 16630
rect 14549 16690 14615 16693
rect 17953 16690 18019 16693
rect 14549 16688 18019 16690
rect 14549 16632 14554 16688
rect 14610 16632 17958 16688
rect 18014 16632 18019 16688
rect 14549 16630 18019 16632
rect 14549 16627 14615 16630
rect 17953 16627 18019 16630
rect 2129 16554 2195 16557
rect 8753 16554 8819 16557
rect 2129 16552 8819 16554
rect 2129 16496 2134 16552
rect 2190 16496 8758 16552
rect 8814 16496 8819 16552
rect 2129 16494 8819 16496
rect 2129 16491 2195 16494
rect 8753 16491 8819 16494
rect 6453 16418 6519 16421
rect 8477 16418 8543 16421
rect 6453 16416 8543 16418
rect 6453 16360 6458 16416
rect 6514 16360 8482 16416
rect 8538 16360 8543 16416
rect 6453 16358 8543 16360
rect 6453 16355 6519 16358
rect 8477 16355 8543 16358
rect 8753 16418 8819 16421
rect 12252 16418 12450 16452
rect 14733 16418 14799 16421
rect 8753 16416 14799 16418
rect 8753 16360 8758 16416
rect 8814 16392 14738 16416
rect 8814 16360 12312 16392
rect 8753 16358 12312 16360
rect 12390 16360 14738 16392
rect 14794 16360 14799 16416
rect 12390 16358 14799 16360
rect 8753 16355 8819 16358
rect 14733 16355 14799 16358
rect 5610 16352 5930 16353
rect 0 16282 480 16312
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 11237 16282 11303 16285
rect 0 16222 4906 16282
rect 0 16192 480 16222
rect 4846 16146 4906 16222
rect 5996 16280 11303 16282
rect 5996 16224 11242 16280
rect 11298 16224 11303 16280
rect 5996 16222 11303 16224
rect 5996 16146 6056 16222
rect 11237 16219 11303 16222
rect 4846 16086 6056 16146
rect 10777 16146 10843 16149
rect 19057 16146 19123 16149
rect 10777 16144 19123 16146
rect 10777 16088 10782 16144
rect 10838 16088 19062 16144
rect 19118 16088 19123 16144
rect 10777 16086 19123 16088
rect 10777 16083 10843 16086
rect 19057 16083 19123 16086
rect 5165 16010 5231 16013
rect 15285 16010 15351 16013
rect 5165 16008 15351 16010
rect 5165 15952 5170 16008
rect 5226 15952 15290 16008
rect 15346 15952 15351 16008
rect 5165 15950 15351 15952
rect 5165 15947 5231 15950
rect 15285 15947 15351 15950
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 19241 16010 19307 16013
rect 17972 16008 19307 16010
rect 17972 15952 19246 16008
rect 19302 15952 19307 16008
rect 17972 15950 19307 15952
rect 17972 15948 17978 15950
rect 19241 15947 19307 15950
rect 10277 15808 10597 15809
rect 0 15738 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 4061 15738 4127 15741
rect 0 15736 4127 15738
rect 0 15680 4066 15736
rect 4122 15680 4127 15736
rect 0 15678 4127 15680
rect 0 15648 480 15678
rect 4061 15675 4127 15678
rect 4521 15738 4587 15741
rect 6913 15738 6979 15741
rect 4521 15736 6979 15738
rect 4521 15680 4526 15736
rect 4582 15680 6918 15736
rect 6974 15680 6979 15736
rect 4521 15678 6979 15680
rect 4521 15675 4587 15678
rect 6913 15675 6979 15678
rect 4061 15602 4127 15605
rect 6637 15602 6703 15605
rect 4061 15600 6703 15602
rect 4061 15544 4066 15600
rect 4122 15544 6642 15600
rect 6698 15544 6703 15600
rect 4061 15542 6703 15544
rect 4061 15539 4127 15542
rect 6637 15539 6703 15542
rect 9489 15602 9555 15605
rect 18045 15602 18111 15605
rect 9489 15600 18111 15602
rect 9489 15544 9494 15600
rect 9550 15544 18050 15600
rect 18106 15544 18111 15600
rect 9489 15542 18111 15544
rect 9489 15539 9555 15542
rect 18045 15539 18111 15542
rect 3509 15466 3575 15469
rect 7189 15466 7255 15469
rect 3509 15464 7255 15466
rect 3509 15408 3514 15464
rect 3570 15408 7194 15464
rect 7250 15408 7255 15464
rect 3509 15406 7255 15408
rect 3509 15403 3575 15406
rect 7189 15403 7255 15406
rect 7741 15466 7807 15469
rect 11789 15466 11855 15469
rect 7741 15464 11855 15466
rect 7741 15408 7746 15464
rect 7802 15408 11794 15464
rect 11850 15408 11855 15464
rect 7741 15406 11855 15408
rect 7741 15403 7807 15406
rect 11789 15403 11855 15406
rect 12433 15466 12499 15469
rect 19425 15466 19491 15469
rect 12433 15464 19491 15466
rect 12433 15408 12438 15464
rect 12494 15408 19430 15464
rect 19486 15408 19491 15464
rect 12433 15406 19491 15408
rect 12433 15403 12499 15406
rect 19425 15403 19491 15406
rect 7281 15330 7347 15333
rect 11697 15330 11763 15333
rect 7281 15328 11763 15330
rect 7281 15272 7286 15328
rect 7342 15272 11702 15328
rect 11758 15272 11763 15328
rect 7281 15270 11763 15272
rect 7281 15267 7347 15270
rect 11697 15267 11763 15270
rect 5610 15264 5930 15265
rect 0 15194 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3969 15194 4035 15197
rect 0 15192 4035 15194
rect 0 15136 3974 15192
rect 4030 15136 4035 15192
rect 0 15134 4035 15136
rect 0 15104 480 15134
rect 3969 15131 4035 15134
rect 3509 15058 3575 15061
rect 11973 15058 12039 15061
rect 3509 15056 12039 15058
rect 3509 15000 3514 15056
rect 3570 15000 11978 15056
rect 12034 15000 12039 15056
rect 3509 14998 12039 15000
rect 3509 14995 3575 14998
rect 11973 14995 12039 14998
rect 3877 14922 3943 14925
rect 4521 14922 4587 14925
rect 8385 14922 8451 14925
rect 3877 14920 8451 14922
rect 3877 14864 3882 14920
rect 3938 14864 4526 14920
rect 4582 14864 8390 14920
rect 8446 14864 8451 14920
rect 3877 14862 8451 14864
rect 3877 14859 3943 14862
rect 4521 14859 4587 14862
rect 8385 14859 8451 14862
rect 16389 14922 16455 14925
rect 22553 14922 22619 14925
rect 16389 14920 22619 14922
rect 16389 14864 16394 14920
rect 16450 14864 22558 14920
rect 22614 14864 22619 14920
rect 16389 14862 22619 14864
rect 16389 14859 16455 14862
rect 22553 14859 22619 14862
rect 841 14786 907 14789
rect 1853 14786 1919 14789
rect 5073 14786 5139 14789
rect 841 14784 5139 14786
rect 841 14728 846 14784
rect 902 14728 1858 14784
rect 1914 14728 5078 14784
rect 5134 14728 5139 14784
rect 841 14726 5139 14728
rect 841 14723 907 14726
rect 1853 14723 1919 14726
rect 5073 14723 5139 14726
rect 5257 14786 5323 14789
rect 7465 14786 7531 14789
rect 5257 14784 7531 14786
rect 5257 14728 5262 14784
rect 5318 14728 7470 14784
rect 7526 14728 7531 14784
rect 5257 14726 7531 14728
rect 5257 14723 5323 14726
rect 7465 14723 7531 14726
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 480 14590
rect 1485 14587 1551 14590
rect 2773 14650 2839 14653
rect 4061 14650 4127 14653
rect 9029 14650 9095 14653
rect 2773 14648 9095 14650
rect 2773 14592 2778 14648
rect 2834 14592 4066 14648
rect 4122 14592 9034 14648
rect 9090 14592 9095 14648
rect 2773 14590 9095 14592
rect 2773 14587 2839 14590
rect 4061 14587 4127 14590
rect 9029 14587 9095 14590
rect 13629 14650 13695 14653
rect 18873 14650 18939 14653
rect 13629 14648 18939 14650
rect 13629 14592 13634 14648
rect 13690 14592 18878 14648
rect 18934 14592 18939 14648
rect 13629 14590 18939 14592
rect 13629 14587 13695 14590
rect 18873 14587 18939 14590
rect 3877 14514 3943 14517
rect 5993 14514 6059 14517
rect 3877 14512 6059 14514
rect 3877 14456 3882 14512
rect 3938 14456 5998 14512
rect 6054 14456 6059 14512
rect 3877 14454 6059 14456
rect 3877 14451 3943 14454
rect 5993 14451 6059 14454
rect 12249 14514 12315 14517
rect 15285 14514 15351 14517
rect 12249 14512 15351 14514
rect 12249 14456 12254 14512
rect 12310 14456 15290 14512
rect 15346 14456 15351 14512
rect 12249 14454 15351 14456
rect 12249 14451 12315 14454
rect 15285 14451 15351 14454
rect 3325 14378 3391 14381
rect 8017 14378 8083 14381
rect 3325 14376 8083 14378
rect 3325 14320 3330 14376
rect 3386 14320 8022 14376
rect 8078 14320 8083 14376
rect 3325 14318 8083 14320
rect 3325 14315 3391 14318
rect 8017 14315 8083 14318
rect 10041 14378 10107 14381
rect 13353 14378 13419 14381
rect 10041 14376 13419 14378
rect 10041 14320 10046 14376
rect 10102 14320 13358 14376
rect 13414 14320 13419 14376
rect 10041 14318 13419 14320
rect 10041 14315 10107 14318
rect 13353 14315 13419 14318
rect 2865 14242 2931 14245
rect 4153 14242 4219 14245
rect 2865 14240 4219 14242
rect 2865 14184 2870 14240
rect 2926 14184 4158 14240
rect 4214 14184 4219 14240
rect 2865 14182 4219 14184
rect 2865 14179 2931 14182
rect 4153 14179 4219 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 1761 14106 1827 14109
rect 3049 14106 3115 14109
rect 1761 14104 3115 14106
rect 1761 14048 1766 14104
rect 1822 14048 3054 14104
rect 3110 14048 3115 14104
rect 1761 14046 3115 14048
rect 1761 14043 1827 14046
rect 3049 14043 3115 14046
rect 0 13970 480 14000
rect 5533 13970 5599 13973
rect 11145 13970 11211 13973
rect 13905 13970 13971 13973
rect 0 13968 5599 13970
rect 0 13912 5538 13968
rect 5594 13912 5599 13968
rect 0 13910 5599 13912
rect 0 13880 480 13910
rect 5533 13907 5599 13910
rect 6134 13968 13971 13970
rect 6134 13912 11150 13968
rect 11206 13912 13910 13968
rect 13966 13912 13971 13968
rect 6134 13910 13971 13912
rect 3601 13834 3667 13837
rect 6134 13834 6194 13910
rect 11145 13907 11211 13910
rect 13905 13907 13971 13910
rect 3601 13832 6194 13834
rect 3601 13776 3606 13832
rect 3662 13776 6194 13832
rect 3601 13774 6194 13776
rect 6269 13834 6335 13837
rect 8569 13834 8635 13837
rect 6269 13832 8635 13834
rect 6269 13776 6274 13832
rect 6330 13776 8574 13832
rect 8630 13776 8635 13832
rect 6269 13774 8635 13776
rect 3601 13771 3667 13774
rect 6269 13771 6335 13774
rect 8569 13771 8635 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3509 13562 3575 13565
rect 9397 13562 9463 13565
rect 10041 13562 10107 13565
rect 3509 13560 10107 13562
rect 3509 13504 3514 13560
rect 3570 13504 9402 13560
rect 9458 13504 10046 13560
rect 10102 13504 10107 13560
rect 3509 13502 10107 13504
rect 3509 13499 3575 13502
rect 9397 13499 9463 13502
rect 10041 13499 10107 13502
rect 0 13426 480 13456
rect 5165 13426 5231 13429
rect 20897 13426 20963 13429
rect 0 13366 1410 13426
rect 0 13336 480 13366
rect 1350 13290 1410 13366
rect 5165 13424 20963 13426
rect 5165 13368 5170 13424
rect 5226 13368 20902 13424
rect 20958 13368 20963 13424
rect 5165 13366 20963 13368
rect 5165 13363 5231 13366
rect 20897 13363 20963 13366
rect 7649 13290 7715 13293
rect 1350 13288 7715 13290
rect 1350 13232 7654 13288
rect 7710 13232 7715 13288
rect 1350 13230 7715 13232
rect 7649 13227 7715 13230
rect 14181 13290 14247 13293
rect 19425 13290 19491 13293
rect 14181 13288 19491 13290
rect 14181 13232 14186 13288
rect 14242 13232 19430 13288
rect 19486 13232 19491 13288
rect 14181 13230 19491 13232
rect 14181 13227 14247 13230
rect 19425 13227 19491 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 0 12882 480 12912
rect 4245 12882 4311 12885
rect 0 12880 4311 12882
rect 0 12824 4250 12880
rect 4306 12824 4311 12880
rect 0 12822 4311 12824
rect 0 12792 480 12822
rect 4245 12819 4311 12822
rect 5809 12882 5875 12885
rect 13813 12882 13879 12885
rect 5809 12880 13879 12882
rect 5809 12824 5814 12880
rect 5870 12824 13818 12880
rect 13874 12824 13879 12880
rect 5809 12822 13879 12824
rect 5809 12819 5875 12822
rect 13813 12819 13879 12822
rect 15101 12882 15167 12885
rect 16021 12882 16087 12885
rect 15101 12880 16087 12882
rect 15101 12824 15106 12880
rect 15162 12824 16026 12880
rect 16082 12824 16087 12880
rect 15101 12822 16087 12824
rect 15101 12819 15167 12822
rect 16021 12819 16087 12822
rect 4061 12746 4127 12749
rect 6085 12746 6151 12749
rect 10777 12746 10843 12749
rect 26233 12746 26299 12749
rect 4061 12744 6151 12746
rect 4061 12688 4066 12744
rect 4122 12688 6090 12744
rect 6146 12688 6151 12744
rect 4061 12686 6151 12688
rect 4061 12683 4127 12686
rect 6085 12683 6151 12686
rect 6502 12744 26299 12746
rect 6502 12688 10782 12744
rect 10838 12688 26238 12744
rect 26294 12688 26299 12744
rect 6502 12686 26299 12688
rect 3233 12610 3299 12613
rect 4981 12610 5047 12613
rect 3233 12608 5047 12610
rect 3233 12552 3238 12608
rect 3294 12552 4986 12608
rect 5042 12552 5047 12608
rect 3233 12550 5047 12552
rect 3233 12547 3299 12550
rect 4981 12547 5047 12550
rect 5257 12610 5323 12613
rect 5625 12610 5691 12613
rect 6502 12610 6562 12686
rect 10777 12683 10843 12686
rect 26233 12683 26299 12686
rect 5257 12608 6562 12610
rect 5257 12552 5262 12608
rect 5318 12552 5630 12608
rect 5686 12552 6562 12608
rect 5257 12550 6562 12552
rect 5257 12547 5323 12550
rect 5625 12547 5691 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 14825 12474 14891 12477
rect 15837 12474 15903 12477
rect 16573 12474 16639 12477
rect 14825 12472 16639 12474
rect 14825 12416 14830 12472
rect 14886 12416 15842 12472
rect 15898 12416 16578 12472
rect 16634 12416 16639 12472
rect 14825 12414 16639 12416
rect 14825 12411 14891 12414
rect 15837 12411 15903 12414
rect 16573 12411 16639 12414
rect 0 12338 480 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 480 12278
rect 1577 12275 1643 12278
rect 11237 12338 11303 12341
rect 21173 12338 21239 12341
rect 11237 12336 21239 12338
rect 11237 12280 11242 12336
rect 11298 12280 21178 12336
rect 21234 12280 21239 12336
rect 11237 12278 21239 12280
rect 11237 12275 11303 12278
rect 21173 12275 21239 12278
rect 22001 12338 22067 12341
rect 24209 12338 24275 12341
rect 22001 12336 24275 12338
rect 22001 12280 22006 12336
rect 22062 12280 24214 12336
rect 24270 12280 24275 12336
rect 22001 12278 24275 12280
rect 22001 12275 22067 12278
rect 24209 12275 24275 12278
rect 1761 12202 1827 12205
rect 13813 12202 13879 12205
rect 1761 12200 13879 12202
rect 1761 12144 1766 12200
rect 1822 12144 13818 12200
rect 13874 12144 13879 12200
rect 1761 12142 13879 12144
rect 1761 12139 1827 12142
rect 13813 12139 13879 12142
rect 13997 12202 14063 12205
rect 17953 12202 18019 12205
rect 13997 12200 18019 12202
rect 13997 12144 14002 12200
rect 14058 12144 17958 12200
rect 18014 12144 18019 12200
rect 13997 12142 18019 12144
rect 13997 12139 14063 12142
rect 17953 12139 18019 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 22277 11930 22343 11933
rect 17910 11928 22343 11930
rect 17910 11872 22282 11928
rect 22338 11872 22343 11928
rect 17910 11870 22343 11872
rect 0 11794 480 11824
rect 6177 11794 6243 11797
rect 0 11792 6243 11794
rect 0 11736 6182 11792
rect 6238 11736 6243 11792
rect 0 11734 6243 11736
rect 0 11704 480 11734
rect 6177 11731 6243 11734
rect 13629 11794 13695 11797
rect 17910 11794 17970 11870
rect 22277 11867 22343 11870
rect 13629 11792 17970 11794
rect 13629 11736 13634 11792
rect 13690 11736 17970 11792
rect 13629 11734 17970 11736
rect 13629 11731 13695 11734
rect 7465 11658 7531 11661
rect 2638 11656 7531 11658
rect 2638 11600 7470 11656
rect 7526 11600 7531 11656
rect 2638 11598 7531 11600
rect 0 11114 480 11144
rect 2405 11114 2471 11117
rect 2638 11114 2698 11598
rect 7465 11595 7531 11598
rect 7925 11658 7991 11661
rect 17769 11658 17835 11661
rect 19517 11658 19583 11661
rect 7925 11656 16636 11658
rect 7925 11600 7930 11656
rect 7986 11600 16636 11656
rect 7925 11598 16636 11600
rect 7925 11595 7991 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 16576 11250 16636 11598
rect 17769 11656 19583 11658
rect 17769 11600 17774 11656
rect 17830 11600 19522 11656
rect 19578 11600 19583 11656
rect 17769 11598 19583 11600
rect 17769 11595 17835 11598
rect 19517 11595 19583 11598
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 20805 11250 20871 11253
rect 16576 11248 20871 11250
rect 16576 11192 20810 11248
rect 20866 11192 20871 11248
rect 16576 11190 20871 11192
rect 20805 11187 20871 11190
rect 3693 11114 3759 11117
rect 0 11054 2330 11114
rect 0 11024 480 11054
rect 2270 10978 2330 11054
rect 2405 11112 2698 11114
rect 2405 11056 2410 11112
rect 2466 11056 2698 11112
rect 2405 11054 2698 11056
rect 2822 11112 3759 11114
rect 2822 11056 3698 11112
rect 3754 11056 3759 11112
rect 2822 11054 3759 11056
rect 2405 11051 2471 11054
rect 2822 10978 2882 11054
rect 3693 11051 3759 11054
rect 13353 11114 13419 11117
rect 22001 11114 22067 11117
rect 13353 11112 22067 11114
rect 13353 11056 13358 11112
rect 13414 11056 22006 11112
rect 22062 11056 22067 11112
rect 13353 11054 22067 11056
rect 13353 11051 13419 11054
rect 22001 11051 22067 11054
rect 2270 10918 2882 10978
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 4061 10706 4127 10709
rect 16757 10706 16823 10709
rect 4061 10704 16823 10706
rect 4061 10648 4066 10704
rect 4122 10648 16762 10704
rect 16818 10648 16823 10704
rect 4061 10646 16823 10648
rect 4061 10643 4127 10646
rect 16757 10643 16823 10646
rect 0 10570 480 10600
rect 1853 10570 1919 10573
rect 0 10568 1919 10570
rect 0 10512 1858 10568
rect 1914 10512 1919 10568
rect 0 10510 1919 10512
rect 0 10480 480 10510
rect 1853 10507 1919 10510
rect 3785 10434 3851 10437
rect 6545 10434 6611 10437
rect 3785 10432 6611 10434
rect 3785 10376 3790 10432
rect 3846 10376 6550 10432
rect 6606 10376 6611 10432
rect 3785 10374 6611 10376
rect 3785 10371 3851 10374
rect 6545 10371 6611 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 7649 10162 7715 10165
rect 16389 10162 16455 10165
rect 7649 10160 16455 10162
rect 7649 10104 7654 10160
rect 7710 10104 16394 10160
rect 16450 10104 16455 10160
rect 7649 10102 16455 10104
rect 7649 10099 7715 10102
rect 16389 10099 16455 10102
rect 0 10026 480 10056
rect 4521 10026 4587 10029
rect 0 10024 4587 10026
rect 0 9968 4526 10024
rect 4582 9968 4587 10024
rect 0 9966 4587 9968
rect 0 9936 480 9966
rect 4521 9963 4587 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 2313 9618 2379 9621
rect 7005 9618 7071 9621
rect 2313 9616 7071 9618
rect 2313 9560 2318 9616
rect 2374 9560 7010 9616
rect 7066 9560 7071 9616
rect 2313 9558 7071 9560
rect 2313 9555 2379 9558
rect 7005 9555 7071 9558
rect 9673 9618 9739 9621
rect 16941 9618 17007 9621
rect 9673 9616 17007 9618
rect 9673 9560 9678 9616
rect 9734 9560 16946 9616
rect 17002 9560 17007 9616
rect 9673 9558 17007 9560
rect 9673 9555 9739 9558
rect 16941 9555 17007 9558
rect 0 9482 480 9512
rect 6361 9482 6427 9485
rect 0 9480 6427 9482
rect 0 9424 6366 9480
rect 6422 9424 6427 9480
rect 0 9422 6427 9424
rect 0 9392 480 9422
rect 6361 9419 6427 9422
rect 12433 9482 12499 9485
rect 18045 9482 18111 9485
rect 12433 9480 18111 9482
rect 12433 9424 12438 9480
rect 12494 9424 18050 9480
rect 18106 9424 18111 9480
rect 12433 9422 18111 9424
rect 12433 9419 12499 9422
rect 18045 9419 18111 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2037 9210 2103 9213
rect 9949 9210 10015 9213
rect 2037 9208 10015 9210
rect 2037 9152 2042 9208
rect 2098 9152 9954 9208
rect 10010 9152 10015 9208
rect 2037 9150 10015 9152
rect 2037 9147 2103 9150
rect 9949 9147 10015 9150
rect 10777 9210 10843 9213
rect 12985 9210 13051 9213
rect 10777 9208 13051 9210
rect 10777 9152 10782 9208
rect 10838 9152 12990 9208
rect 13046 9152 13051 9208
rect 10777 9150 13051 9152
rect 10777 9147 10843 9150
rect 12985 9147 13051 9150
rect 0 8938 480 8968
rect 7741 8938 7807 8941
rect 0 8936 7807 8938
rect 0 8880 7746 8936
rect 7802 8880 7807 8936
rect 0 8878 7807 8880
rect 0 8848 480 8878
rect 7741 8875 7807 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 1669 8530 1735 8533
rect 9857 8530 9923 8533
rect 1669 8528 9923 8530
rect 1669 8472 1674 8528
rect 1730 8472 9862 8528
rect 9918 8472 9923 8528
rect 1669 8470 9923 8472
rect 1669 8467 1735 8470
rect 9857 8467 9923 8470
rect 10593 8394 10659 8397
rect 4846 8392 10659 8394
rect 4846 8336 10598 8392
rect 10654 8336 10659 8392
rect 4846 8334 10659 8336
rect 0 8258 480 8288
rect 4846 8258 4906 8334
rect 10593 8331 10659 8334
rect 0 8198 4906 8258
rect 0 8168 480 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 4061 7986 4127 7989
rect 15837 7986 15903 7989
rect 4061 7984 15903 7986
rect 4061 7928 4066 7984
rect 4122 7928 15842 7984
rect 15898 7928 15903 7984
rect 4061 7926 15903 7928
rect 4061 7923 4127 7926
rect 15837 7923 15903 7926
rect 9622 7788 9628 7852
rect 9692 7850 9698 7852
rect 12525 7850 12591 7853
rect 9692 7848 12591 7850
rect 9692 7792 12530 7848
rect 12586 7792 12591 7848
rect 9692 7790 12591 7792
rect 9692 7788 9698 7790
rect 12525 7787 12591 7790
rect 0 7714 480 7744
rect 0 7654 4906 7714
rect 0 7624 480 7654
rect 4846 7442 4906 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 13445 7442 13511 7445
rect 4846 7440 13511 7442
rect 4846 7384 13450 7440
rect 13506 7384 13511 7440
rect 4846 7382 13511 7384
rect 13445 7379 13511 7382
rect 0 7170 480 7200
rect 4061 7170 4127 7173
rect 0 7168 4127 7170
rect 0 7112 4066 7168
rect 4122 7112 4127 7168
rect 0 7110 4127 7112
rect 0 7080 480 7110
rect 4061 7107 4127 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 4061 6898 4127 6901
rect 9489 6898 9555 6901
rect 4061 6896 9555 6898
rect 4061 6840 4066 6896
rect 4122 6840 9494 6896
rect 9550 6840 9555 6896
rect 4061 6838 9555 6840
rect 4061 6835 4127 6838
rect 9489 6835 9555 6838
rect 3877 6762 3943 6765
rect 11513 6762 11579 6765
rect 3877 6760 11579 6762
rect 3877 6704 3882 6760
rect 3938 6704 11518 6760
rect 11574 6704 11579 6760
rect 3877 6702 11579 6704
rect 3877 6699 3943 6702
rect 11513 6699 11579 6702
rect 0 6626 480 6656
rect 4797 6626 4863 6629
rect 0 6624 4863 6626
rect 0 6568 4802 6624
rect 4858 6568 4863 6624
rect 0 6566 4863 6568
rect 0 6536 480 6566
rect 4797 6563 4863 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 9489 6354 9555 6357
rect 9622 6354 9628 6356
rect 9489 6352 9628 6354
rect 9489 6296 9494 6352
rect 9550 6296 9628 6352
rect 9489 6294 9628 6296
rect 9489 6291 9555 6294
rect 9622 6292 9628 6294
rect 9692 6292 9698 6356
rect 11421 6218 11487 6221
rect 4662 6216 11487 6218
rect 4662 6160 11426 6216
rect 11482 6160 11487 6216
rect 4662 6158 11487 6160
rect 0 6082 480 6112
rect 4662 6082 4722 6158
rect 11421 6155 11487 6158
rect 0 6022 4722 6082
rect 0 5992 480 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 5610 5472 5930 5473
rect 0 5402 480 5432
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 3969 5402 4035 5405
rect 0 5400 4035 5402
rect 0 5344 3974 5400
rect 4030 5344 4035 5400
rect 0 5342 4035 5344
rect 0 5312 480 5342
rect 3969 5339 4035 5342
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3785 4858 3851 4861
rect 0 4856 3851 4858
rect 0 4800 3790 4856
rect 3846 4800 3851 4856
rect 0 4798 3851 4800
rect 0 4768 480 4798
rect 3785 4795 3851 4798
rect 5610 4384 5930 4385
rect 0 4314 480 4344
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3877 3770 3943 3773
rect 0 3768 3943 3770
rect 0 3712 3882 3768
rect 3938 3712 3943 3768
rect 0 3710 3943 3712
rect 0 3680 480 3710
rect 3877 3707 3943 3710
rect 12065 3498 12131 3501
rect 23197 3498 23263 3501
rect 12065 3496 23263 3498
rect 12065 3440 12070 3496
rect 12126 3440 23202 3496
rect 23258 3440 23263 3496
rect 12065 3438 23263 3440
rect 12065 3435 12131 3438
rect 23197 3435 23263 3438
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 0 3166 3066 3226
rect 0 3136 480 3166
rect 3006 2954 3066 3166
rect 14825 2954 14891 2957
rect 3006 2952 14891 2954
rect 3006 2896 14830 2952
rect 14886 2896 14891 2952
rect 3006 2894 14891 2896
rect 14825 2891 14891 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2546 480 2576
rect 15929 2546 15995 2549
rect 0 2544 15995 2546
rect 0 2488 15934 2544
rect 15990 2488 15995 2544
rect 0 2486 15995 2488
rect 0 2456 480 2486
rect 15929 2483 15995 2486
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 0 2002 480 2032
rect 0 1942 1594 2002
rect 0 1912 480 1942
rect 1534 1730 1594 1942
rect 13537 1730 13603 1733
rect 1534 1728 13603 1730
rect 1534 1672 13542 1728
rect 13598 1672 13603 1728
rect 1534 1670 13603 1672
rect 13537 1667 13603 1670
rect 0 1458 480 1488
rect 11145 1458 11211 1461
rect 0 1456 11211 1458
rect 0 1400 11150 1456
rect 11206 1400 11211 1456
rect 0 1398 11211 1400
rect 0 1368 480 1398
rect 11145 1395 11211 1398
rect 0 914 480 944
rect 10041 914 10107 917
rect 0 912 10107 914
rect 0 856 10046 912
rect 10102 856 10107 912
rect 0 854 10107 856
rect 0 824 480 854
rect 10041 851 10107 854
rect 0 370 480 400
rect 2957 370 3023 373
rect 0 368 3023 370
rect 0 312 2962 368
rect 3018 312 3023 368
rect 0 310 3023 312
rect 0 280 480 310
rect 2957 307 3023 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 6132 17172 6196 17236
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 17908 15948 17972 16012
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 9628 7788 9692 7852
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 9628 6292 9692 6356
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 6131 17236 6197 17237
rect 6131 17172 6132 17236
rect 6196 17172 6197 17236
rect 6131 17171 6197 17172
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 6134 16098 6194 17171
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 9630 6357 9690 7787
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 9627 6356 9693 6357
rect 9627 6292 9628 6356
rect 9692 6292 9693 6356
rect 9627 6291 9693 6292
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 6046 15862 6282 16098
rect 17822 16012 18058 16098
rect 17822 15948 17908 16012
rect 17908 15948 17972 16012
rect 17972 15948 18058 16012
rect 17822 15862 18058 15948
<< metal5 >>
rect 6004 16098 18100 16140
rect 6004 15862 6046 16098
rect 6282 15862 17822 16098
rect 18058 15862 18100 16098
rect 6004 15820 18100 15862
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_112
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_124
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_136
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_148
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_119
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_97
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 1786 592
use scs8hd_conb_1  _038_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12696 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_124
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_17.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_48
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _036_
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_70
timestamp 1586364061
transform 1 0 7544 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_97
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_14.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_101
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_buf_1  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_17
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_26
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_62
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_66
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_70
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_116
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 130 592
use scs8hd_conb_1  _039_
timestamp 1586364061
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_149
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_162
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 314 592
use scs8hd_buf_1  mux_left_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_39
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_conb_1  _054_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_50
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7636 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_28.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_30.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_conb_1  _037_
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_131
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_137
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 1786 592
use scs8hd_buf_1  mux_top_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_164
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_187
timestamp 1586364061
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_203
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_215
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_243
timestamp 1586364061
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_89
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_146
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 18308 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_181
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_219
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_243
timestamp 1586364061
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _053_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_conb_1  _044_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_52
timestamp 1586364061
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_26.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_60
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _046_
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_98
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_30.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_30.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_30.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_146
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_150
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_167
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_207
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_30
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_40
timestamp 1586364061
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _045_
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_28.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _047_
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 590 592
use scs8hd_conb_1  _048_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_28.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_203
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_28.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_225
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_229
timestamp 1586364061
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_241
timestamp 1586364061
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2760 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_16
timestamp 1586364061
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _086_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_24
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_71
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_28.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_28.mux_l2_in_0_
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_30.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_32.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_177
timestamp 1586364061
transform 1 0 17388 0 -1 12512
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_200
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_212
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  mux_top_track_30.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21804 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_223
timestamp 1586364061
transform 1 0 21620 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_228
timestamp 1586364061
transform 1 0 22080 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_240
timestamp 1586364061
transform 1 0 23184 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_264
timestamp 1586364061
transform 1 0 25392 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_272
timestamp 1586364061
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _087_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_20_28
timestamp 1586364061
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_24
timestamp 1586364061
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_20
timestamp 1586364061
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3128 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_48
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 5888 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_26.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  _085_
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_26.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_85
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 866 592
use scs8hd_conb_1  _035_
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11776 0 -1 13600
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_135
timestamp 1586364061
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_147
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_139
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  mux_top_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_163
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_176
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 774 592
use scs8hd_conb_1  _040_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_203
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_32.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22264 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_32.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_229
timestamp 1586364061
transform 1 0 22172 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_233
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_237
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_254
timestamp 1586364061
transform 1 0 24472 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_266
timestamp 1586364061
transform 1 0 25576 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7544 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _043_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_120
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_133
timestamp 1586364061
transform 1 0 13340 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_163
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_167
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_conb_1  _052_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_46
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_50
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_73
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_77
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use scs8hd_conb_1  _041_
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_131
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_135
timestamp 1586364061
transform 1 0 13524 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 314 592
use scs8hd_conb_1  _049_
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_34.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_170
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_181
timestamp 1586364061
transform 1 0 17756 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_193
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_205
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_213
timestamp 1586364061
transform 1 0 20700 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _078_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 1786 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_38
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_buf_2  _084_
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_42
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_50
timestamp 1586364061
transform 1 0 5704 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_54
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_85
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use scs8hd_conb_1  _042_
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_34.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_34.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_202
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_206
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_214
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_229
timestamp 1586364061
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4600 0 -1 15776
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_36
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_57
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_61
timestamp 1586364061
transform 1 0 6716 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_78
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_82
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10396 0 -1 15776
box -38 -48 1786 592
use scs8hd_mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_120
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_125
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_146
timestamp 1586364061
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_157
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_34.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 1786 592
use scs8hd_decap_12  FILLER_24_184
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_196
timestamp 1586364061
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _096_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_208
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_231
timestamp 1586364061
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_243
timestamp 1586364061
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_255
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_267
timestamp 1586364061
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_77
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 314 592
use scs8hd_conb_1  _034_
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_83
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_87
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _080_
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_100
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_104
timestamp 1586364061
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_107
timestamp 1586364061
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_116
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _050_
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_172
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_176
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use scs8hd_buf_1  mux_left_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_202
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_226
timestamp 1586364061
transform 1 0 21896 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_238
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _075_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _074_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_14
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_14
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_11
timestamp 1586364061
transform 1 0 2116 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _077_
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use scs8hd_buf_2  _076_
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_23
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_24
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_48
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_44
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5336 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_50
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_54
timestamp 1586364061
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use scs8hd_mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_67
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 866 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_84
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_97
timestamp 1586364061
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_90
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  _081_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_38.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use scs8hd_mux2_1  mux_top_track_36.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_147
timestamp 1586364061
transform 1 0 14628 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_143
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_36.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_158
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14996 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_top_track_36.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_162
timestamp 1586364061
transform 1 0 16008 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 774 592
use scs8hd_buf_1  mux_left_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_187
timestamp 1586364061
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_191
timestamp 1586364061
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_203
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_215
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_239
timestamp 1586364061
transform 1 0 23092 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  FILLER_28_9
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_21
timestamp 1586364061
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_25
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_buf_2  _079_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_85
timestamp 1586364061
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_27.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_136
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_1  mux_top_track_36.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_buf_1  mux_top_track_36.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_36.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 590 592
use scs8hd_buf_1  mux_left_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_174
timestamp 1586364061
transform 1 0 17112 0 -1 17952
box -38 -48 774 592
use scs8hd_conb_1  _066_
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_185
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_197
timestamp 1586364061
transform 1 0 19228 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_209
timestamp 1586364061
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 1786 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_8
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_31
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_48
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_52
timestamp 1586364061
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_56
timestamp 1586364061
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9292 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_85
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_100
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _056_
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_38.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_38.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use scs8hd_buf_2  _089_
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_160
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_180
timestamp 1586364061
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_16
timestamp 1586364061
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _082_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_20
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_24
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_28
timestamp 1586364061
transform 1 0 3680 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_36
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_42
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_63
timestamp 1586364061
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_67
timestamp 1586364061
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_90
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_134
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use scs8hd_conb_1  _051_
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_173
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_185
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_197
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_209
timestamp 1586364061
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_14
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_18
timestamp 1586364061
transform 1 0 2760 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_31
timestamp 1586364061
transform 1 0 3956 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_49
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_left_track_27.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_81
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_136
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 406 592
use scs8hd_mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 774 592
use scs8hd_conb_1  _064_
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_162
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_174
timestamp 1586364061
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_38.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24104 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_248
timestamp 1586364061
transform 1 0 23920 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_252
timestamp 1586364061
transform 1 0 24288 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_264
timestamp 1586364061
transform 1 0 25392 0 1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 20128
box -38 -48 1786 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_38
timestamp 1586364061
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 4784 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_49
timestamp 1586364061
transform 1 0 5612 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_53
timestamp 1586364061
transform 1 0 5980 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_57
timestamp 1586364061
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6716 0 -1 20128
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_27.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_90
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_107
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_111
timestamp 1586364061
transform 1 0 11316 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_32_138
timestamp 1586364061
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use scs8hd_conb_1  _063_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_157
timestamp 1586364061
transform 1 0 15548 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_169
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_181
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1932 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_buf_2  _071_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_11
timestamp 1586364061
transform 1 0 2116 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2300 0 -1 21216
box -38 -48 222 592
use scs8hd_buf_2  _072_
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_28
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_32
timestamp 1586364061
transform 1 0 4048 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_45
timestamp 1586364061
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_55
timestamp 1586364061
transform 1 0 6164 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_51
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6348 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6532 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 1786 592
use scs8hd_buf_1  mux_left_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 6992 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_67
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_71
timestamp 1586364061
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_78
timestamp 1586364061
transform 1 0 8280 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_88
timestamp 1586364061
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_107
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_102
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_115
timestamp 1586364061
transform 1 0 11684 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _057_
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_132
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_142
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_146
timestamp 1586364061
transform 1 0 14536 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_161
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_173
timestamp 1586364061
transform 1 0 17020 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_181
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _069_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_55
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_79
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8648 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8464 0 1 21216
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_101
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_116
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12972 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_148
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_160
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_172
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_16
timestamp 1586364061
transform 1 0 2576 0 -1 22304
box -38 -48 222 592
use scs8hd_conb_1  _055_
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 4600 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_20
timestamp 1586364061
transform 1 0 2944 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_25
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_29
timestamp 1586364061
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_35
timestamp 1586364061
transform 1 0 4324 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6440 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_40
timestamp 1586364061
transform 1 0 4784 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_36_52
timestamp 1586364061
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  mux_left_track_27.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 8004 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_69
timestamp 1586364061
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_73
timestamp 1586364061
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_27.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_88
timestamp 1586364061
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_97
timestamp 1586364061
transform 1 0 10028 0 -1 22304
box -38 -48 406 592
use scs8hd_conb_1  _059_
timestamp 1586364061
transform 1 0 9752 0 -1 22304
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_101
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_104
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_114
timestamp 1586364061
transform 1 0 11592 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_118
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_138
timestamp 1586364061
transform 1 0 13800 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_150
timestamp 1586364061
transform 1 0 14904 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 1786 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_30
timestamp 1586364061
transform 1 0 3864 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_36
timestamp 1586364061
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_40
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7728 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 7544 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_67
timestamp 1586364061
transform 1 0 7268 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_91
timestamp 1586364061
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_99
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_111
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _062_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_left_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_131
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 15456 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_154
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 590 592
use scs8hd_buf_1  mux_top_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16284 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_164
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_192
timestamp 1586364061
transform 1 0 18768 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_195
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_26.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_207
timestamp 1586364061
transform 1 0 20148 0 1 22304
box -38 -48 774 592
use scs8hd_decap_12  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_34.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_34.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_249
timestamp 1586364061
transform 1 0 24012 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_261
timestamp 1586364061
transform 1 0 25116 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_273
timestamp 1586364061
transform 1 0 26220 0 1 22304
box -38 -48 406 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 2024 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4600 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 4416 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3036 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_57
timestamp 1586364061
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_61
timestamp 1586364061
transform 1 0 6716 0 -1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 11408 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_110
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_114
timestamp 1586364061
transform 1 0 11592 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_137
timestamp 1586364061
transform 1 0 13708 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _106_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_149
timestamp 1586364061
transform 1 0 14812 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_38_158
timestamp 1586364061
transform 1 0 15640 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_172
timestamp 1586364061
transform 1 0 16928 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_1  mux_top_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17848 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_1  mux_top_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_180
timestamp 1586364061
transform 1 0 17664 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_185
timestamp 1586364061
transform 1 0 18124 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_196
timestamp 1586364061
transform 1 0 19136 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_1  mux_top_track_26.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_208
timestamp 1586364061
transform 1 0 20240 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_8  FILLER_38_218
timestamp 1586364061
transform 1 0 21160 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _093_
timestamp 1586364061
transform 1 0 22172 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_38_226
timestamp 1586364061
transform 1 0 21896 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_233
timestamp 1586364061
transform 1 0 22540 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_2  _090_
timestamp 1586364061
transform 1 0 23828 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_245
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_7
timestamp 1586364061
transform 1 0 1748 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_9
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 2024 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2300 0 1 23392
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_40_21
timestamp 1586364061
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_25
timestamp 1586364061
transform 1 0 3404 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_37
timestamp 1586364061
transform 1 0 4508 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 4324 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4784 0 -1 24480
box -38 -48 1786 592
use scs8hd_mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_55
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_59
timestamp 1586364061
transform 1 0 6532 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_64
timestamp 1586364061
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_79
timestamp 1586364061
transform 1 0 8372 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7544 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_12  FILLER_40_79
timestamp 1586364061
transform 1 0 8372 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_87
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use scs8hd_conb_1  _060_
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_91
timestamp 1586364061
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_91
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9844 0 1 23392
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11408 0 -1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_106
timestamp 1586364061
transform 1 0 10856 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_4  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_conb_1  _058_
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_6  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13800 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 1786 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 15456 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_157
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_161
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_172
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_176
timestamp 1586364061
transform 1 0 17296 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_173
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_169
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 17112 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_160
timestamp 1586364061
transform 1 0 15824 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 19320 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 18216 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_182
timestamp 1586364061
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_190
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_194
timestamp 1586364061
transform 1 0 18952 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_206
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_202
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _097_
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _094_
timestamp 1586364061
transform 1 0 21620 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _095_
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_226
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_230
timestamp 1586364061
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_234
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_240
timestamp 1586364061
transform 1 0 23184 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_buf_2  _092_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _091_
timestamp 1586364061
transform 1 0 23276 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _088_
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_257
timestamp 1586364061
transform 1 0 24748 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_245
timestamp 1586364061
transform 1 0 23644 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_261
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_265
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_40_269
timestamp 1586364061
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_1  mux_left_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2392 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 1840 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 2208 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_6
timestamp 1586364061
transform 1 0 1656 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_10
timestamp 1586364061
transform 1 0 2024 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 3956 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_23
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _073_
timestamp 1586364061
transform 1 0 5520 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 6072 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5336 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_44
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_52
timestamp 1586364061
transform 1 0 5888 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_56
timestamp 1586364061
transform 1 0 6256 0 1 24480
box -38 -48 406 592
use scs8hd_conb_1  _061_
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use scs8hd_mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7268 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_60
timestamp 1586364061
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_65
timestamp 1586364061
transform 1 0 7084 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_69
timestamp 1586364061
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9568 0 1 24480
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9384 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_82
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_88
timestamp 1586364061
transform 1 0 9200 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_111
timestamp 1586364061
transform 1 0 11316 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_115
timestamp 1586364061
transform 1 0 11684 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_144
timestamp 1586364061
transform 1 0 14352 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_156
timestamp 1586364061
transform 1 0 15456 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_168
timestamp 1586364061
transform 1 0 16560 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_41_180
timestamp 1586364061
transform 1 0 17664 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_buf_2  _068_
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use scs8hd_buf_2  _070_
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_7
timestamp 1586364061
transform 1 0 1748 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_19
timestamp 1586364061
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use scs8hd_mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4324 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_conb_1  _065_
timestamp 1586364061
transform 1 0 7912 0 -1 25568
box -38 -48 314 592
use scs8hd_conb_1  _067_
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_66
timestamp 1586364061
transform 1 0 7176 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_77
timestamp 1586364061
transform 1 0 8188 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_81
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_42_153
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 13910 0 13966 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 23202 0 23258 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 8848 480 8968 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 10480 480 10600 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 2456 480 2576 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 17960 480 18080 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21360 480 21480 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21904 480 22024 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 13336 480 13456 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16192 480 16312 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 82 nsew default input
rlabel metal3 s 0 23672 480 23792 6 left_top_grid_pin_42_
port 83 nsew default input
rlabel metal3 s 0 24216 480 24336 6 left_top_grid_pin_43_
port 84 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 85 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 86 nsew default input
rlabel metal3 s 0 25984 480 26104 6 left_top_grid_pin_46_
port 87 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 88 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 89 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 90 nsew default input
rlabel metal2 s 4618 0 4674 480 6 prog_clk
port 91 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 92 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 93 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 94 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_37_
port 95 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_38_
port 96 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 97 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_40_
port 98 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_41_
port 99 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 100 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 101 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 27678 28000
<< end >>
