magic
tech EFS8A
magscale 1 2
timestamp 1602532674
<< locali >>
rect 8251 23137 8378 23171
rect 7699 19941 7744 19975
rect 1547 19465 1685 19499
rect 6837 18139 6871 18377
rect 14841 18071 14875 18241
rect 3341 14875 3375 15113
rect 4905 15011 4939 15113
rect 12995 14569 13001 14603
rect 12995 14501 13029 14569
rect 8309 13719 8343 13821
rect 24627 13345 24662 13379
rect 11437 13175 11471 13345
rect 14565 10591 14599 10761
rect 5267 9129 5273 9163
rect 5267 9061 5301 9129
rect 5359 8279 5393 8347
rect 5359 8245 5365 8279
rect 16991 6817 17026 6851
rect 4019 5729 4146 5763
rect 2559 4777 2605 4811
rect 1443 4641 1478 4675
rect 2455 4641 2490 4675
<< viali >>
rect 10241 24157 10275 24191
rect 6193 23817 6227 23851
rect 10241 23817 10275 23851
rect 13369 23817 13403 23851
rect 15853 23817 15887 23851
rect 21005 23817 21039 23851
rect 25145 23817 25179 23851
rect 1869 23681 1903 23715
rect 1476 23613 1510 23647
rect 5708 23613 5742 23647
rect 10057 23613 10091 23647
rect 11228 23613 11262 23647
rect 11621 23613 11655 23647
rect 12884 23613 12918 23647
rect 15368 23613 15402 23647
rect 20821 23613 20855 23647
rect 21373 23613 21407 23647
rect 24644 23613 24678 23647
rect 24731 23545 24765 23579
rect 1547 23477 1581 23511
rect 5779 23477 5813 23511
rect 10701 23477 10735 23511
rect 11299 23477 11333 23511
rect 12955 23477 12989 23511
rect 15439 23477 15473 23511
rect 23029 23273 23063 23307
rect 10885 23205 10919 23239
rect 12449 23205 12483 23239
rect 4112 23137 4146 23171
rect 8217 23137 8251 23171
rect 9756 23137 9790 23171
rect 22845 23137 22879 23171
rect 10793 23069 10827 23103
rect 11069 23069 11103 23103
rect 12357 23069 12391 23103
rect 12909 23001 12943 23035
rect 4215 22933 4249 22967
rect 8447 22933 8481 22967
rect 9827 22933 9861 22967
rect 10425 22933 10459 22967
rect 4077 22729 4111 22763
rect 8861 22729 8895 22763
rect 9321 22729 9355 22763
rect 9781 22729 9815 22763
rect 12265 22729 12299 22763
rect 13461 22729 13495 22763
rect 10425 22593 10459 22627
rect 11069 22593 11103 22627
rect 12541 22593 12575 22627
rect 12817 22593 12851 22627
rect 6653 22525 6687 22559
rect 7113 22525 7147 22559
rect 8677 22525 8711 22559
rect 10517 22457 10551 22491
rect 12633 22457 12667 22491
rect 7481 22389 7515 22423
rect 8309 22389 8343 22423
rect 10149 22389 10183 22423
rect 11345 22389 11379 22423
rect 11897 22389 11931 22423
rect 22845 22389 22879 22423
rect 11253 22185 11287 22219
rect 12817 22185 12851 22219
rect 7573 22117 7607 22151
rect 10241 22117 10275 22151
rect 12541 22117 12575 22151
rect 1476 22049 1510 22083
rect 4512 22049 4546 22083
rect 10885 22049 10919 22083
rect 12357 22049 12391 22083
rect 17024 22049 17058 22083
rect 6377 21981 6411 22015
rect 7481 21981 7515 22015
rect 1547 21913 1581 21947
rect 8033 21913 8067 21947
rect 8493 21913 8527 21947
rect 17095 21913 17129 21947
rect 4583 21845 4617 21879
rect 5181 21845 5215 21879
rect 1593 21641 1627 21675
rect 4537 21641 4571 21675
rect 7849 21641 7883 21675
rect 8217 21641 8251 21675
rect 10149 21641 10183 21675
rect 17049 21641 17083 21675
rect 5273 21505 5307 21539
rect 5549 21505 5583 21539
rect 6929 21505 6963 21539
rect 7573 21505 7607 21539
rect 8493 21505 8527 21539
rect 8769 21505 8803 21539
rect 10977 21505 11011 21539
rect 5365 21369 5399 21403
rect 7021 21369 7055 21403
rect 8585 21369 8619 21403
rect 9781 21369 9815 21403
rect 10701 21369 10735 21403
rect 10793 21369 10827 21403
rect 4997 21301 5031 21335
rect 6653 21301 6687 21335
rect 10517 21301 10551 21335
rect 11897 21301 11931 21335
rect 6929 21097 6963 21131
rect 8493 21097 8527 21131
rect 5641 21029 5675 21063
rect 7021 21029 7055 21063
rect 10517 21029 10551 21063
rect 6193 20961 6227 20995
rect 7665 20961 7699 20995
rect 11989 20961 12023 20995
rect 24660 20961 24694 20995
rect 4077 20893 4111 20927
rect 5549 20893 5583 20927
rect 8585 20893 8619 20927
rect 10425 20893 10459 20927
rect 11897 20893 11931 20927
rect 10977 20825 11011 20859
rect 5181 20757 5215 20791
rect 12909 20757 12943 20791
rect 24731 20757 24765 20791
rect 1593 20553 1627 20587
rect 4629 20553 4663 20587
rect 6285 20553 6319 20587
rect 7757 20553 7791 20587
rect 10977 20553 11011 20587
rect 24777 20553 24811 20587
rect 25237 20553 25271 20587
rect 5825 20485 5859 20519
rect 10609 20485 10643 20519
rect 11253 20485 11287 20519
rect 11989 20485 12023 20519
rect 4353 20417 4387 20451
rect 5273 20417 5307 20451
rect 12909 20417 12943 20451
rect 13185 20417 13219 20451
rect 1409 20349 1443 20383
rect 1961 20349 1995 20383
rect 4261 20349 4295 20383
rect 6837 20349 6871 20383
rect 8401 20349 8435 20383
rect 8620 20349 8654 20383
rect 9229 20349 9263 20383
rect 9689 20349 9723 20383
rect 24593 20349 24627 20383
rect 5365 20281 5399 20315
rect 7199 20281 7233 20315
rect 9505 20281 9539 20315
rect 10010 20281 10044 20315
rect 12725 20281 12759 20315
rect 13001 20281 13035 20315
rect 3525 20213 3559 20247
rect 5089 20213 5123 20247
rect 6653 20213 6687 20247
rect 8723 20213 8757 20247
rect 24409 20213 24443 20247
rect 1823 20009 1857 20043
rect 6377 20009 6411 20043
rect 7297 20009 7331 20043
rect 8309 20009 8343 20043
rect 10609 20009 10643 20043
rect 12357 20009 12391 20043
rect 5819 19941 5853 19975
rect 7665 19941 7699 19975
rect 10010 19941 10044 19975
rect 11758 19941 11792 19975
rect 13185 19941 13219 19975
rect 1752 19873 1786 19907
rect 2764 19873 2798 19907
rect 4445 19873 4479 19907
rect 13737 19873 13771 19907
rect 5457 19805 5491 19839
rect 7389 19805 7423 19839
rect 9689 19805 9723 19839
rect 11437 19805 11471 19839
rect 2835 19669 2869 19703
rect 4629 19669 4663 19703
rect 5181 19669 5215 19703
rect 6837 19669 6871 19703
rect 12817 19669 12851 19703
rect 1685 19465 1719 19499
rect 3065 19465 3099 19499
rect 7849 19465 7883 19499
rect 9873 19465 9907 19499
rect 11437 19465 11471 19499
rect 13737 19465 13771 19499
rect 8677 19397 8711 19431
rect 10241 19397 10275 19431
rect 5917 19329 5951 19363
rect 9597 19329 9631 19363
rect 13185 19329 13219 19363
rect 1476 19261 1510 19295
rect 2672 19261 2706 19295
rect 4169 19261 4203 19295
rect 5181 19261 5215 19295
rect 5733 19261 5767 19295
rect 6653 19261 6687 19295
rect 7113 19261 7147 19295
rect 7297 19261 7331 19295
rect 8861 19261 8895 19295
rect 9321 19261 9355 19295
rect 10425 19261 10459 19295
rect 10885 19261 10919 19295
rect 12817 19193 12851 19227
rect 12909 19193 12943 19227
rect 1961 19125 1995 19159
rect 2329 19125 2363 19159
rect 2743 19125 2777 19159
rect 3433 19125 3467 19159
rect 4353 19125 4387 19159
rect 4629 19125 4663 19159
rect 4997 19125 5031 19159
rect 6285 19125 6319 19159
rect 6929 19125 6963 19159
rect 8217 19125 8251 19159
rect 10701 19125 10735 19159
rect 11805 19125 11839 19159
rect 1593 18921 1627 18955
rect 5365 18921 5399 18955
rect 5733 18921 5767 18955
rect 9505 18921 9539 18955
rect 12173 18921 12207 18955
rect 12817 18921 12851 18955
rect 24777 18921 24811 18955
rect 4997 18853 5031 18887
rect 6009 18853 6043 18887
rect 7573 18853 7607 18887
rect 10701 18853 10735 18887
rect 11574 18853 11608 18887
rect 1409 18785 1443 18819
rect 2973 18785 3007 18819
rect 4905 18785 4939 18819
rect 9689 18785 9723 18819
rect 10149 18785 10183 18819
rect 13185 18785 13219 18819
rect 15368 18785 15402 18819
rect 24593 18785 24627 18819
rect 5917 18717 5951 18751
rect 6193 18717 6227 18751
rect 7205 18717 7239 18751
rect 7481 18717 7515 18751
rect 7757 18717 7791 18751
rect 10425 18717 10459 18751
rect 11253 18717 11287 18751
rect 13829 18717 13863 18751
rect 11069 18649 11103 18683
rect 15439 18649 15473 18683
rect 3157 18581 3191 18615
rect 6929 18581 6963 18615
rect 8861 18581 8895 18615
rect 1593 18377 1627 18411
rect 2053 18377 2087 18411
rect 2329 18377 2363 18411
rect 3433 18377 3467 18411
rect 4997 18377 5031 18411
rect 6193 18377 6227 18411
rect 6837 18377 6871 18411
rect 8309 18377 8343 18411
rect 9873 18377 9907 18411
rect 11437 18377 11471 18411
rect 11805 18377 11839 18411
rect 13185 18377 13219 18411
rect 25421 18377 25455 18411
rect 4353 18309 4387 18343
rect 5917 18241 5951 18275
rect 1409 18173 1443 18207
rect 2564 18173 2598 18207
rect 2973 18173 3007 18207
rect 4169 18173 4203 18207
rect 5825 18173 5859 18207
rect 7941 18309 7975 18343
rect 24731 18309 24765 18343
rect 7021 18241 7055 18275
rect 7665 18241 7699 18275
rect 9229 18241 9263 18275
rect 14657 18241 14691 18275
rect 14841 18241 14875 18275
rect 25145 18241 25179 18275
rect 12484 18173 12518 18207
rect 2651 18105 2685 18139
rect 6837 18105 6871 18139
rect 7113 18105 7147 18139
rect 8953 18105 8987 18139
rect 9045 18105 9079 18139
rect 10517 18105 10551 18139
rect 10609 18105 10643 18139
rect 11161 18105 11195 18139
rect 12173 18105 12207 18139
rect 14013 18105 14047 18139
rect 14105 18105 14139 18139
rect 15393 18173 15427 18207
rect 15577 18173 15611 18207
rect 24660 18173 24694 18207
rect 15485 18105 15519 18139
rect 4629 18037 4663 18071
rect 6653 18037 6687 18071
rect 8769 18037 8803 18071
rect 10241 18037 10275 18071
rect 12587 18037 12621 18071
rect 13829 18037 13863 18071
rect 14841 18037 14875 18071
rect 15025 18037 15059 18071
rect 4905 17833 4939 17867
rect 6469 17833 6503 17867
rect 7481 17833 7515 17867
rect 11989 17833 12023 17867
rect 5641 17765 5675 17799
rect 6193 17765 6227 17799
rect 7021 17765 7055 17799
rect 10241 17765 10275 17799
rect 13001 17765 13035 17799
rect 13093 17765 13127 17799
rect 15485 17765 15519 17799
rect 2605 17697 2639 17731
rect 4077 17697 4111 17731
rect 8033 17697 8067 17731
rect 8493 17697 8527 17731
rect 10333 17697 10367 17731
rect 11805 17697 11839 17731
rect 5549 17629 5583 17663
rect 8769 17629 8803 17663
rect 15393 17629 15427 17663
rect 15669 17629 15703 17663
rect 13553 17561 13587 17595
rect 1593 17493 1627 17527
rect 2237 17493 2271 17527
rect 4261 17493 4295 17527
rect 5273 17493 5307 17527
rect 9873 17493 9907 17527
rect 12541 17493 12575 17527
rect 14013 17493 14047 17527
rect 14381 17493 14415 17527
rect 6193 17289 6227 17323
rect 6561 17289 6595 17323
rect 7757 17289 7791 17323
rect 10333 17289 10367 17323
rect 10609 17289 10643 17323
rect 11897 17289 11931 17323
rect 13461 17289 13495 17323
rect 14105 17289 14139 17323
rect 15393 17289 15427 17323
rect 13737 17221 13771 17255
rect 9229 17153 9263 17187
rect 11161 17153 11195 17187
rect 14657 17153 14691 17187
rect 1685 17085 1719 17119
rect 3617 17085 3651 17119
rect 4169 17085 4203 17119
rect 5181 17085 5215 17119
rect 5733 17085 5767 17119
rect 5917 17085 5951 17119
rect 6837 17085 6871 17119
rect 9137 17085 9171 17119
rect 9873 17085 9907 17119
rect 12541 17085 12575 17119
rect 3525 17017 3559 17051
rect 4353 17017 4387 17051
rect 7158 17017 7192 17051
rect 10885 17017 10919 17051
rect 10977 17017 11011 17051
rect 12862 17017 12896 17051
rect 14381 17017 14415 17051
rect 14473 17017 14507 17051
rect 1869 16949 1903 16983
rect 2697 16949 2731 16983
rect 4629 16949 4663 16983
rect 5089 16949 5123 16983
rect 8033 16949 8067 16983
rect 8493 16949 8527 16983
rect 12173 16949 12207 16983
rect 15669 16949 15703 16983
rect 3709 16745 3743 16779
rect 5181 16745 5215 16779
rect 6193 16745 6227 16779
rect 6837 16745 6871 16779
rect 7021 16745 7055 16779
rect 10609 16745 10643 16779
rect 12909 16745 12943 16779
rect 15393 16745 15427 16779
rect 5635 16677 5669 16711
rect 7941 16677 7975 16711
rect 8217 16677 8251 16711
rect 8769 16677 8803 16711
rect 10010 16677 10044 16711
rect 10885 16677 10919 16711
rect 12310 16677 12344 16711
rect 13921 16677 13955 16711
rect 1476 16609 1510 16643
rect 2973 16609 3007 16643
rect 4112 16609 4146 16643
rect 5273 16609 5307 16643
rect 13185 16609 13219 16643
rect 15577 16609 15611 16643
rect 15761 16609 15795 16643
rect 3157 16541 3191 16575
rect 8125 16541 8159 16575
rect 9689 16541 9723 16575
rect 11989 16541 12023 16575
rect 1547 16405 1581 16439
rect 1961 16405 1995 16439
rect 4215 16405 4249 16439
rect 7481 16405 7515 16439
rect 2973 16201 3007 16235
rect 3617 16201 3651 16235
rect 5365 16201 5399 16235
rect 9321 16201 9355 16235
rect 11345 16201 11379 16235
rect 12633 16201 12667 16235
rect 11069 16133 11103 16167
rect 7389 16065 7423 16099
rect 9689 16065 9723 16099
rect 13277 16065 13311 16099
rect 15485 16065 15519 16099
rect 1961 15997 1995 16031
rect 4077 15997 4111 16031
rect 4261 15997 4295 16031
rect 4905 15997 4939 16031
rect 8217 15997 8251 16031
rect 8769 15997 8803 16031
rect 9045 15997 9079 16031
rect 10149 15997 10183 16031
rect 14841 15997 14875 16031
rect 14933 15997 14967 16031
rect 15393 15997 15427 16031
rect 24660 15997 24694 16031
rect 25053 15997 25087 16031
rect 5733 15929 5767 15963
rect 8033 15929 8067 15963
rect 10470 15929 10504 15963
rect 11989 15929 12023 15963
rect 13461 15929 13495 15963
rect 13553 15929 13587 15963
rect 14105 15929 14139 15963
rect 1593 15861 1627 15895
rect 2145 15861 2179 15895
rect 6837 15861 6871 15895
rect 7757 15861 7791 15895
rect 14381 15861 14415 15895
rect 15945 15861 15979 15895
rect 24731 15861 24765 15895
rect 1777 15657 1811 15691
rect 4261 15657 4295 15691
rect 5457 15657 5491 15691
rect 8769 15657 8803 15691
rect 10517 15657 10551 15691
rect 2145 15589 2179 15623
rect 4537 15589 4571 15623
rect 4629 15589 4663 15623
rect 9321 15589 9355 15623
rect 10241 15589 10275 15623
rect 11345 15589 11379 15623
rect 13829 15589 13863 15623
rect 15301 15589 15335 15623
rect 6377 15521 6411 15555
rect 7665 15521 7699 15555
rect 8493 15521 8527 15555
rect 8677 15521 8711 15555
rect 9689 15521 9723 15555
rect 15393 15521 15427 15555
rect 24593 15521 24627 15555
rect 2053 15453 2087 15487
rect 5181 15453 5215 15487
rect 6101 15453 6135 15487
rect 11253 15453 11287 15487
rect 11529 15453 11563 15487
rect 13093 15453 13127 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 2605 15385 2639 15419
rect 14933 15385 14967 15419
rect 24777 15385 24811 15419
rect 7481 15317 7515 15351
rect 9873 15317 9907 15351
rect 13369 15317 13403 15351
rect 1961 15113 1995 15147
rect 3341 15113 3375 15147
rect 3433 15113 3467 15147
rect 4629 15113 4663 15147
rect 4905 15113 4939 15147
rect 6561 15113 6595 15147
rect 9137 15113 9171 15147
rect 10333 15113 10367 15147
rect 13737 15113 13771 15147
rect 15393 15113 15427 15147
rect 23811 15113 23845 15147
rect 24685 15113 24719 15147
rect 3065 15045 3099 15079
rect 2145 14977 2179 15011
rect 2605 14977 2639 15011
rect 4261 15045 4295 15079
rect 8217 15045 8251 15079
rect 3709 14977 3743 15011
rect 4905 14977 4939 15011
rect 5273 14977 5307 15011
rect 9689 14977 9723 15011
rect 11805 14977 11839 15011
rect 12817 14977 12851 15011
rect 5917 14909 5951 14943
rect 7665 14909 7699 14943
rect 8217 14909 8251 14943
rect 8401 14909 8435 14943
rect 15577 14909 15611 14943
rect 16221 14909 16255 14943
rect 16589 14909 16623 14943
rect 23740 14909 23774 14943
rect 24133 14909 24167 14943
rect 2237 14841 2271 14875
rect 3341 14841 3375 14875
rect 3801 14841 3835 14875
rect 5365 14841 5399 14875
rect 6285 14841 6319 14875
rect 9413 14841 9447 14875
rect 9505 14841 9539 14875
rect 10885 14841 10919 14875
rect 12541 14841 12575 14875
rect 12633 14841 12667 14875
rect 14105 14841 14139 14875
rect 14197 14841 14231 14875
rect 14749 14841 14783 14875
rect 5089 14773 5123 14807
rect 7205 14773 7239 14807
rect 8769 14773 8803 14807
rect 11437 14773 11471 14807
rect 12265 14773 12299 14807
rect 2053 14569 2087 14603
rect 3157 14569 3191 14603
rect 3709 14569 3743 14603
rect 4997 14569 5031 14603
rect 5273 14569 5307 14603
rect 6377 14569 6411 14603
rect 6745 14569 6779 14603
rect 7297 14569 7331 14603
rect 11161 14569 11195 14603
rect 12541 14569 12575 14603
rect 13001 14569 13035 14603
rect 13553 14569 13587 14603
rect 14013 14569 14047 14603
rect 15025 14569 15059 14603
rect 1685 14501 1719 14535
rect 2599 14501 2633 14535
rect 4439 14501 4473 14535
rect 10603 14501 10637 14535
rect 5892 14433 5926 14467
rect 7481 14433 7515 14467
rect 8033 14433 8067 14467
rect 8217 14433 8251 14467
rect 10241 14433 10275 14467
rect 15301 14433 15335 14467
rect 15393 14433 15427 14467
rect 2237 14365 2271 14399
rect 4077 14365 4111 14399
rect 7113 14365 7147 14399
rect 12633 14365 12667 14399
rect 14749 14365 14783 14399
rect 16865 14365 16899 14399
rect 5733 14229 5767 14263
rect 5963 14229 5997 14263
rect 8677 14229 8711 14263
rect 9321 14229 9355 14263
rect 12081 14229 12115 14263
rect 2697 14025 2731 14059
rect 3893 14025 3927 14059
rect 5457 14025 5491 14059
rect 6285 14025 6319 14059
rect 7757 14025 7791 14059
rect 9229 14025 9263 14059
rect 13829 14025 13863 14059
rect 15669 14025 15703 14059
rect 6561 13957 6595 13991
rect 8861 13957 8895 13991
rect 10333 13957 10367 13991
rect 16037 13957 16071 13991
rect 1685 13889 1719 13923
rect 3525 13889 3559 13923
rect 6837 13889 6871 13923
rect 8732 13889 8766 13923
rect 8953 13889 8987 13923
rect 10701 13889 10735 13923
rect 14749 13889 14783 13923
rect 15025 13889 15059 13923
rect 2329 13821 2363 13855
rect 4261 13821 4295 13855
rect 4445 13821 4479 13855
rect 4721 13821 4755 13855
rect 4997 13821 5031 13855
rect 5549 13821 5583 13855
rect 8309 13821 8343 13855
rect 11069 13821 11103 13855
rect 11253 13821 11287 13855
rect 11529 13821 11563 13855
rect 12909 13821 12943 13855
rect 16313 13821 16347 13855
rect 18245 13821 18279 13855
rect 18797 13821 18831 13855
rect 1777 13753 1811 13787
rect 3157 13753 3191 13787
rect 7158 13753 7192 13787
rect 8125 13753 8159 13787
rect 8585 13753 8619 13787
rect 12173 13753 12207 13787
rect 12725 13753 12759 13787
rect 13230 13753 13264 13787
rect 14565 13753 14599 13787
rect 14841 13753 14875 13787
rect 16221 13753 16255 13787
rect 5733 13685 5767 13719
rect 8309 13685 8343 13719
rect 8401 13685 8435 13719
rect 9873 13685 9907 13719
rect 11897 13685 11931 13719
rect 14197 13685 14231 13719
rect 18429 13685 18463 13719
rect 1685 13481 1719 13515
rect 3249 13481 3283 13515
rect 4169 13481 4203 13515
rect 11989 13481 12023 13515
rect 15393 13481 15427 13515
rect 17003 13481 17037 13515
rect 2053 13413 2087 13447
rect 2605 13413 2639 13447
rect 10695 13413 10729 13447
rect 12265 13413 12299 13447
rect 12817 13413 12851 13447
rect 13093 13413 13127 13447
rect 14381 13413 14415 13447
rect 4169 13345 4203 13379
rect 4537 13345 4571 13379
rect 5641 13345 5675 13379
rect 7113 13345 7147 13379
rect 11253 13345 11287 13379
rect 11437 13345 11471 13379
rect 13645 13345 13679 13379
rect 15301 13345 15335 13379
rect 15761 13345 15795 13379
rect 16932 13345 16966 13379
rect 24593 13345 24627 13379
rect 1961 13277 1995 13311
rect 3617 13277 3651 13311
rect 7481 13277 7515 13311
rect 7573 13277 7607 13311
rect 10333 13277 10367 13311
rect 2973 13209 3007 13243
rect 7278 13209 7312 13243
rect 8677 13209 8711 13243
rect 9965 13209 9999 13243
rect 12173 13277 12207 13311
rect 14013 13277 14047 13311
rect 13810 13209 13844 13243
rect 14657 13209 14691 13243
rect 5825 13141 5859 13175
rect 6285 13141 6319 13175
rect 7021 13141 7055 13175
rect 7389 13141 7423 13175
rect 8217 13141 8251 13175
rect 9045 13141 9079 13175
rect 11437 13141 11471 13175
rect 11529 13141 11563 13175
rect 13461 13141 13495 13175
rect 13921 13141 13955 13175
rect 24731 13141 24765 13175
rect 1869 12937 1903 12971
rect 3341 12937 3375 12971
rect 4077 12937 4111 12971
rect 7205 12937 7239 12971
rect 8677 12937 8711 12971
rect 11345 12937 11379 12971
rect 14178 12937 14212 12971
rect 14473 12937 14507 12971
rect 24685 12937 24719 12971
rect 2329 12869 2363 12903
rect 3709 12869 3743 12903
rect 6285 12869 6319 12903
rect 8309 12869 8343 12903
rect 9762 12869 9796 12903
rect 9873 12869 9907 12903
rect 10977 12869 11011 12903
rect 13093 12869 13127 12903
rect 13737 12869 13771 12903
rect 14289 12869 14323 12903
rect 15301 12869 15335 12903
rect 1547 12801 1581 12835
rect 4445 12801 4479 12835
rect 8180 12801 8214 12835
rect 8401 12801 8435 12835
rect 9965 12801 9999 12835
rect 10701 12801 10735 12835
rect 12541 12801 12575 12835
rect 14381 12801 14415 12835
rect 16589 12801 16623 12835
rect 1460 12733 1494 12767
rect 2421 12733 2455 12767
rect 4813 12733 4847 12767
rect 5181 12733 5215 12767
rect 5457 12733 5491 12767
rect 7021 12733 7055 12767
rect 11161 12733 11195 12767
rect 11621 12733 11655 12767
rect 14013 12733 14047 12767
rect 15577 12733 15611 12767
rect 16037 12733 16071 12767
rect 16957 12733 16991 12767
rect 2742 12665 2776 12699
rect 7481 12665 7515 12699
rect 8033 12665 8067 12699
rect 9597 12665 9631 12699
rect 10333 12665 10367 12699
rect 12265 12665 12299 12699
rect 12633 12665 12667 12699
rect 4997 12597 5031 12631
rect 6653 12597 6687 12631
rect 7941 12597 7975 12631
rect 9137 12597 9171 12631
rect 9505 12597 9539 12631
rect 15669 12597 15703 12631
rect 17325 12597 17359 12631
rect 1685 12393 1719 12427
rect 6285 12393 6319 12427
rect 7849 12393 7883 12427
rect 10885 12393 10919 12427
rect 11897 12393 11931 12427
rect 12633 12393 12667 12427
rect 16313 12393 16347 12427
rect 1961 12325 1995 12359
rect 2421 12325 2455 12359
rect 2513 12325 2547 12359
rect 11253 12325 11287 12359
rect 13185 12325 13219 12359
rect 13553 12325 13587 12359
rect 13829 12325 13863 12359
rect 15117 12325 15151 12359
rect 15485 12325 15519 12359
rect 4077 12257 4111 12291
rect 4537 12257 4571 12291
rect 5641 12257 5675 12291
rect 7205 12257 7239 12291
rect 9689 12257 9723 12291
rect 11621 12257 11655 12291
rect 12081 12257 12115 12291
rect 17877 12257 17911 12291
rect 2697 12189 2731 12223
rect 4629 12189 4663 12223
rect 6009 12189 6043 12223
rect 7573 12189 7607 12223
rect 10057 12189 10091 12223
rect 13737 12189 13771 12223
rect 14013 12189 14047 12223
rect 15393 12189 15427 12223
rect 16865 12189 16899 12223
rect 5806 12121 5840 12155
rect 9965 12121 9999 12155
rect 14657 12121 14691 12155
rect 15945 12121 15979 12155
rect 3433 12053 3467 12087
rect 5181 12053 5215 12087
rect 5917 12053 5951 12087
rect 6653 12053 6687 12087
rect 7021 12053 7055 12087
rect 7343 12053 7377 12087
rect 7481 12053 7515 12087
rect 8217 12053 8251 12087
rect 8677 12053 8711 12087
rect 9045 12053 9079 12087
rect 9413 12053 9447 12087
rect 9827 12053 9861 12087
rect 10149 12053 10183 12087
rect 18061 12053 18095 12087
rect 2789 11849 2823 11883
rect 4169 11849 4203 11883
rect 4537 11849 4571 11883
rect 5825 11849 5859 11883
rect 6975 11849 7009 11883
rect 7389 11849 7423 11883
rect 8585 11849 8619 11883
rect 9137 11849 9171 11883
rect 9597 11849 9631 11883
rect 12173 11849 12207 11883
rect 12909 11849 12943 11883
rect 14749 11849 14783 11883
rect 24731 11849 24765 11883
rect 2513 11781 2547 11815
rect 6193 11781 6227 11815
rect 8401 11781 8435 11815
rect 10609 11781 10643 11815
rect 15485 11781 15519 11815
rect 1501 11713 1535 11747
rect 2973 11713 3007 11747
rect 6561 11713 6595 11747
rect 8493 11713 8527 11747
rect 11805 11713 11839 11747
rect 14933 11713 14967 11747
rect 15945 11713 15979 11747
rect 16405 11713 16439 11747
rect 4721 11645 4755 11679
rect 5273 11645 5307 11679
rect 6872 11645 6906 11679
rect 8272 11645 8306 11679
rect 9689 11645 9723 11679
rect 10793 11645 10827 11679
rect 11253 11645 11287 11679
rect 13093 11645 13127 11679
rect 16313 11645 16347 11679
rect 16497 11645 16531 11679
rect 24660 11645 24694 11679
rect 25145 11645 25179 11679
rect 1593 11577 1627 11611
rect 2145 11577 2179 11611
rect 3335 11577 3369 11611
rect 8125 11577 8159 11611
rect 10149 11577 10183 11611
rect 11529 11577 11563 11611
rect 13414 11577 13448 11611
rect 15002 11577 15036 11611
rect 3893 11509 3927 11543
rect 4813 11509 4847 11543
rect 7941 11509 7975 11543
rect 9873 11509 9907 11543
rect 14013 11509 14047 11543
rect 14381 11509 14415 11543
rect 18245 11509 18279 11543
rect 2329 11305 2363 11339
rect 3433 11305 3467 11339
rect 7297 11305 7331 11339
rect 9965 11305 9999 11339
rect 13737 11305 13771 11339
rect 13921 11305 13955 11339
rect 14933 11305 14967 11339
rect 15393 11305 15427 11339
rect 2513 11237 2547 11271
rect 2605 11237 2639 11271
rect 3157 11237 3191 11271
rect 4398 11237 4432 11271
rect 5641 11237 5675 11271
rect 8585 11237 8619 11271
rect 11345 11237 11379 11271
rect 12535 11237 12569 11271
rect 16865 11237 16899 11271
rect 1476 11169 1510 11203
rect 4077 11169 4111 11203
rect 5825 11169 5859 11203
rect 6377 11169 6411 11203
rect 6929 11169 6963 11203
rect 7849 11169 7883 11203
rect 10701 11169 10735 11203
rect 11069 11169 11103 11203
rect 12173 11169 12207 11203
rect 15301 11169 15335 11203
rect 15761 11169 15795 11203
rect 16957 11169 16991 11203
rect 3893 11101 3927 11135
rect 6285 11101 6319 11135
rect 7996 11101 8030 11135
rect 8217 11101 8251 11135
rect 1547 11033 1581 11067
rect 7665 11033 7699 11067
rect 1961 10965 1995 10999
rect 4997 10965 5031 10999
rect 5273 10965 5307 10999
rect 8125 10965 8159 10999
rect 8861 10965 8895 10999
rect 9505 10965 9539 10999
rect 10241 10965 10275 10999
rect 13093 10965 13127 10999
rect 14473 10965 14507 10999
rect 4169 10761 4203 10795
rect 4537 10761 4571 10795
rect 5917 10761 5951 10795
rect 6653 10761 6687 10795
rect 9965 10761 9999 10795
rect 10241 10761 10275 10795
rect 10701 10761 10735 10795
rect 12265 10761 12299 10795
rect 12817 10761 12851 10795
rect 14565 10761 14599 10795
rect 14657 10761 14691 10795
rect 15853 10761 15887 10795
rect 16543 10761 16577 10795
rect 3617 10693 3651 10727
rect 7573 10693 7607 10727
rect 8355 10693 8389 10727
rect 8493 10693 8527 10727
rect 9689 10693 9723 10727
rect 13185 10693 13219 10727
rect 3065 10625 3099 10659
rect 6193 10625 6227 10659
rect 6837 10625 6871 10659
rect 8582 10625 8616 10659
rect 9321 10625 9355 10659
rect 14289 10625 14323 10659
rect 16865 10693 16899 10727
rect 2053 10557 2087 10591
rect 4629 10557 4663 10591
rect 5181 10557 5215 10591
rect 8217 10557 8251 10591
rect 9781 10557 9815 10591
rect 10977 10557 11011 10591
rect 11253 10557 11287 10591
rect 11805 10557 11839 10591
rect 14013 10557 14047 10591
rect 14565 10557 14599 10591
rect 14841 10557 14875 10591
rect 15301 10557 15335 10591
rect 16221 10557 16255 10591
rect 16440 10557 16474 10591
rect 17233 10557 17267 10591
rect 23740 10557 23774 10591
rect 24133 10557 24167 10591
rect 3157 10489 3191 10523
rect 8953 10489 8987 10523
rect 11529 10489 11563 10523
rect 13369 10489 13403 10523
rect 13461 10489 13495 10523
rect 1685 10421 1719 10455
rect 2421 10421 2455 10455
rect 2881 10421 2915 10455
rect 4721 10421 4755 10455
rect 7849 10421 7883 10455
rect 14933 10421 14967 10455
rect 23811 10421 23845 10455
rect 4721 10217 4755 10251
rect 6377 10217 6411 10251
rect 9321 10217 9355 10251
rect 12265 10217 12299 10251
rect 12909 10217 12943 10251
rect 1777 10149 1811 10183
rect 2973 10149 3007 10183
rect 7021 10149 7055 10183
rect 10425 10149 10459 10183
rect 10885 10149 10919 10183
rect 2697 10081 2731 10115
rect 4905 10081 4939 10115
rect 5181 10081 5215 10115
rect 6193 10081 6227 10115
rect 7573 10081 7607 10115
rect 7720 10081 7754 10115
rect 9689 10081 9723 10115
rect 11345 10081 11379 10115
rect 13093 10081 13127 10115
rect 13277 10081 13311 10115
rect 15945 10081 15979 10115
rect 1685 10013 1719 10047
rect 3709 10013 3743 10047
rect 7481 10013 7515 10047
rect 7941 10013 7975 10047
rect 10057 10013 10091 10047
rect 11253 10013 11287 10047
rect 2237 9945 2271 9979
rect 4353 9945 4387 9979
rect 8953 9945 8987 9979
rect 9965 9945 9999 9979
rect 3433 9877 3467 9911
rect 7849 9877 7883 9911
rect 8033 9877 8067 9911
rect 8585 9877 8619 9911
rect 9854 9877 9888 9911
rect 14841 9877 14875 9911
rect 15577 9877 15611 9911
rect 1685 9673 1719 9707
rect 3801 9673 3835 9707
rect 5917 9673 5951 9707
rect 6561 9673 6595 9707
rect 12173 9673 12207 9707
rect 14381 9673 14415 9707
rect 16129 9673 16163 9707
rect 4261 9605 4295 9639
rect 11621 9605 11655 9639
rect 12909 9605 12943 9639
rect 16497 9605 16531 9639
rect 2145 9537 2179 9571
rect 4813 9537 4847 9571
rect 6285 9537 6319 9571
rect 10701 9537 10735 9571
rect 13093 9537 13127 9571
rect 15209 9537 15243 9571
rect 15669 9537 15703 9571
rect 6837 9469 6871 9503
rect 7389 9469 7423 9503
rect 9137 9469 9171 9503
rect 9505 9469 9539 9503
rect 14013 9469 14047 9503
rect 14933 9469 14967 9503
rect 1961 9401 1995 9435
rect 2466 9401 2500 9435
rect 4629 9401 4663 9435
rect 4905 9401 4939 9435
rect 5457 9401 5491 9435
rect 9781 9401 9815 9435
rect 10793 9401 10827 9435
rect 11345 9401 11379 9435
rect 13414 9401 13448 9435
rect 15301 9401 15335 9435
rect 3065 9333 3099 9367
rect 6929 9333 6963 9367
rect 7849 9333 7883 9367
rect 8309 9333 8343 9367
rect 8953 9333 8987 9367
rect 10149 9333 10183 9367
rect 10517 9333 10551 9367
rect 4721 9129 4755 9163
rect 5273 9129 5307 9163
rect 9045 9129 9079 9163
rect 12449 9129 12483 9163
rect 12817 9129 12851 9163
rect 14013 9129 14047 9163
rect 2053 9061 2087 9095
rect 2605 9061 2639 9095
rect 7205 9061 7239 9095
rect 11345 9061 11379 9095
rect 13414 9061 13448 9095
rect 15485 9061 15519 9095
rect 6653 8993 6687 9027
rect 6837 8993 6871 9027
rect 8033 8993 8067 9027
rect 8585 8993 8619 9027
rect 9689 8993 9723 9027
rect 16957 8993 16991 9027
rect 1961 8925 1995 8959
rect 4905 8925 4939 8959
rect 8769 8925 8803 8959
rect 11253 8925 11287 8959
rect 11897 8925 11931 8959
rect 13093 8925 13127 8959
rect 15117 8925 15151 8959
rect 15393 8925 15427 8959
rect 16037 8925 16071 8959
rect 16865 8925 16899 8959
rect 10149 8857 10183 8891
rect 1685 8789 1719 8823
rect 5825 8789 5859 8823
rect 7665 8789 7699 8823
rect 9873 8789 9907 8823
rect 10517 8789 10551 8823
rect 10885 8789 10919 8823
rect 14289 8789 14323 8823
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 8493 8585 8527 8619
rect 9505 8585 9539 8619
rect 9781 8585 9815 8619
rect 12173 8585 12207 8619
rect 13645 8585 13679 8619
rect 15577 8585 15611 8619
rect 16957 8585 16991 8619
rect 25145 8585 25179 8619
rect 6653 8517 6687 8551
rect 3433 8449 3467 8483
rect 3985 8449 4019 8483
rect 7205 8449 7239 8483
rect 7941 8449 7975 8483
rect 9965 8449 9999 8483
rect 12449 8449 12483 8483
rect 14565 8449 14599 8483
rect 16129 8449 16163 8483
rect 1777 8381 1811 8415
rect 2237 8381 2271 8415
rect 4997 8381 5031 8415
rect 8401 8381 8435 8415
rect 8953 8381 8987 8415
rect 13369 8381 13403 8415
rect 24660 8381 24694 8415
rect 2145 8313 2179 8347
rect 2599 8313 2633 8347
rect 6929 8313 6963 8347
rect 7021 8313 7055 8347
rect 10286 8313 10320 8347
rect 12811 8313 12845 8347
rect 14289 8313 14323 8347
rect 14381 8313 14415 8347
rect 15301 8313 15335 8347
rect 15853 8313 15887 8347
rect 15945 8313 15979 8347
rect 3157 8245 3191 8279
rect 5365 8245 5399 8279
rect 5917 8245 5951 8279
rect 6285 8245 6319 8279
rect 8217 8245 8251 8279
rect 10885 8245 10919 8279
rect 11161 8245 11195 8279
rect 11621 8245 11655 8279
rect 14105 8245 14139 8279
rect 24731 8245 24765 8279
rect 2605 8041 2639 8075
rect 4629 8041 4663 8075
rect 5733 8041 5767 8075
rect 7297 8041 7331 8075
rect 8953 8041 8987 8075
rect 9965 8041 9999 8075
rect 13093 8041 13127 8075
rect 15117 8041 15151 8075
rect 16865 8041 16899 8075
rect 1777 7973 1811 8007
rect 4905 7973 4939 8007
rect 5457 7973 5491 8007
rect 6469 7973 6503 8007
rect 10654 7973 10688 8007
rect 12265 7973 12299 8007
rect 13829 7973 13863 8007
rect 14381 7973 14415 8007
rect 15485 7973 15519 8007
rect 8493 7905 8527 7939
rect 10333 7905 10367 7939
rect 11253 7905 11287 7939
rect 24660 7905 24694 7939
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 4813 7837 4847 7871
rect 6377 7837 6411 7871
rect 6745 7837 6779 7871
rect 7665 7837 7699 7871
rect 7849 7837 7883 7871
rect 9229 7837 9263 7871
rect 12173 7837 12207 7871
rect 12817 7837 12851 7871
rect 13737 7837 13771 7871
rect 15393 7837 15427 7871
rect 15669 7837 15703 7871
rect 2973 7769 3007 7803
rect 3341 7701 3375 7735
rect 24731 7701 24765 7735
rect 2789 7497 2823 7531
rect 3157 7497 3191 7531
rect 6101 7497 6135 7531
rect 6377 7497 6411 7531
rect 9597 7497 9631 7531
rect 10333 7497 10367 7531
rect 10885 7497 10919 7531
rect 11897 7497 11931 7531
rect 15393 7497 15427 7531
rect 16129 7497 16163 7531
rect 7389 7429 7423 7463
rect 24731 7429 24765 7463
rect 1777 7361 1811 7395
rect 2053 7361 2087 7395
rect 9873 7361 9907 7395
rect 12817 7361 12851 7395
rect 13737 7361 13771 7395
rect 14013 7361 14047 7395
rect 3341 7293 3375 7327
rect 4445 7293 4479 7327
rect 4997 7293 5031 7327
rect 5549 7293 5583 7327
rect 7757 7293 7791 7327
rect 7941 7293 7975 7327
rect 9413 7293 9447 7327
rect 10701 7293 10735 7327
rect 14105 7293 14139 7327
rect 15644 7293 15678 7327
rect 16405 7293 16439 7327
rect 24660 7293 24694 7327
rect 25145 7293 25179 7327
rect 1869 7225 1903 7259
rect 3249 7225 3283 7259
rect 8585 7225 8619 7259
rect 12541 7225 12575 7259
rect 12633 7225 12667 7259
rect 4813 7157 4847 7191
rect 5089 7157 5123 7191
rect 6837 7157 6871 7191
rect 12173 7157 12207 7191
rect 15715 7157 15749 7191
rect 25513 7157 25547 7191
rect 2145 6953 2179 6987
rect 4813 6953 4847 6987
rect 8677 6953 8711 6987
rect 9873 6953 9907 6987
rect 10701 6953 10735 6987
rect 10977 6953 11011 6987
rect 12541 6953 12575 6987
rect 12817 6953 12851 6987
rect 14105 6953 14139 6987
rect 2599 6885 2633 6919
rect 4997 6885 5031 6919
rect 8309 6885 8343 6919
rect 12173 6885 12207 6919
rect 2237 6817 2271 6851
rect 5641 6817 5675 6851
rect 6561 6817 6595 6851
rect 7573 6817 7607 6851
rect 9689 6817 9723 6851
rect 12081 6817 12115 6851
rect 13036 6817 13070 6851
rect 15853 6817 15887 6851
rect 16957 6817 16991 6851
rect 7720 6749 7754 6783
rect 7941 6749 7975 6783
rect 13645 6749 13679 6783
rect 6377 6681 6411 6715
rect 17095 6681 17129 6715
rect 1777 6613 1811 6647
rect 3157 6613 3191 6647
rect 6745 6613 6779 6647
rect 7481 6613 7515 6647
rect 7849 6613 7883 6647
rect 13139 6613 13173 6647
rect 16037 6613 16071 6647
rect 5917 6409 5951 6443
rect 7665 6409 7699 6443
rect 7987 6409 8021 6443
rect 8125 6409 8159 6443
rect 8493 6409 8527 6443
rect 11529 6409 11563 6443
rect 13001 6409 13035 6443
rect 15853 6409 15887 6443
rect 9229 6341 9263 6375
rect 21005 6341 21039 6375
rect 2145 6273 2179 6307
rect 3065 6273 3099 6307
rect 4813 6273 4847 6307
rect 7205 6273 7239 6307
rect 8217 6273 8251 6307
rect 12449 6273 12483 6307
rect 3341 6205 3375 6239
rect 4721 6205 4755 6239
rect 4905 6205 4939 6239
rect 20821 6205 20855 6239
rect 21373 6205 21407 6239
rect 1777 6137 1811 6171
rect 1869 6137 1903 6171
rect 3249 6137 3283 6171
rect 7849 6137 7883 6171
rect 8861 6137 8895 6171
rect 2789 6069 2823 6103
rect 6653 6069 6687 6103
rect 9781 6069 9815 6103
rect 17049 6069 17083 6103
rect 3065 5865 3099 5899
rect 4215 5865 4249 5899
rect 8309 5865 8343 5899
rect 8677 5865 8711 5899
rect 1869 5797 1903 5831
rect 2697 5797 2731 5831
rect 7573 5797 7607 5831
rect 3985 5729 4019 5763
rect 7665 5729 7699 5763
rect 1777 5661 1811 5695
rect 2145 5661 2179 5695
rect 8033 5661 8067 5695
rect 7830 5593 7864 5627
rect 7941 5525 7975 5559
rect 2237 5321 2271 5355
rect 3065 5321 3099 5355
rect 8769 5321 8803 5355
rect 4077 5253 4111 5287
rect 8401 5253 8435 5287
rect 1547 5185 1581 5219
rect 1460 5117 1494 5151
rect 1869 5117 1903 5151
rect 2697 5117 2731 5151
rect 2881 5117 2915 5151
rect 7021 5117 7055 5151
rect 8677 5117 8711 5151
rect 6561 5049 6595 5083
rect 7665 5049 7699 5083
rect 8493 5049 8527 5083
rect 7941 4981 7975 5015
rect 9413 4981 9447 5015
rect 1869 4777 1903 4811
rect 2605 4777 2639 4811
rect 7205 4777 7239 4811
rect 8677 4777 8711 4811
rect 1547 4709 1581 4743
rect 1409 4641 1443 4675
rect 2421 4641 2455 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 7665 4573 7699 4607
rect 8309 4437 8343 4471
rect 2421 4233 2455 4267
rect 7665 4233 7699 4267
rect 1547 4165 1581 4199
rect 7297 4165 7331 4199
rect 10609 4097 10643 4131
rect 1444 4029 1478 4063
rect 1869 4029 1903 4063
rect 10517 3961 10551 3995
rect 10930 3961 10964 3995
rect 11529 3893 11563 3927
rect 1593 3689 1627 3723
rect 10701 3689 10735 3723
rect 11529 3621 11563 3655
rect 12081 3621 12115 3655
rect 13461 3553 13495 3587
rect 11437 3485 11471 3519
rect 12909 3485 12943 3519
rect 12541 3349 12575 3383
rect 1547 3145 1581 3179
rect 10379 3145 10413 3179
rect 11437 3145 11471 3179
rect 13461 3145 13495 3179
rect 14473 3145 14507 3179
rect 12541 3009 12575 3043
rect 13185 3009 13219 3043
rect 1444 2941 1478 2975
rect 1869 2941 1903 2975
rect 10308 2941 10342 2975
rect 14080 2941 14114 2975
rect 12633 2873 12667 2907
rect 10793 2805 10827 2839
rect 11713 2805 11747 2839
rect 12265 2805 12299 2839
rect 14151 2805 14185 2839
rect 1547 2601 1581 2635
rect 5871 2601 5905 2635
rect 9919 2601 9953 2635
rect 11667 2601 11701 2635
rect 1476 2465 1510 2499
rect 5800 2465 5834 2499
rect 9816 2465 9850 2499
rect 10241 2465 10275 2499
rect 11596 2465 11630 2499
rect 14105 2465 14139 2499
rect 14657 2465 14691 2499
rect 19048 2465 19082 2499
rect 1869 2397 1903 2431
rect 6285 2261 6319 2295
rect 12081 2261 12115 2295
rect 14289 2261 14323 2295
rect 19119 2261 19153 2295
rect 19533 2261 19567 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10229 24191 10287 24197
rect 10229 24188 10241 24191
rect 10192 24160 10241 24188
rect 10192 24148 10198 24160
rect 10229 24157 10241 24160
rect 10275 24157 10287 24191
rect 10229 24151 10287 24157
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 6181 23851 6239 23857
rect 6181 23817 6193 23851
rect 6227 23848 6239 23851
rect 6914 23848 6920 23860
rect 6227 23820 6920 23848
rect 6227 23817 6239 23820
rect 6181 23811 6239 23817
rect 1302 23672 1308 23724
rect 1360 23712 1366 23724
rect 1857 23715 1915 23721
rect 1857 23712 1869 23715
rect 1360 23684 1869 23712
rect 1360 23672 1366 23684
rect 1479 23653 1507 23684
rect 1857 23681 1869 23684
rect 1903 23681 1915 23715
rect 1857 23675 1915 23681
rect 1464 23647 1522 23653
rect 1464 23613 1476 23647
rect 1510 23613 1522 23647
rect 1464 23607 1522 23613
rect 5696 23647 5754 23653
rect 5696 23613 5708 23647
rect 5742 23644 5754 23647
rect 6196 23644 6224 23811
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 10229 23851 10287 23857
rect 10229 23817 10241 23851
rect 10275 23848 10287 23851
rect 10870 23848 10876 23860
rect 10275 23820 10876 23848
rect 10275 23817 10287 23820
rect 10229 23811 10287 23817
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 13357 23851 13415 23857
rect 13357 23817 13369 23851
rect 13403 23848 13415 23851
rect 14826 23848 14832 23860
rect 13403 23820 14832 23848
rect 13403 23817 13415 23820
rect 13357 23811 13415 23817
rect 5742 23616 6224 23644
rect 10045 23647 10103 23653
rect 5742 23613 5754 23616
rect 5696 23607 5754 23613
rect 10045 23613 10057 23647
rect 10091 23644 10103 23647
rect 10091 23616 10732 23644
rect 10091 23613 10103 23616
rect 10045 23607 10103 23613
rect 1118 23468 1124 23520
rect 1176 23508 1182 23520
rect 1535 23511 1593 23517
rect 1535 23508 1547 23511
rect 1176 23480 1547 23508
rect 1176 23468 1182 23480
rect 1535 23477 1547 23480
rect 1581 23477 1593 23511
rect 1535 23471 1593 23477
rect 5442 23468 5448 23520
rect 5500 23508 5506 23520
rect 10704 23517 10732 23616
rect 11054 23604 11060 23656
rect 11112 23644 11118 23656
rect 11216 23647 11274 23653
rect 11216 23644 11228 23647
rect 11112 23616 11228 23644
rect 11112 23604 11118 23616
rect 11216 23613 11228 23616
rect 11262 23644 11274 23647
rect 11609 23647 11667 23653
rect 11609 23644 11621 23647
rect 11262 23616 11621 23644
rect 11262 23613 11274 23616
rect 11216 23607 11274 23613
rect 11609 23613 11621 23616
rect 11655 23613 11667 23647
rect 11609 23607 11667 23613
rect 12872 23647 12930 23653
rect 12872 23613 12884 23647
rect 12918 23644 12930 23647
rect 13372 23644 13400 23811
rect 14826 23808 14832 23820
rect 14884 23808 14890 23860
rect 15841 23851 15899 23857
rect 15841 23817 15853 23851
rect 15887 23848 15899 23851
rect 16850 23848 16856 23860
rect 15887 23820 16856 23848
rect 15887 23817 15899 23820
rect 15841 23811 15899 23817
rect 12918 23616 13400 23644
rect 15356 23647 15414 23653
rect 12918 23613 12930 23616
rect 12872 23607 12930 23613
rect 15356 23613 15368 23647
rect 15402 23644 15414 23647
rect 15856 23644 15884 23811
rect 16850 23808 16856 23820
rect 16908 23808 16914 23860
rect 20993 23851 21051 23857
rect 20993 23817 21005 23851
rect 21039 23848 21051 23851
rect 22830 23848 22836 23860
rect 21039 23820 22836 23848
rect 21039 23817 21051 23820
rect 20993 23811 21051 23817
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 15402 23616 15884 23644
rect 15402 23613 15414 23616
rect 15356 23607 15414 23613
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 19392 23616 20821 23644
rect 19392 23604 19398 23616
rect 20809 23613 20821 23616
rect 20855 23644 20867 23647
rect 21361 23647 21419 23653
rect 21361 23644 21373 23647
rect 20855 23616 21373 23644
rect 20855 23613 20867 23616
rect 20809 23607 20867 23613
rect 21361 23613 21373 23616
rect 21407 23613 21419 23647
rect 21361 23607 21419 23613
rect 24632 23647 24690 23653
rect 24632 23613 24644 23647
rect 24678 23644 24690 23647
rect 25130 23644 25136 23656
rect 24678 23616 25136 23644
rect 24678 23613 24690 23616
rect 24632 23607 24690 23613
rect 25130 23604 25136 23616
rect 25188 23604 25194 23656
rect 21174 23536 21180 23588
rect 21232 23576 21238 23588
rect 24719 23579 24777 23585
rect 24719 23576 24731 23579
rect 21232 23548 24731 23576
rect 21232 23536 21238 23548
rect 24719 23545 24731 23548
rect 24765 23545 24777 23579
rect 24719 23539 24777 23545
rect 5767 23511 5825 23517
rect 5767 23508 5779 23511
rect 5500 23480 5779 23508
rect 5500 23468 5506 23480
rect 5767 23477 5779 23480
rect 5813 23477 5825 23511
rect 5767 23471 5825 23477
rect 10689 23511 10747 23517
rect 10689 23477 10701 23511
rect 10735 23508 10747 23511
rect 11287 23511 11345 23517
rect 11287 23508 11299 23511
rect 10735 23480 11299 23508
rect 10735 23477 10747 23480
rect 10689 23471 10747 23477
rect 11287 23477 11299 23480
rect 11333 23477 11345 23511
rect 11287 23471 11345 23477
rect 12526 23468 12532 23520
rect 12584 23508 12590 23520
rect 12943 23511 13001 23517
rect 12943 23508 12955 23511
rect 12584 23480 12955 23508
rect 12584 23468 12590 23480
rect 12943 23477 12955 23480
rect 12989 23477 13001 23511
rect 12943 23471 13001 23477
rect 14366 23468 14372 23520
rect 14424 23508 14430 23520
rect 15427 23511 15485 23517
rect 15427 23508 15439 23511
rect 14424 23480 15439 23508
rect 14424 23468 14430 23480
rect 15427 23477 15439 23480
rect 15473 23477 15485 23511
rect 15427 23471 15485 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 23017 23307 23075 23313
rect 23017 23273 23029 23307
rect 23063 23304 23075 23307
rect 24854 23304 24860 23316
rect 23063 23276 24860 23304
rect 23063 23273 23075 23276
rect 23017 23267 23075 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 10870 23236 10876 23248
rect 10831 23208 10876 23236
rect 10870 23196 10876 23208
rect 10928 23196 10934 23248
rect 12434 23236 12440 23248
rect 12395 23208 12440 23236
rect 12434 23196 12440 23208
rect 12492 23196 12498 23248
rect 106 23128 112 23180
rect 164 23168 170 23180
rect 4062 23168 4068 23180
rect 4120 23177 4126 23180
rect 4120 23171 4158 23177
rect 164 23140 4068 23168
rect 164 23128 170 23140
rect 4062 23128 4068 23140
rect 4146 23137 4158 23171
rect 4120 23131 4158 23137
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23168 8263 23171
rect 8294 23168 8300 23180
rect 8251 23140 8300 23168
rect 8251 23137 8263 23140
rect 8205 23131 8263 23137
rect 4120 23128 4126 23131
rect 8294 23128 8300 23140
rect 8352 23128 8358 23180
rect 9744 23171 9802 23177
rect 9744 23137 9756 23171
rect 9790 23168 9802 23171
rect 9858 23168 9864 23180
rect 9790 23140 9864 23168
rect 9790 23137 9802 23140
rect 9744 23131 9802 23137
rect 9858 23128 9864 23140
rect 9916 23128 9922 23180
rect 22830 23168 22836 23180
rect 22791 23140 22836 23168
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 10778 23100 10784 23112
rect 10739 23072 10784 23100
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11054 23100 11060 23112
rect 11015 23072 11060 23100
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23100 12403 23103
rect 13446 23100 13452 23112
rect 12391 23072 13452 23100
rect 12391 23069 12403 23072
rect 12345 23063 12403 23069
rect 13446 23060 13452 23072
rect 13504 23060 13510 23112
rect 10796 23032 10824 23060
rect 12802 23032 12808 23044
rect 10796 23004 12808 23032
rect 12802 22992 12808 23004
rect 12860 23032 12866 23044
rect 12897 23035 12955 23041
rect 12897 23032 12909 23035
rect 12860 23004 12909 23032
rect 12860 22992 12866 23004
rect 12897 23001 12909 23004
rect 12943 23001 12955 23035
rect 12897 22995 12955 23001
rect 3234 22924 3240 22976
rect 3292 22964 3298 22976
rect 4203 22967 4261 22973
rect 4203 22964 4215 22967
rect 3292 22936 4215 22964
rect 3292 22924 3298 22936
rect 4203 22933 4215 22936
rect 4249 22933 4261 22967
rect 4203 22927 4261 22933
rect 8435 22967 8493 22973
rect 8435 22933 8447 22967
rect 8481 22964 8493 22967
rect 9214 22964 9220 22976
rect 8481 22936 9220 22964
rect 8481 22933 8493 22936
rect 8435 22927 8493 22933
rect 9214 22924 9220 22936
rect 9272 22924 9278 22976
rect 9306 22924 9312 22976
rect 9364 22964 9370 22976
rect 9815 22967 9873 22973
rect 9815 22964 9827 22967
rect 9364 22936 9827 22964
rect 9364 22924 9370 22936
rect 9815 22933 9827 22936
rect 9861 22933 9873 22967
rect 9815 22927 9873 22933
rect 10134 22924 10140 22976
rect 10192 22964 10198 22976
rect 10410 22964 10416 22976
rect 10192 22936 10416 22964
rect 10192 22924 10198 22936
rect 10410 22924 10416 22936
rect 10468 22924 10474 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 4062 22760 4068 22772
rect 4023 22732 4068 22760
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 8846 22760 8852 22772
rect 8807 22732 8852 22760
rect 8846 22720 8852 22732
rect 8904 22720 8910 22772
rect 9306 22760 9312 22772
rect 9267 22732 9312 22760
rect 9306 22720 9312 22732
rect 9364 22720 9370 22772
rect 9769 22763 9827 22769
rect 9769 22729 9781 22763
rect 9815 22760 9827 22763
rect 9858 22760 9864 22772
rect 9815 22732 9864 22760
rect 9815 22729 9827 22732
rect 9769 22723 9827 22729
rect 9858 22720 9864 22732
rect 9916 22720 9922 22772
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12434 22760 12440 22772
rect 12299 22732 12440 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 13446 22760 13452 22772
rect 13407 22732 13452 22760
rect 13446 22720 13452 22732
rect 13504 22720 13510 22772
rect 10410 22624 10416 22636
rect 10371 22596 10416 22624
rect 10410 22584 10416 22596
rect 10468 22584 10474 22636
rect 11054 22624 11060 22636
rect 11015 22596 11060 22624
rect 11054 22584 11060 22596
rect 11112 22584 11118 22636
rect 12526 22624 12532 22636
rect 12487 22596 12532 22624
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 12802 22624 12808 22636
rect 12763 22596 12808 22624
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 6641 22559 6699 22565
rect 6641 22525 6653 22559
rect 6687 22556 6699 22559
rect 7101 22559 7159 22565
rect 7101 22556 7113 22559
rect 6687 22528 7113 22556
rect 6687 22525 6699 22528
rect 6641 22519 6699 22525
rect 7101 22525 7113 22528
rect 7147 22556 7159 22559
rect 7742 22556 7748 22568
rect 7147 22528 7748 22556
rect 7147 22525 7159 22528
rect 7101 22519 7159 22525
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 8665 22559 8723 22565
rect 8665 22525 8677 22559
rect 8711 22556 8723 22559
rect 9306 22556 9312 22568
rect 8711 22528 9312 22556
rect 8711 22525 8723 22528
rect 8665 22519 8723 22525
rect 9306 22516 9312 22528
rect 9364 22516 9370 22568
rect 10505 22491 10563 22497
rect 10505 22457 10517 22491
rect 10551 22457 10563 22491
rect 10505 22451 10563 22457
rect 12621 22491 12679 22497
rect 12621 22457 12633 22491
rect 12667 22457 12679 22491
rect 12621 22451 12679 22457
rect 7466 22420 7472 22432
rect 7427 22392 7472 22420
rect 7466 22380 7472 22392
rect 7524 22380 7530 22432
rect 8294 22420 8300 22432
rect 8255 22392 8300 22420
rect 8294 22380 8300 22392
rect 8352 22380 8358 22432
rect 10134 22420 10140 22432
rect 10095 22392 10140 22420
rect 10134 22380 10140 22392
rect 10192 22420 10198 22432
rect 10520 22420 10548 22451
rect 10192 22392 10548 22420
rect 10192 22380 10198 22392
rect 10870 22380 10876 22432
rect 10928 22420 10934 22432
rect 11333 22423 11391 22429
rect 11333 22420 11345 22423
rect 10928 22392 11345 22420
rect 10928 22380 10934 22392
rect 11333 22389 11345 22392
rect 11379 22389 11391 22423
rect 11333 22383 11391 22389
rect 11885 22423 11943 22429
rect 11885 22389 11897 22423
rect 11931 22420 11943 22423
rect 12342 22420 12348 22432
rect 11931 22392 12348 22420
rect 11931 22389 11943 22392
rect 11885 22383 11943 22389
rect 12342 22380 12348 22392
rect 12400 22420 12406 22432
rect 12636 22420 12664 22451
rect 22830 22420 22836 22432
rect 12400 22392 12664 22420
rect 22791 22392 22836 22420
rect 12400 22380 12406 22392
rect 22830 22380 22836 22392
rect 22888 22380 22894 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 10778 22176 10784 22228
rect 10836 22216 10842 22228
rect 11241 22219 11299 22225
rect 11241 22216 11253 22219
rect 10836 22188 11253 22216
rect 10836 22176 10842 22188
rect 11241 22185 11253 22188
rect 11287 22185 11299 22219
rect 11241 22179 11299 22185
rect 12618 22176 12624 22228
rect 12676 22216 12682 22228
rect 12805 22219 12863 22225
rect 12805 22216 12817 22219
rect 12676 22188 12817 22216
rect 12676 22176 12682 22188
rect 12805 22185 12817 22188
rect 12851 22185 12863 22219
rect 12805 22179 12863 22185
rect 1210 22108 1216 22160
rect 1268 22148 1274 22160
rect 1268 22120 1507 22148
rect 1268 22108 1274 22120
rect 1479 22089 1507 22120
rect 7466 22108 7472 22160
rect 7524 22148 7530 22160
rect 7561 22151 7619 22157
rect 7561 22148 7573 22151
rect 7524 22120 7573 22148
rect 7524 22108 7530 22120
rect 7561 22117 7573 22120
rect 7607 22117 7619 22151
rect 7561 22111 7619 22117
rect 10134 22108 10140 22160
rect 10192 22148 10198 22160
rect 10229 22151 10287 22157
rect 10229 22148 10241 22151
rect 10192 22120 10241 22148
rect 10192 22108 10198 22120
rect 10229 22117 10241 22120
rect 10275 22117 10287 22151
rect 10229 22111 10287 22117
rect 12434 22108 12440 22160
rect 12492 22148 12498 22160
rect 12529 22151 12587 22157
rect 12529 22148 12541 22151
rect 12492 22120 12541 22148
rect 12492 22108 12498 22120
rect 12529 22117 12541 22120
rect 12575 22117 12587 22151
rect 12529 22111 12587 22117
rect 4522 22089 4528 22092
rect 1464 22083 1522 22089
rect 1464 22049 1476 22083
rect 1510 22049 1522 22083
rect 4500 22083 4528 22089
rect 4500 22080 4512 22083
rect 4435 22052 4512 22080
rect 1464 22043 1522 22049
rect 4500 22049 4512 22052
rect 4580 22080 4586 22092
rect 4890 22080 4896 22092
rect 4580 22052 4896 22080
rect 4500 22043 4528 22049
rect 4522 22040 4528 22043
rect 4580 22040 4586 22052
rect 4890 22040 4896 22052
rect 4948 22040 4954 22092
rect 10870 22080 10876 22092
rect 10831 22052 10876 22080
rect 10870 22040 10876 22052
rect 10928 22040 10934 22092
rect 12342 22080 12348 22092
rect 12303 22052 12348 22080
rect 12342 22040 12348 22052
rect 12400 22040 12406 22092
rect 17034 22089 17040 22092
rect 17012 22083 17040 22089
rect 17012 22080 17024 22083
rect 16947 22052 17024 22080
rect 17012 22049 17024 22052
rect 17092 22080 17098 22092
rect 18874 22080 18880 22092
rect 17092 22052 18880 22080
rect 17012 22043 17040 22049
rect 17034 22040 17040 22043
rect 17092 22040 17098 22052
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 22012 6423 22015
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 6411 21984 7481 22012
rect 6411 21981 6423 21984
rect 6365 21975 6423 21981
rect 7469 21981 7481 21984
rect 7515 22012 7527 22015
rect 8202 22012 8208 22024
rect 7515 21984 8208 22012
rect 7515 21981 7527 21984
rect 7469 21975 7527 21981
rect 8202 21972 8208 21984
rect 8260 21972 8266 22024
rect 1535 21947 1593 21953
rect 1535 21913 1547 21947
rect 1581 21944 1593 21947
rect 6914 21944 6920 21956
rect 1581 21916 6920 21944
rect 1581 21913 1593 21916
rect 1535 21907 1593 21913
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 7558 21904 7564 21956
rect 7616 21944 7622 21956
rect 8021 21947 8079 21953
rect 8021 21944 8033 21947
rect 7616 21916 8033 21944
rect 7616 21904 7622 21916
rect 8021 21913 8033 21916
rect 8067 21944 8079 21947
rect 8294 21944 8300 21956
rect 8067 21916 8300 21944
rect 8067 21913 8079 21916
rect 8021 21907 8079 21913
rect 8294 21904 8300 21916
rect 8352 21904 8358 21956
rect 8478 21944 8484 21956
rect 8391 21916 8484 21944
rect 8478 21904 8484 21916
rect 8536 21944 8542 21956
rect 17083 21947 17141 21953
rect 17083 21944 17095 21947
rect 8536 21916 17095 21944
rect 8536 21904 8542 21916
rect 17083 21913 17095 21916
rect 17129 21913 17141 21947
rect 17083 21907 17141 21913
rect 4571 21879 4629 21885
rect 4571 21845 4583 21879
rect 4617 21876 4629 21879
rect 5169 21879 5227 21885
rect 5169 21876 5181 21879
rect 4617 21848 5181 21876
rect 4617 21845 4629 21848
rect 4571 21839 4629 21845
rect 5169 21845 5181 21848
rect 5215 21876 5227 21879
rect 5258 21876 5264 21888
rect 5215 21848 5264 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1210 21632 1216 21684
rect 1268 21672 1274 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 1268 21644 1593 21672
rect 1268 21632 1274 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 4522 21672 4528 21684
rect 4483 21644 4528 21672
rect 1581 21635 1639 21641
rect 4522 21632 4528 21644
rect 4580 21632 4586 21684
rect 7466 21632 7472 21684
rect 7524 21672 7530 21684
rect 7837 21675 7895 21681
rect 7837 21672 7849 21675
rect 7524 21644 7849 21672
rect 7524 21632 7530 21644
rect 7837 21641 7849 21644
rect 7883 21641 7895 21675
rect 8202 21672 8208 21684
rect 8163 21644 8208 21672
rect 7837 21635 7895 21641
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 10137 21675 10195 21681
rect 10137 21641 10149 21675
rect 10183 21672 10195 21675
rect 10870 21672 10876 21684
rect 10183 21644 10876 21672
rect 10183 21641 10195 21644
rect 10137 21635 10195 21641
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 17034 21672 17040 21684
rect 16995 21644 17040 21672
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 7754 21576 8800 21604
rect 5258 21536 5264 21548
rect 5219 21508 5264 21536
rect 5258 21496 5264 21508
rect 5316 21496 5322 21548
rect 5534 21536 5540 21548
rect 5495 21508 5540 21536
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 6914 21536 6920 21548
rect 6875 21508 6920 21536
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7561 21539 7619 21545
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 7754 21536 7782 21576
rect 8478 21536 8484 21548
rect 7607 21508 7782 21536
rect 8439 21508 8484 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 8478 21496 8484 21508
rect 8536 21496 8542 21548
rect 8772 21545 8800 21576
rect 8757 21539 8815 21545
rect 8757 21505 8769 21539
rect 8803 21536 8815 21539
rect 9122 21536 9128 21548
rect 8803 21508 9128 21536
rect 8803 21505 8815 21508
rect 8757 21499 8815 21505
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10962 21536 10968 21548
rect 9916 21508 10968 21536
rect 9916 21496 9922 21508
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 5353 21403 5411 21409
rect 5353 21369 5365 21403
rect 5399 21369 5411 21403
rect 5353 21363 5411 21369
rect 4982 21332 4988 21344
rect 4943 21304 4988 21332
rect 4982 21292 4988 21304
rect 5040 21332 5046 21344
rect 5368 21332 5396 21363
rect 7006 21360 7012 21412
rect 7064 21400 7070 21412
rect 8570 21400 8576 21412
rect 7064 21372 7109 21400
rect 8531 21372 8576 21400
rect 7064 21360 7070 21372
rect 8570 21360 8576 21372
rect 8628 21360 8634 21412
rect 9769 21403 9827 21409
rect 9769 21369 9781 21403
rect 9815 21400 9827 21403
rect 10686 21400 10692 21412
rect 9815 21372 10692 21400
rect 9815 21369 9827 21372
rect 9769 21363 9827 21369
rect 10686 21360 10692 21372
rect 10744 21360 10750 21412
rect 10781 21403 10839 21409
rect 10781 21369 10793 21403
rect 10827 21400 10839 21403
rect 11974 21400 11980 21412
rect 10827 21372 11980 21400
rect 10827 21369 10839 21372
rect 10781 21363 10839 21369
rect 5040 21304 5396 21332
rect 6641 21335 6699 21341
rect 5040 21292 5046 21304
rect 6641 21301 6653 21335
rect 6687 21332 6699 21335
rect 7024 21332 7052 21360
rect 6687 21304 7052 21332
rect 10505 21335 10563 21341
rect 6687 21301 6699 21304
rect 6641 21295 6699 21301
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 10796 21332 10824 21363
rect 11974 21360 11980 21372
rect 12032 21360 12038 21412
rect 10551 21304 10824 21332
rect 11885 21335 11943 21341
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 11885 21301 11897 21335
rect 11931 21332 11943 21335
rect 12342 21332 12348 21344
rect 11931 21304 12348 21332
rect 11931 21301 11943 21304
rect 11885 21295 11943 21301
rect 12342 21292 12348 21304
rect 12400 21292 12406 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 6914 21128 6920 21140
rect 6875 21100 6920 21128
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 8481 21131 8539 21137
rect 8481 21097 8493 21131
rect 8527 21128 8539 21131
rect 8570 21128 8576 21140
rect 8527 21100 8576 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 5629 21063 5687 21069
rect 5629 21029 5641 21063
rect 5675 21060 5687 21063
rect 6270 21060 6276 21072
rect 5675 21032 6276 21060
rect 5675 21029 5687 21032
rect 5629 21023 5687 21029
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 7006 21060 7012 21072
rect 6967 21032 7012 21060
rect 7006 21020 7012 21032
rect 7064 21020 7070 21072
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20992 6239 20995
rect 7558 20992 7564 21004
rect 6227 20964 7564 20992
rect 6227 20961 6239 20964
rect 6181 20955 6239 20961
rect 7558 20952 7564 20964
rect 7616 20952 7622 21004
rect 7653 20995 7711 21001
rect 7653 20961 7665 20995
rect 7699 20992 7711 20995
rect 8294 20992 8300 21004
rect 7699 20964 8300 20992
rect 7699 20961 7711 20964
rect 7653 20955 7711 20961
rect 8294 20952 8300 20964
rect 8352 20992 8358 21004
rect 8496 20992 8524 21091
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 10505 21063 10563 21069
rect 10505 21029 10517 21063
rect 10551 21060 10563 21063
rect 10551 21032 11376 21060
rect 10551 21029 10563 21032
rect 10505 21023 10563 21029
rect 8352 20964 8524 20992
rect 8352 20952 8358 20964
rect 11348 20936 11376 21032
rect 11974 20992 11980 21004
rect 11935 20964 11980 20992
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 24648 20995 24706 21001
rect 24648 20961 24660 20995
rect 24694 20992 24706 20995
rect 25222 20992 25228 21004
rect 24694 20964 25228 20992
rect 24694 20961 24706 20964
rect 24648 20955 24706 20961
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4065 20927 4123 20933
rect 4065 20924 4077 20927
rect 4028 20896 4077 20924
rect 4028 20884 4034 20896
rect 4065 20893 4077 20896
rect 4111 20893 4123 20927
rect 5534 20924 5540 20936
rect 5495 20896 5540 20924
rect 4065 20887 4123 20893
rect 5534 20884 5540 20896
rect 5592 20884 5598 20936
rect 8573 20927 8631 20933
rect 8573 20893 8585 20927
rect 8619 20924 8631 20927
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 8619 20896 10425 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 10413 20893 10425 20896
rect 10459 20924 10471 20927
rect 11238 20924 11244 20936
rect 10459 20896 11244 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 11885 20927 11943 20933
rect 11885 20924 11897 20927
rect 11388 20896 11897 20924
rect 11388 20884 11394 20896
rect 11885 20893 11897 20896
rect 11931 20893 11943 20927
rect 11885 20887 11943 20893
rect 10962 20856 10968 20868
rect 10923 20828 10968 20856
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 5166 20788 5172 20800
rect 5127 20760 5172 20788
rect 5166 20748 5172 20760
rect 5224 20748 5230 20800
rect 12894 20788 12900 20800
rect 12855 20760 12900 20788
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 18598 20748 18604 20800
rect 18656 20788 18662 20800
rect 24719 20791 24777 20797
rect 24719 20788 24731 20791
rect 18656 20760 24731 20788
rect 18656 20748 18662 20760
rect 24719 20757 24731 20760
rect 24765 20757 24777 20791
rect 24719 20751 24777 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 4617 20587 4675 20593
rect 4617 20553 4629 20587
rect 4663 20584 4675 20587
rect 5534 20584 5540 20596
rect 4663 20556 5540 20584
rect 4663 20553 4675 20556
rect 4617 20547 4675 20553
rect 5534 20544 5540 20556
rect 5592 20584 5598 20596
rect 6270 20584 6276 20596
rect 5592 20556 5856 20584
rect 6183 20556 6276 20584
rect 5592 20544 5598 20556
rect 4706 20476 4712 20528
rect 4764 20516 4770 20528
rect 5166 20516 5172 20528
rect 4764 20488 5172 20516
rect 4764 20476 4770 20488
rect 5166 20476 5172 20488
rect 5224 20516 5230 20528
rect 5828 20525 5856 20556
rect 6270 20544 6276 20556
rect 6328 20584 6334 20596
rect 7742 20584 7748 20596
rect 6328 20556 7748 20584
rect 6328 20544 6334 20556
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 10965 20587 11023 20593
rect 10965 20553 10977 20587
rect 11011 20584 11023 20587
rect 11330 20584 11336 20596
rect 11011 20556 11336 20584
rect 11011 20553 11023 20556
rect 10965 20547 11023 20553
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 24762 20584 24768 20596
rect 24723 20556 24768 20584
rect 24762 20544 24768 20556
rect 24820 20544 24826 20596
rect 25222 20584 25228 20596
rect 25135 20556 25228 20584
rect 25222 20544 25228 20556
rect 25280 20584 25286 20596
rect 26878 20584 26884 20596
rect 25280 20556 26884 20584
rect 25280 20544 25286 20556
rect 26878 20544 26884 20556
rect 26936 20544 26942 20596
rect 5813 20519 5871 20525
rect 5224 20488 5304 20516
rect 5224 20476 5230 20488
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 4982 20448 4988 20460
rect 4387 20420 4988 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 4982 20408 4988 20420
rect 5040 20408 5046 20460
rect 5276 20457 5304 20488
rect 5813 20485 5825 20519
rect 5859 20485 5871 20519
rect 5813 20479 5871 20485
rect 10597 20519 10655 20525
rect 10597 20485 10609 20519
rect 10643 20516 10655 20519
rect 10870 20516 10876 20528
rect 10643 20488 10876 20516
rect 10643 20485 10655 20488
rect 10597 20479 10655 20485
rect 10870 20476 10876 20488
rect 10928 20476 10934 20528
rect 11238 20516 11244 20528
rect 11199 20488 11244 20516
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 11974 20516 11980 20528
rect 11935 20488 11980 20516
rect 11974 20476 11980 20488
rect 12032 20476 12038 20528
rect 12636 20488 13216 20516
rect 5261 20451 5319 20457
rect 5261 20417 5273 20451
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 10778 20408 10784 20460
rect 10836 20448 10842 20460
rect 12636 20448 12664 20488
rect 13188 20460 13216 20488
rect 12894 20448 12900 20460
rect 10836 20420 12664 20448
rect 12855 20420 12900 20448
rect 10836 20408 10842 20420
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13170 20448 13176 20460
rect 13083 20420 13176 20448
rect 13170 20408 13176 20420
rect 13228 20408 13234 20460
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1670 20380 1676 20392
rect 1443 20352 1676 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1670 20340 1676 20352
rect 1728 20380 1734 20392
rect 1949 20383 2007 20389
rect 1949 20380 1961 20383
rect 1728 20352 1961 20380
rect 1728 20340 1734 20352
rect 1949 20349 1961 20352
rect 1995 20349 2007 20383
rect 1949 20343 2007 20349
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20349 4307 20383
rect 4249 20343 4307 20349
rect 3513 20247 3571 20253
rect 3513 20213 3525 20247
rect 3559 20244 3571 20247
rect 4264 20244 4292 20343
rect 6730 20340 6736 20392
rect 6788 20380 6794 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6788 20352 6837 20380
rect 6788 20340 6794 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7742 20340 7748 20392
rect 7800 20380 7806 20392
rect 8389 20383 8447 20389
rect 8389 20380 8401 20383
rect 7800 20352 8401 20380
rect 7800 20340 7806 20352
rect 8389 20349 8401 20352
rect 8435 20380 8447 20383
rect 8608 20383 8666 20389
rect 8608 20380 8620 20383
rect 8435 20352 8620 20380
rect 8435 20349 8447 20352
rect 8389 20343 8447 20349
rect 8608 20349 8620 20352
rect 8654 20349 8666 20383
rect 8608 20343 8666 20349
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 9677 20383 9735 20389
rect 9677 20380 9689 20383
rect 9263 20352 9689 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 9677 20349 9689 20352
rect 9723 20380 9735 20383
rect 10686 20380 10692 20392
rect 9723 20352 10692 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 24581 20383 24639 20389
rect 24581 20380 24593 20383
rect 24412 20352 24593 20380
rect 5350 20312 5356 20324
rect 5311 20284 5356 20312
rect 5350 20272 5356 20284
rect 5408 20272 5414 20324
rect 7187 20315 7245 20321
rect 7187 20312 7199 20315
rect 6656 20284 7199 20312
rect 5077 20247 5135 20253
rect 5077 20244 5089 20247
rect 3559 20216 5089 20244
rect 3559 20213 3571 20216
rect 3513 20207 3571 20213
rect 5077 20213 5089 20216
rect 5123 20244 5135 20247
rect 5368 20244 5396 20272
rect 5123 20216 5396 20244
rect 5123 20213 5135 20216
rect 5077 20207 5135 20213
rect 6270 20204 6276 20256
rect 6328 20244 6334 20256
rect 6656 20253 6684 20284
rect 7187 20281 7199 20284
rect 7233 20312 7245 20315
rect 9493 20315 9551 20321
rect 9493 20312 9505 20315
rect 7233 20284 9505 20312
rect 7233 20281 7245 20284
rect 7187 20275 7245 20281
rect 9493 20281 9505 20284
rect 9539 20312 9551 20315
rect 9858 20312 9864 20324
rect 9539 20284 9864 20312
rect 9539 20281 9551 20284
rect 9493 20275 9551 20281
rect 9858 20272 9864 20284
rect 9916 20312 9922 20324
rect 9998 20315 10056 20321
rect 9998 20312 10010 20315
rect 9916 20284 10010 20312
rect 9916 20272 9922 20284
rect 9998 20281 10010 20284
rect 10044 20281 10056 20315
rect 9998 20275 10056 20281
rect 12713 20315 12771 20321
rect 12713 20281 12725 20315
rect 12759 20312 12771 20315
rect 12986 20312 12992 20324
rect 12759 20284 12992 20312
rect 12759 20281 12771 20284
rect 12713 20275 12771 20281
rect 12986 20272 12992 20284
rect 13044 20272 13050 20324
rect 6641 20247 6699 20253
rect 6641 20244 6653 20247
rect 6328 20216 6653 20244
rect 6328 20204 6334 20216
rect 6641 20213 6653 20216
rect 6687 20213 6699 20247
rect 6641 20207 6699 20213
rect 8711 20247 8769 20253
rect 8711 20213 8723 20247
rect 8757 20244 8769 20247
rect 9398 20244 9404 20256
rect 8757 20216 9404 20244
rect 8757 20213 8769 20216
rect 8711 20207 8769 20213
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 24412 20253 24440 20352
rect 24581 20349 24593 20352
rect 24627 20349 24639 20383
rect 24581 20343 24639 20349
rect 24397 20247 24455 20253
rect 24397 20244 24409 20247
rect 18656 20216 24409 20244
rect 18656 20204 18662 20216
rect 24397 20213 24409 20216
rect 24443 20213 24455 20247
rect 24397 20207 24455 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1811 20043 1869 20049
rect 1811 20009 1823 20043
rect 1857 20040 1869 20043
rect 1946 20040 1952 20052
rect 1857 20012 1952 20040
rect 1857 20009 1869 20012
rect 1811 20003 1869 20009
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 5350 20000 5356 20052
rect 5408 20040 5414 20052
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 5408 20012 6377 20040
rect 5408 20000 5414 20012
rect 6365 20009 6377 20012
rect 6411 20009 6423 20043
rect 6365 20003 6423 20009
rect 7285 20043 7343 20049
rect 7285 20009 7297 20043
rect 7331 20040 7343 20043
rect 8294 20040 8300 20052
rect 7331 20012 8300 20040
rect 7331 20009 7343 20012
rect 7285 20003 7343 20009
rect 8294 20000 8300 20012
rect 8352 20000 8358 20052
rect 10597 20043 10655 20049
rect 10597 20009 10609 20043
rect 10643 20040 10655 20043
rect 11974 20040 11980 20052
rect 10643 20012 11980 20040
rect 10643 20009 10655 20012
rect 10597 20003 10655 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12342 20040 12348 20052
rect 12303 20012 12348 20040
rect 12342 20000 12348 20012
rect 12400 20000 12406 20052
rect 5807 19975 5865 19981
rect 5807 19941 5819 19975
rect 5853 19972 5865 19975
rect 6270 19972 6276 19984
rect 5853 19944 6276 19972
rect 5853 19941 5865 19944
rect 5807 19935 5865 19941
rect 6270 19932 6276 19944
rect 6328 19932 6334 19984
rect 7650 19972 7656 19984
rect 7611 19944 7656 19972
rect 7650 19932 7656 19944
rect 7708 19932 7714 19984
rect 9858 19932 9864 19984
rect 9916 19972 9922 19984
rect 9998 19975 10056 19981
rect 9998 19972 10010 19975
rect 9916 19944 10010 19972
rect 9916 19932 9922 19944
rect 9998 19941 10010 19944
rect 10044 19941 10056 19975
rect 9998 19935 10056 19941
rect 11422 19932 11428 19984
rect 11480 19972 11486 19984
rect 11746 19975 11804 19981
rect 11746 19972 11758 19975
rect 11480 19944 11758 19972
rect 11480 19932 11486 19944
rect 11746 19941 11758 19944
rect 11792 19941 11804 19975
rect 11746 19935 11804 19941
rect 12986 19932 12992 19984
rect 13044 19972 13050 19984
rect 13173 19975 13231 19981
rect 13173 19972 13185 19975
rect 13044 19944 13185 19972
rect 13044 19932 13050 19944
rect 13173 19941 13185 19944
rect 13219 19941 13231 19975
rect 13173 19935 13231 19941
rect 1740 19907 1798 19913
rect 1740 19873 1752 19907
rect 1786 19904 1798 19907
rect 1946 19904 1952 19916
rect 1786 19876 1952 19904
rect 1786 19873 1798 19876
rect 1740 19867 1798 19873
rect 1946 19864 1952 19876
rect 2004 19864 2010 19916
rect 2752 19907 2810 19913
rect 2752 19873 2764 19907
rect 2798 19904 2810 19907
rect 3418 19904 3424 19916
rect 2798 19876 3424 19904
rect 2798 19873 2810 19876
rect 2752 19867 2810 19873
rect 3418 19864 3424 19876
rect 3476 19864 3482 19916
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 4614 19904 4620 19916
rect 4479 19876 4620 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4614 19864 4620 19876
rect 4672 19864 4678 19916
rect 13722 19904 13728 19916
rect 13683 19876 13728 19904
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 5442 19836 5448 19848
rect 5403 19808 5448 19836
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19836 7435 19839
rect 8202 19836 8208 19848
rect 7423 19808 8208 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9674 19836 9680 19848
rect 9635 19808 9680 19836
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 11425 19839 11483 19845
rect 11425 19805 11437 19839
rect 11471 19836 11483 19839
rect 11698 19836 11704 19848
rect 11471 19808 11704 19836
rect 11471 19805 11483 19808
rect 11425 19799 11483 19805
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 2038 19660 2044 19712
rect 2096 19700 2102 19712
rect 2823 19703 2881 19709
rect 2823 19700 2835 19703
rect 2096 19672 2835 19700
rect 2096 19660 2102 19672
rect 2823 19669 2835 19672
rect 2869 19669 2881 19703
rect 2823 19663 2881 19669
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 4617 19703 4675 19709
rect 4617 19700 4629 19703
rect 3936 19672 4629 19700
rect 3936 19660 3942 19672
rect 4617 19669 4629 19672
rect 4663 19669 4675 19703
rect 5166 19700 5172 19712
rect 5127 19672 5172 19700
rect 4617 19663 4675 19669
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 6825 19703 6883 19709
rect 6825 19700 6837 19703
rect 6788 19672 6837 19700
rect 6788 19660 6794 19672
rect 6825 19669 6837 19672
rect 6871 19669 6883 19703
rect 12802 19700 12808 19712
rect 12763 19672 12808 19700
rect 6825 19663 6883 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1670 19496 1676 19508
rect 1631 19468 1676 19496
rect 1670 19456 1676 19468
rect 1728 19456 1734 19508
rect 2866 19456 2872 19508
rect 2924 19496 2930 19508
rect 3053 19499 3111 19505
rect 3053 19496 3065 19499
rect 2924 19468 3065 19496
rect 2924 19456 2930 19468
rect 3053 19465 3065 19468
rect 3099 19465 3111 19499
rect 3053 19459 3111 19465
rect 6270 19456 6276 19508
rect 6328 19496 6334 19508
rect 7650 19496 7656 19508
rect 6328 19468 7656 19496
rect 6328 19456 6334 19468
rect 7650 19456 7656 19468
rect 7708 19496 7714 19508
rect 7837 19499 7895 19505
rect 7837 19496 7849 19499
rect 7708 19468 7849 19496
rect 7708 19456 7714 19468
rect 7837 19465 7849 19468
rect 7883 19465 7895 19499
rect 9858 19496 9864 19508
rect 9819 19468 9864 19496
rect 7837 19459 7895 19465
rect 9858 19456 9864 19468
rect 9916 19496 9922 19508
rect 11422 19496 11428 19508
rect 9916 19468 11428 19496
rect 9916 19456 9922 19468
rect 11422 19456 11428 19468
rect 11480 19456 11486 19508
rect 13722 19496 13728 19508
rect 13683 19468 13728 19496
rect 13722 19456 13728 19468
rect 13780 19456 13786 19508
rect 5166 19388 5172 19440
rect 5224 19428 5230 19440
rect 8665 19431 8723 19437
rect 8665 19428 8677 19431
rect 5224 19400 8677 19428
rect 5224 19388 5230 19400
rect 8665 19397 8677 19400
rect 8711 19428 8723 19431
rect 10229 19431 10287 19437
rect 10229 19428 10241 19431
rect 8711 19400 10241 19428
rect 8711 19397 8723 19400
rect 8665 19391 8723 19397
rect 10229 19397 10241 19400
rect 10275 19397 10287 19431
rect 10229 19391 10287 19397
rect 934 19320 940 19372
rect 992 19360 998 19372
rect 992 19346 4108 19360
rect 992 19332 4068 19346
rect 992 19320 998 19332
rect 4001 19306 4068 19332
rect 1464 19295 1522 19301
rect 1464 19261 1476 19295
rect 1510 19292 1522 19295
rect 2660 19295 2718 19301
rect 1510 19264 2360 19292
rect 1510 19261 1522 19264
rect 1464 19255 1522 19261
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 2332 19165 2360 19264
rect 2660 19261 2672 19295
rect 2706 19292 2718 19295
rect 2866 19292 2872 19304
rect 2706 19264 2872 19292
rect 2706 19261 2718 19264
rect 2660 19255 2718 19261
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 4062 19294 4068 19306
rect 4120 19294 4126 19346
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 5905 19363 5963 19369
rect 4396 19332 5850 19360
rect 4396 19320 4402 19332
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4212 19264 4257 19292
rect 4212 19252 4218 19264
rect 4430 19252 4436 19304
rect 4488 19292 4494 19304
rect 5166 19292 5172 19304
rect 4488 19264 5172 19292
rect 4488 19252 4494 19264
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19261 5779 19295
rect 5822 19292 5850 19332
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 6730 19360 6736 19372
rect 5951 19332 6736 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 6730 19320 6736 19332
rect 6788 19320 6794 19372
rect 8018 19360 8024 19372
rect 7116 19332 8024 19360
rect 7116 19301 7144 19332
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 6641 19295 6699 19301
rect 6641 19292 6653 19295
rect 5822 19264 6653 19292
rect 5721 19255 5779 19261
rect 6641 19261 6653 19264
rect 6687 19292 6699 19295
rect 7101 19295 7159 19301
rect 7101 19292 7113 19295
rect 6687 19264 7113 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7101 19261 7113 19264
rect 7147 19261 7159 19295
rect 7282 19292 7288 19304
rect 7243 19264 7288 19292
rect 7101 19255 7159 19261
rect 4264 19196 4660 19224
rect 2317 19159 2375 19165
rect 2317 19125 2329 19159
rect 2363 19156 2375 19159
rect 2406 19156 2412 19168
rect 2363 19128 2412 19156
rect 2363 19125 2375 19128
rect 2317 19119 2375 19125
rect 2406 19116 2412 19128
rect 2464 19116 2470 19168
rect 2731 19159 2789 19165
rect 2731 19125 2743 19159
rect 2777 19156 2789 19159
rect 2958 19156 2964 19168
rect 2777 19128 2964 19156
rect 2777 19125 2789 19128
rect 2731 19119 2789 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3418 19156 3424 19168
rect 3379 19128 3424 19156
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 4264 19156 4292 19196
rect 4632 19168 4660 19196
rect 5350 19184 5356 19236
rect 5408 19224 5414 19236
rect 5736 19224 5764 19255
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 8680 19292 8708 19391
rect 9585 19363 9643 19369
rect 9585 19329 9597 19363
rect 9631 19360 9643 19363
rect 9674 19360 9680 19372
rect 9631 19332 9680 19360
rect 9631 19329 9643 19332
rect 9585 19323 9643 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 8849 19295 8907 19301
rect 8849 19292 8861 19295
rect 8680 19264 8861 19292
rect 8849 19261 8861 19264
rect 8895 19261 8907 19295
rect 9306 19292 9312 19304
rect 9267 19264 9312 19292
rect 8849 19255 8907 19261
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 10244 19292 10272 19391
rect 13170 19360 13176 19372
rect 13131 19332 13176 19360
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 10413 19295 10471 19301
rect 10413 19292 10425 19295
rect 10244 19264 10425 19292
rect 10413 19261 10425 19264
rect 10459 19261 10471 19295
rect 10870 19292 10876 19304
rect 10831 19264 10876 19292
rect 10413 19255 10471 19261
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 7300 19224 7328 19252
rect 12802 19224 12808 19236
rect 5408 19196 7328 19224
rect 12763 19196 12808 19224
rect 5408 19184 5414 19196
rect 12802 19184 12808 19196
rect 12860 19184 12866 19236
rect 12894 19184 12900 19236
rect 12952 19224 12958 19236
rect 13722 19224 13728 19236
rect 12952 19196 13728 19224
rect 12952 19184 12958 19196
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 4120 19128 4292 19156
rect 4341 19159 4399 19165
rect 4120 19116 4126 19128
rect 4341 19125 4353 19159
rect 4387 19156 4399 19159
rect 4430 19156 4436 19168
rect 4387 19128 4436 19156
rect 4387 19125 4399 19128
rect 4341 19119 4399 19125
rect 4430 19116 4436 19128
rect 4488 19116 4494 19168
rect 4614 19156 4620 19168
rect 4575 19128 4620 19156
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4856 19128 4997 19156
rect 4856 19116 4862 19128
rect 4985 19125 4997 19128
rect 5031 19125 5043 19159
rect 6270 19156 6276 19168
rect 6231 19128 6276 19156
rect 4985 19119 5043 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 6914 19156 6920 19168
rect 6875 19128 6920 19156
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 8202 19156 8208 19168
rect 8163 19128 8208 19156
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 10686 19156 10692 19168
rect 10647 19128 10692 19156
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 11698 19116 11704 19168
rect 11756 19156 11762 19168
rect 11793 19159 11851 19165
rect 11793 19156 11805 19159
rect 11756 19128 11805 19156
rect 11756 19116 11762 19128
rect 11793 19125 11805 19128
rect 11839 19125 11851 19159
rect 11793 19119 11851 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 5350 18952 5356 18964
rect 5311 18924 5356 18952
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 5721 18955 5779 18961
rect 5721 18952 5733 18955
rect 5500 18924 5733 18952
rect 5500 18912 5506 18924
rect 5721 18921 5733 18924
rect 5767 18952 5779 18955
rect 6914 18952 6920 18964
rect 5767 18924 6920 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 9493 18955 9551 18961
rect 9493 18921 9505 18955
rect 9539 18952 9551 18955
rect 9674 18952 9680 18964
rect 9539 18924 9680 18952
rect 9539 18921 9551 18924
rect 9493 18915 9551 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 12805 18955 12863 18961
rect 12805 18952 12817 18955
rect 12207 18924 12817 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 12805 18921 12817 18924
rect 12851 18952 12863 18955
rect 12894 18952 12900 18964
rect 12851 18924 12900 18952
rect 12851 18921 12863 18924
rect 12805 18915 12863 18921
rect 12894 18912 12900 18924
rect 12952 18912 12958 18964
rect 24762 18952 24768 18964
rect 24723 18924 24768 18952
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 4985 18887 5043 18893
rect 4985 18853 4997 18887
rect 5031 18884 5043 18887
rect 5994 18884 6000 18896
rect 5031 18856 6000 18884
rect 5031 18853 5043 18856
rect 4985 18847 5043 18853
rect 5994 18844 6000 18856
rect 6052 18844 6058 18896
rect 7558 18884 7564 18896
rect 7519 18856 7564 18884
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 8478 18844 8484 18896
rect 8536 18884 8542 18896
rect 10689 18887 10747 18893
rect 10689 18884 10701 18887
rect 8536 18856 10701 18884
rect 8536 18844 8542 18856
rect 10689 18853 10701 18856
rect 10735 18884 10747 18887
rect 10870 18884 10876 18896
rect 10735 18856 10876 18884
rect 10735 18853 10747 18856
rect 10689 18847 10747 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11422 18844 11428 18896
rect 11480 18884 11486 18896
rect 11562 18887 11620 18893
rect 11562 18884 11574 18887
rect 11480 18856 11574 18884
rect 11480 18844 11486 18856
rect 11562 18853 11574 18856
rect 11608 18853 11620 18887
rect 11562 18847 11620 18853
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1762 18816 1768 18828
rect 1443 18788 1768 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1762 18776 1768 18788
rect 1820 18816 1826 18828
rect 2314 18816 2320 18828
rect 1820 18788 2320 18816
rect 1820 18776 1826 18788
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18816 3019 18819
rect 3050 18816 3056 18828
rect 3007 18788 3056 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 3050 18776 3056 18788
rect 3108 18776 3114 18828
rect 4890 18816 4896 18828
rect 4851 18788 4896 18816
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 8168 18788 9689 18816
rect 8168 18776 8174 18788
rect 9677 18785 9689 18788
rect 9723 18816 9735 18819
rect 9858 18816 9864 18828
rect 9723 18788 9864 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 10137 18819 10195 18825
rect 10137 18785 10149 18819
rect 10183 18785 10195 18819
rect 13170 18816 13176 18828
rect 13131 18788 13176 18816
rect 10137 18779 10195 18785
rect 5534 18708 5540 18760
rect 5592 18748 5598 18760
rect 5905 18751 5963 18757
rect 5905 18748 5917 18751
rect 5592 18720 5917 18748
rect 5592 18708 5598 18720
rect 5905 18717 5917 18720
rect 5951 18717 5963 18751
rect 6178 18748 6184 18760
rect 6139 18720 6184 18748
rect 5905 18711 5963 18717
rect 6178 18708 6184 18720
rect 6236 18748 6242 18760
rect 7193 18751 7251 18757
rect 7193 18748 7205 18751
rect 6236 18720 7205 18748
rect 6236 18708 6242 18720
rect 7193 18717 7205 18720
rect 7239 18717 7251 18751
rect 7466 18748 7472 18760
rect 7427 18720 7472 18748
rect 7193 18711 7251 18717
rect 7466 18708 7472 18720
rect 7524 18708 7530 18760
rect 7742 18748 7748 18760
rect 7703 18720 7748 18748
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 9306 18748 9312 18760
rect 8864 18720 9312 18748
rect 3145 18615 3203 18621
rect 3145 18581 3157 18615
rect 3191 18612 3203 18615
rect 5074 18612 5080 18624
rect 3191 18584 5080 18612
rect 3191 18581 3203 18584
rect 3145 18575 3203 18581
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7282 18612 7288 18624
rect 6963 18584 7288 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7282 18572 7288 18584
rect 7340 18612 7346 18624
rect 7834 18612 7840 18624
rect 7340 18584 7840 18612
rect 7340 18572 7346 18584
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 8864 18621 8892 18720
rect 9306 18708 9312 18720
rect 9364 18748 9370 18760
rect 10152 18748 10180 18779
rect 13170 18776 13176 18788
rect 13228 18776 13234 18828
rect 15356 18819 15414 18825
rect 15356 18785 15368 18819
rect 15402 18816 15414 18819
rect 15654 18816 15660 18828
rect 15402 18788 15660 18816
rect 15402 18785 15414 18788
rect 15356 18779 15414 18785
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 24578 18816 24584 18828
rect 24539 18788 24584 18816
rect 24578 18776 24584 18788
rect 24636 18816 24642 18828
rect 25406 18816 25412 18828
rect 24636 18788 25412 18816
rect 24636 18776 24642 18788
rect 25406 18776 25412 18788
rect 25464 18776 25470 18828
rect 9364 18720 10180 18748
rect 10413 18751 10471 18757
rect 9364 18708 9370 18720
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10459 18720 11253 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 11241 18717 11253 18720
rect 11287 18748 11299 18751
rect 11790 18748 11796 18760
rect 11287 18720 11796 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 13872 18720 13917 18748
rect 13872 18708 13878 18720
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 11057 18683 11115 18689
rect 11057 18680 11069 18683
rect 10560 18652 11069 18680
rect 10560 18640 10566 18652
rect 11057 18649 11069 18652
rect 11103 18649 11115 18683
rect 11057 18643 11115 18649
rect 15427 18683 15485 18689
rect 15427 18649 15439 18683
rect 15473 18680 15485 18683
rect 18230 18680 18236 18692
rect 15473 18652 18236 18680
rect 15473 18649 15485 18652
rect 15427 18643 15485 18649
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 8849 18615 8907 18621
rect 8849 18612 8861 18615
rect 8720 18584 8861 18612
rect 8720 18572 8726 18584
rect 8849 18581 8861 18584
rect 8895 18581 8907 18615
rect 8849 18575 8907 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 2038 18408 2044 18420
rect 1999 18380 2044 18408
rect 2038 18368 2044 18380
rect 2096 18368 2102 18420
rect 2314 18408 2320 18420
rect 2275 18380 2320 18408
rect 2314 18368 2320 18380
rect 2372 18368 2378 18420
rect 3050 18368 3056 18420
rect 3108 18408 3114 18420
rect 3421 18411 3479 18417
rect 3421 18408 3433 18411
rect 3108 18380 3433 18408
rect 3108 18368 3114 18380
rect 3421 18377 3433 18380
rect 3467 18408 3479 18411
rect 4154 18408 4160 18420
rect 3467 18380 4160 18408
rect 3467 18377 3479 18380
rect 3421 18371 3479 18377
rect 4154 18368 4160 18380
rect 4212 18408 4218 18420
rect 4798 18408 4804 18420
rect 4212 18380 4804 18408
rect 4212 18368 4218 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 4985 18411 5043 18417
rect 4985 18408 4997 18411
rect 4948 18380 4997 18408
rect 4948 18368 4954 18380
rect 4985 18377 4997 18380
rect 5031 18377 5043 18411
rect 4985 18371 5043 18377
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6181 18411 6239 18417
rect 6181 18408 6193 18411
rect 6052 18380 6193 18408
rect 6052 18368 6058 18380
rect 6181 18377 6193 18380
rect 6227 18377 6239 18411
rect 6181 18371 6239 18377
rect 6825 18411 6883 18417
rect 6825 18377 6837 18411
rect 6871 18408 6883 18411
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 6871 18380 8309 18408
rect 6871 18377 6883 18380
rect 6825 18371 6883 18377
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 9858 18408 9864 18420
rect 9819 18380 9864 18408
rect 8297 18371 8355 18377
rect 4338 18340 4344 18352
rect 4299 18312 4344 18340
rect 4338 18300 4344 18312
rect 4396 18300 4402 18352
rect 7558 18340 7564 18352
rect 6012 18312 7564 18340
rect 5905 18275 5963 18281
rect 5905 18241 5917 18275
rect 5951 18272 5963 18275
rect 6012 18272 6040 18312
rect 7558 18300 7564 18312
rect 7616 18340 7622 18352
rect 7929 18343 7987 18349
rect 7929 18340 7941 18343
rect 7616 18312 7941 18340
rect 7616 18300 7622 18312
rect 7929 18309 7941 18312
rect 7975 18309 7987 18343
rect 7929 18303 7987 18309
rect 5951 18244 6040 18272
rect 5951 18241 5963 18244
rect 5905 18235 5963 18241
rect 6178 18232 6184 18284
rect 6236 18272 6242 18284
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6236 18244 7021 18272
rect 6236 18232 6242 18244
rect 7009 18241 7021 18244
rect 7055 18241 7067 18275
rect 7009 18235 7067 18241
rect 7653 18275 7711 18281
rect 7653 18241 7665 18275
rect 7699 18272 7711 18275
rect 7742 18272 7748 18284
rect 7699 18244 7748 18272
rect 7699 18241 7711 18244
rect 7653 18235 7711 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 2038 18204 2044 18216
rect 1443 18176 2044 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 2038 18164 2044 18176
rect 2096 18164 2102 18216
rect 2498 18204 2504 18216
rect 2462 18176 2504 18204
rect 2498 18164 2504 18176
rect 2556 18213 2562 18216
rect 2556 18207 2610 18213
rect 2556 18173 2564 18207
rect 2598 18204 2610 18207
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2598 18176 2973 18204
rect 2598 18173 2610 18176
rect 2556 18167 2610 18173
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18204 4215 18207
rect 4246 18204 4252 18216
rect 4203 18176 4252 18204
rect 4203 18173 4215 18176
rect 4157 18167 4215 18173
rect 2556 18164 2562 18167
rect 4246 18164 4252 18176
rect 4304 18164 4310 18216
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 4948 18176 5825 18204
rect 4948 18164 4954 18176
rect 5813 18173 5825 18176
rect 5859 18204 5871 18207
rect 6638 18204 6644 18216
rect 5859 18176 6644 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 6638 18164 6644 18176
rect 6696 18164 6702 18216
rect 2639 18139 2697 18145
rect 2639 18105 2651 18139
rect 2685 18136 2697 18139
rect 6825 18139 6883 18145
rect 6825 18136 6837 18139
rect 2685 18108 6837 18136
rect 2685 18105 2697 18108
rect 2639 18099 2697 18105
rect 6825 18105 6837 18108
rect 6871 18105 6883 18139
rect 6825 18099 6883 18105
rect 7098 18096 7104 18148
rect 7156 18136 7162 18148
rect 8312 18136 8340 18371
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 11422 18408 11428 18420
rect 11383 18380 11428 18408
rect 11422 18368 11428 18380
rect 11480 18368 11486 18420
rect 11790 18408 11796 18420
rect 11751 18380 11796 18408
rect 11790 18368 11796 18380
rect 11848 18368 11854 18420
rect 13170 18408 13176 18420
rect 13131 18380 13176 18408
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 25406 18408 25412 18420
rect 25367 18380 25412 18408
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 24578 18300 24584 18352
rect 24636 18340 24642 18352
rect 24719 18343 24777 18349
rect 24719 18340 24731 18343
rect 24636 18312 24731 18340
rect 24636 18300 24642 18312
rect 24719 18309 24731 18312
rect 24765 18309 24777 18343
rect 24719 18303 24777 18309
rect 8754 18232 8760 18284
rect 8812 18272 8818 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 8812 18244 9229 18272
rect 8812 18232 8818 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18272 14703 18275
rect 14829 18275 14887 18281
rect 14829 18272 14841 18275
rect 14691 18244 14841 18272
rect 14691 18241 14703 18244
rect 14645 18235 14703 18241
rect 14829 18241 14841 18244
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 25133 18275 25191 18281
rect 25133 18241 25145 18275
rect 25179 18272 25191 18275
rect 27614 18272 27620 18284
rect 25179 18244 27620 18272
rect 25179 18241 25191 18244
rect 25133 18235 25191 18241
rect 12472 18207 12530 18213
rect 12472 18173 12484 18207
rect 12518 18173 12530 18207
rect 15381 18207 15439 18213
rect 15381 18204 15393 18207
rect 12472 18167 12530 18173
rect 14752 18176 15393 18204
rect 8941 18139 8999 18145
rect 8941 18136 8953 18139
rect 7156 18108 7201 18136
rect 8312 18108 8953 18136
rect 7156 18096 7162 18108
rect 8941 18105 8953 18108
rect 8987 18105 8999 18139
rect 8941 18099 8999 18105
rect 9033 18139 9091 18145
rect 9033 18105 9045 18139
rect 9079 18136 9091 18139
rect 9214 18136 9220 18148
rect 9079 18108 9220 18136
rect 9079 18105 9091 18108
rect 9033 18099 9091 18105
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4614 18068 4620 18080
rect 4304 18040 4620 18068
rect 4304 18028 4310 18040
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 6638 18068 6644 18080
rect 6599 18040 6644 18068
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 8757 18071 8815 18077
rect 8757 18037 8769 18071
rect 8803 18068 8815 18071
rect 9048 18068 9076 18099
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 10042 18096 10048 18148
rect 10100 18136 10106 18148
rect 10502 18136 10508 18148
rect 10100 18108 10508 18136
rect 10100 18096 10106 18108
rect 10502 18096 10508 18108
rect 10560 18096 10566 18148
rect 10597 18139 10655 18145
rect 10597 18105 10609 18139
rect 10643 18105 10655 18139
rect 11146 18136 11152 18148
rect 11107 18108 11152 18136
rect 10597 18099 10655 18105
rect 8803 18040 9076 18068
rect 8803 18037 8815 18040
rect 8757 18031 8815 18037
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 10192 18040 10241 18068
rect 10192 18028 10198 18040
rect 10229 18037 10241 18040
rect 10275 18068 10287 18071
rect 10612 18068 10640 18099
rect 11146 18096 11152 18108
rect 11204 18136 11210 18148
rect 12161 18139 12219 18145
rect 12161 18136 12173 18139
rect 11204 18108 12173 18136
rect 11204 18096 11210 18108
rect 12161 18105 12173 18108
rect 12207 18136 12219 18139
rect 12487 18136 12515 18167
rect 13998 18136 14004 18148
rect 12207 18108 12515 18136
rect 13959 18108 14004 18136
rect 12207 18105 12219 18108
rect 12161 18099 12219 18105
rect 13998 18096 14004 18108
rect 14056 18096 14062 18148
rect 14093 18139 14151 18145
rect 14093 18105 14105 18139
rect 14139 18105 14151 18139
rect 14093 18099 14151 18105
rect 10275 18040 10640 18068
rect 10275 18037 10287 18040
rect 10229 18031 10287 18037
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 12575 18071 12633 18077
rect 12575 18068 12587 18071
rect 11940 18040 12587 18068
rect 11940 18028 11946 18040
rect 12575 18037 12587 18040
rect 12621 18037 12633 18071
rect 12575 18031 12633 18037
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 13504 18040 13829 18068
rect 13504 18028 13510 18040
rect 13817 18037 13829 18040
rect 13863 18068 13875 18071
rect 14108 18068 14136 18099
rect 14752 18068 14780 18176
rect 15381 18173 15393 18176
rect 15427 18204 15439 18207
rect 15565 18207 15623 18213
rect 15565 18204 15577 18207
rect 15427 18176 15577 18204
rect 15427 18173 15439 18176
rect 15381 18167 15439 18173
rect 15565 18173 15577 18176
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 24648 18207 24706 18213
rect 24648 18173 24660 18207
rect 24694 18204 24706 18207
rect 25148 18204 25176 18235
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 24694 18176 25176 18204
rect 24694 18173 24706 18176
rect 24648 18167 24706 18173
rect 15470 18136 15476 18148
rect 15431 18108 15476 18136
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 13863 18040 14780 18068
rect 14829 18071 14887 18077
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 14829 18037 14841 18071
rect 14875 18068 14887 18071
rect 15013 18071 15071 18077
rect 15013 18068 15025 18071
rect 14875 18040 15025 18068
rect 14875 18037 14887 18040
rect 14829 18031 14887 18037
rect 15013 18037 15025 18040
rect 15059 18068 15071 18071
rect 15654 18068 15660 18080
rect 15059 18040 15660 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 4890 17864 4896 17876
rect 4851 17836 4896 17864
rect 4890 17824 4896 17836
rect 4948 17824 4954 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 5592 17836 6469 17864
rect 5592 17824 5598 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 6457 17827 6515 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 11977 17867 12035 17873
rect 11977 17833 11989 17867
rect 12023 17864 12035 17867
rect 12710 17864 12716 17876
rect 12023 17836 12716 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 4982 17756 4988 17808
rect 5040 17796 5046 17808
rect 5629 17799 5687 17805
rect 5629 17796 5641 17799
rect 5040 17768 5641 17796
rect 5040 17756 5046 17768
rect 5629 17765 5641 17768
rect 5675 17796 5687 17799
rect 5994 17796 6000 17808
rect 5675 17768 6000 17796
rect 5675 17765 5687 17768
rect 5629 17759 5687 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 6178 17796 6184 17808
rect 6139 17768 6184 17796
rect 6178 17756 6184 17768
rect 6236 17756 6242 17808
rect 7009 17799 7067 17805
rect 7009 17765 7021 17799
rect 7055 17796 7067 17799
rect 10042 17796 10048 17808
rect 7055 17768 10048 17796
rect 7055 17765 7067 17768
rect 7009 17759 7067 17765
rect 10042 17756 10048 17768
rect 10100 17756 10106 17808
rect 10134 17756 10140 17808
rect 10192 17796 10198 17808
rect 10229 17799 10287 17805
rect 10229 17796 10241 17799
rect 10192 17768 10241 17796
rect 10192 17756 10198 17768
rect 10229 17765 10241 17768
rect 10275 17765 10287 17799
rect 12986 17796 12992 17808
rect 12947 17768 12992 17796
rect 10229 17759 10287 17765
rect 12986 17756 12992 17768
rect 13044 17756 13050 17808
rect 13081 17799 13139 17805
rect 13081 17765 13093 17799
rect 13127 17796 13139 17799
rect 13170 17796 13176 17808
rect 13127 17768 13176 17796
rect 13127 17765 13139 17768
rect 13081 17759 13139 17765
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 15470 17796 15476 17808
rect 15431 17768 15476 17796
rect 15470 17756 15476 17768
rect 15528 17756 15534 17808
rect 2593 17731 2651 17737
rect 2593 17697 2605 17731
rect 2639 17728 2651 17731
rect 2866 17728 2872 17740
rect 2639 17700 2872 17728
rect 2639 17697 2651 17700
rect 2593 17691 2651 17697
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4246 17728 4252 17740
rect 4111 17700 4252 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4246 17688 4252 17700
rect 4304 17688 4310 17740
rect 8018 17728 8024 17740
rect 7979 17700 8024 17728
rect 8018 17688 8024 17700
rect 8076 17688 8082 17740
rect 8478 17728 8484 17740
rect 8439 17700 8484 17728
rect 8478 17688 8484 17700
rect 8536 17688 8542 17740
rect 10318 17728 10324 17740
rect 10279 17700 10324 17728
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17728 11851 17731
rect 11882 17728 11888 17740
rect 11839 17700 11888 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 5537 17663 5595 17669
rect 5537 17660 5549 17663
rect 5224 17632 5549 17660
rect 5224 17620 5230 17632
rect 5537 17629 5549 17632
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17660 8815 17663
rect 11698 17660 11704 17672
rect 8803 17632 11704 17660
rect 8803 17629 8815 17632
rect 8757 17623 8815 17629
rect 11698 17620 11704 17632
rect 11756 17620 11762 17672
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17629 15439 17663
rect 15654 17660 15660 17672
rect 15615 17632 15660 17660
rect 15381 17623 15439 17629
rect 13541 17595 13599 17601
rect 13541 17561 13553 17595
rect 13587 17592 13599 17595
rect 15396 17592 15424 17623
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 15562 17592 15568 17604
rect 13587 17564 13814 17592
rect 15396 17564 15568 17592
rect 13587 17561 13599 17564
rect 13541 17555 13599 17561
rect 1486 17484 1492 17536
rect 1544 17524 1550 17536
rect 1581 17527 1639 17533
rect 1581 17524 1593 17527
rect 1544 17496 1593 17524
rect 1544 17484 1550 17496
rect 1581 17493 1593 17496
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2225 17527 2283 17533
rect 2225 17524 2237 17527
rect 2096 17496 2237 17524
rect 2096 17484 2102 17496
rect 2225 17493 2237 17496
rect 2271 17493 2283 17527
rect 2225 17487 2283 17493
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 4249 17527 4307 17533
rect 4249 17524 4261 17527
rect 4212 17496 4261 17524
rect 4212 17484 4218 17496
rect 4249 17493 4261 17496
rect 4295 17493 4307 17527
rect 5258 17524 5264 17536
rect 5219 17496 5264 17524
rect 4249 17487 4307 17493
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 9861 17527 9919 17533
rect 9861 17524 9873 17527
rect 8720 17496 9873 17524
rect 8720 17484 8726 17496
rect 9861 17493 9873 17496
rect 9907 17493 9919 17527
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 9861 17487 9919 17493
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13786 17524 13814 17564
rect 15562 17552 15568 17564
rect 15620 17552 15626 17604
rect 13998 17524 14004 17536
rect 13786 17496 14004 17524
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 14369 17527 14427 17533
rect 14369 17493 14381 17527
rect 14415 17524 14427 17527
rect 14642 17524 14648 17536
rect 14415 17496 14648 17524
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 14642 17484 14648 17496
rect 14700 17484 14706 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 5994 17280 6000 17332
rect 6052 17320 6058 17332
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 6052 17292 6193 17320
rect 6052 17280 6058 17292
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 6270 17280 6276 17332
rect 6328 17320 6334 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6328 17292 6561 17320
rect 6328 17280 6334 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 6564 17184 6592 17283
rect 6638 17280 6644 17332
rect 6696 17320 6702 17332
rect 7098 17320 7104 17332
rect 6696 17292 7104 17320
rect 6696 17280 6702 17292
rect 7098 17280 7104 17292
rect 7156 17320 7162 17332
rect 7745 17323 7803 17329
rect 7745 17320 7757 17323
rect 7156 17292 7757 17320
rect 7156 17280 7162 17292
rect 7745 17289 7757 17292
rect 7791 17289 7803 17323
rect 10318 17320 10324 17332
rect 10279 17292 10324 17320
rect 7745 17283 7803 17289
rect 10318 17280 10324 17292
rect 10376 17320 10382 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 10376 17292 10609 17320
rect 10376 17280 10382 17292
rect 10597 17289 10609 17292
rect 10643 17320 10655 17323
rect 10962 17320 10968 17332
rect 10643 17292 10968 17320
rect 10643 17289 10655 17292
rect 10597 17283 10655 17289
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 11882 17320 11888 17332
rect 11843 17292 11888 17320
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 14093 17323 14151 17329
rect 14093 17320 14105 17323
rect 13872 17292 14105 17320
rect 13872 17280 13878 17292
rect 14093 17289 14105 17292
rect 14139 17320 14151 17323
rect 14458 17320 14464 17332
rect 14139 17292 14464 17320
rect 14139 17289 14151 17292
rect 14093 17283 14151 17289
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 15381 17323 15439 17329
rect 15381 17289 15393 17323
rect 15427 17320 15439 17323
rect 15470 17320 15476 17332
rect 15427 17292 15476 17320
rect 15427 17289 15439 17292
rect 15381 17283 15439 17289
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 13170 17212 13176 17264
rect 13228 17252 13234 17264
rect 13725 17255 13783 17261
rect 13725 17252 13737 17255
rect 13228 17224 13737 17252
rect 13228 17212 13234 17224
rect 13725 17221 13737 17224
rect 13771 17221 13783 17255
rect 13725 17215 13783 17221
rect 9214 17184 9220 17196
rect 4172 17156 5304 17184
rect 6564 17156 7189 17184
rect 9175 17156 9220 17184
rect 1486 17076 1492 17128
rect 1544 17116 1550 17128
rect 1673 17119 1731 17125
rect 1673 17116 1685 17119
rect 1544 17088 1685 17116
rect 1544 17076 1550 17088
rect 1673 17085 1685 17088
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 3605 17119 3663 17125
rect 3605 17085 3617 17119
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17048 3571 17051
rect 3620 17048 3648 17079
rect 3694 17076 3700 17128
rect 3752 17116 3758 17128
rect 4172 17125 4200 17156
rect 5276 17128 5304 17156
rect 4157 17119 4215 17125
rect 4157 17116 4169 17119
rect 3752 17088 4169 17116
rect 3752 17076 3758 17088
rect 4157 17085 4169 17088
rect 4203 17085 4215 17119
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 4157 17079 4215 17085
rect 5092 17088 5181 17116
rect 3878 17048 3884 17060
rect 3559 17020 3884 17048
rect 3559 17017 3571 17020
rect 3513 17011 3571 17017
rect 3878 17008 3884 17020
rect 3936 17008 3942 17060
rect 4338 17048 4344 17060
rect 4299 17020 4344 17048
rect 4338 17008 4344 17020
rect 4396 17008 4402 17060
rect 5092 16992 5120 17088
rect 5169 17085 5181 17088
rect 5215 17085 5227 17119
rect 5169 17079 5227 17085
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 5721 17119 5779 17125
rect 5721 17116 5733 17119
rect 5316 17088 5733 17116
rect 5316 17076 5322 17088
rect 5721 17085 5733 17088
rect 5767 17085 5779 17119
rect 5721 17079 5779 17085
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 6822 17116 6828 17128
rect 5951 17088 6828 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 5736 17048 5764 17079
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6086 17048 6092 17060
rect 5736 17020 6092 17048
rect 6086 17008 6092 17020
rect 6144 17008 6150 17060
rect 7161 17057 7189 17156
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 11146 17184 11152 17196
rect 11107 17156 11152 17184
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 13998 17144 14004 17196
rect 14056 17184 14062 17196
rect 14645 17187 14703 17193
rect 14645 17184 14657 17187
rect 14056 17156 14657 17184
rect 14056 17144 14062 17156
rect 14645 17153 14657 17156
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 9125 17119 9183 17125
rect 9125 17116 9137 17119
rect 8352 17088 9137 17116
rect 8352 17076 8358 17088
rect 9125 17085 9137 17088
rect 9171 17116 9183 17119
rect 9858 17116 9864 17128
rect 9171 17088 9864 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 12526 17116 12532 17128
rect 12487 17088 12532 17116
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 7146 17051 7204 17057
rect 7146 17017 7158 17051
rect 7192 17017 7204 17051
rect 7146 17011 7204 17017
rect 8754 17008 8760 17060
rect 8812 17048 8818 17060
rect 10870 17048 10876 17060
rect 8812 17020 10876 17048
rect 8812 17008 8818 17020
rect 10870 17008 10876 17020
rect 10928 17008 10934 17060
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 12850 17051 12908 17057
rect 12850 17048 12862 17051
rect 11020 17020 11065 17048
rect 12176 17020 12862 17048
rect 11020 17008 11026 17020
rect 12176 16992 12204 17020
rect 12850 17017 12862 17020
rect 12896 17017 12908 17051
rect 12850 17011 12908 17017
rect 14369 17051 14427 17057
rect 14369 17017 14381 17051
rect 14415 17017 14427 17051
rect 14369 17011 14427 17017
rect 1854 16980 1860 16992
rect 1815 16952 1860 16980
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 2685 16983 2743 16989
rect 2685 16949 2697 16983
rect 2731 16980 2743 16983
rect 2866 16980 2872 16992
rect 2731 16952 2872 16980
rect 2731 16949 2743 16952
rect 2685 16943 2743 16949
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 4246 16940 4252 16992
rect 4304 16980 4310 16992
rect 4617 16983 4675 16989
rect 4617 16980 4629 16983
rect 4304 16952 4629 16980
rect 4304 16940 4310 16952
rect 4617 16949 4629 16952
rect 4663 16949 4675 16983
rect 5074 16980 5080 16992
rect 5035 16952 5080 16980
rect 4617 16943 4675 16949
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 8018 16980 8024 16992
rect 7340 16952 8024 16980
rect 7340 16940 7346 16952
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 8478 16980 8484 16992
rect 8439 16952 8484 16980
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 12158 16980 12164 16992
rect 12119 16952 12164 16980
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 14384 16980 14412 17011
rect 14458 17008 14464 17060
rect 14516 17048 14522 17060
rect 14516 17020 14561 17048
rect 14516 17008 14522 17020
rect 14642 16980 14648 16992
rect 14384 16952 14648 16980
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 15654 16980 15660 16992
rect 15615 16952 15660 16980
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3694 16776 3700 16788
rect 3655 16748 3700 16776
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 5166 16776 5172 16788
rect 5127 16748 5172 16776
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 5994 16736 6000 16788
rect 6052 16776 6058 16788
rect 6181 16779 6239 16785
rect 6181 16776 6193 16779
rect 6052 16748 6193 16776
rect 6052 16736 6058 16748
rect 6181 16745 6193 16748
rect 6227 16745 6239 16779
rect 6822 16776 6828 16788
rect 6783 16748 6828 16776
rect 6181 16739 6239 16745
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7009 16779 7067 16785
rect 7009 16745 7021 16779
rect 7055 16776 7067 16779
rect 7466 16776 7472 16788
rect 7055 16748 7472 16776
rect 7055 16745 7067 16748
rect 7009 16739 7067 16745
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 10597 16779 10655 16785
rect 10597 16745 10609 16779
rect 10643 16776 10655 16779
rect 10962 16776 10968 16788
rect 10643 16748 10968 16776
rect 10643 16745 10655 16748
rect 10597 16739 10655 16745
rect 10962 16736 10968 16748
rect 11020 16736 11026 16788
rect 12897 16779 12955 16785
rect 12897 16745 12909 16779
rect 12943 16776 12955 16779
rect 13170 16776 13176 16788
rect 12943 16748 13176 16776
rect 12943 16745 12955 16748
rect 12897 16739 12955 16745
rect 13170 16736 13176 16748
rect 13228 16736 13234 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 13786 16748 15393 16776
rect 5350 16668 5356 16720
rect 5408 16708 5414 16720
rect 5623 16711 5681 16717
rect 5623 16708 5635 16711
rect 5408 16680 5635 16708
rect 5408 16668 5414 16680
rect 5623 16677 5635 16680
rect 5669 16708 5681 16711
rect 6270 16708 6276 16720
rect 5669 16680 6276 16708
rect 5669 16677 5681 16680
rect 5623 16671 5681 16677
rect 6270 16668 6276 16680
rect 6328 16708 6334 16720
rect 6546 16708 6552 16720
rect 6328 16680 6552 16708
rect 6328 16668 6334 16680
rect 6546 16668 6552 16680
rect 6604 16668 6610 16720
rect 7929 16711 7987 16717
rect 7929 16677 7941 16711
rect 7975 16708 7987 16711
rect 8205 16711 8263 16717
rect 8205 16708 8217 16711
rect 7975 16680 8217 16708
rect 7975 16677 7987 16680
rect 7929 16671 7987 16677
rect 8205 16677 8217 16680
rect 8251 16708 8263 16711
rect 8294 16708 8300 16720
rect 8251 16680 8300 16708
rect 8251 16677 8263 16680
rect 8205 16671 8263 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 8754 16708 8760 16720
rect 8715 16680 8760 16708
rect 8754 16668 8760 16680
rect 8812 16668 8818 16720
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 9998 16711 10056 16717
rect 9998 16708 10010 16711
rect 9640 16680 10010 16708
rect 9640 16668 9646 16680
rect 9998 16677 10010 16680
rect 10044 16677 10056 16711
rect 10870 16708 10876 16720
rect 10831 16680 10876 16708
rect 9998 16671 10056 16677
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 12158 16668 12164 16720
rect 12216 16708 12222 16720
rect 12298 16711 12356 16717
rect 12298 16708 12310 16711
rect 12216 16680 12310 16708
rect 12216 16668 12222 16680
rect 12298 16677 12310 16680
rect 12344 16677 12356 16711
rect 12298 16671 12356 16677
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 1578 16640 1584 16652
rect 1510 16612 1584 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2958 16640 2964 16652
rect 2919 16612 2964 16640
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3602 16600 3608 16652
rect 3660 16640 3666 16652
rect 4100 16643 4158 16649
rect 4100 16640 4112 16643
rect 3660 16612 4112 16640
rect 3660 16600 3666 16612
rect 4100 16609 4112 16612
rect 4146 16609 4158 16643
rect 4100 16603 4158 16609
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 5261 16643 5319 16649
rect 5261 16640 5273 16643
rect 4396 16612 5273 16640
rect 4396 16600 4402 16612
rect 5261 16609 5273 16612
rect 5307 16640 5319 16643
rect 5442 16640 5448 16652
rect 5307 16612 5448 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 12986 16600 12992 16652
rect 13044 16640 13050 16652
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 13044 16612 13185 16640
rect 13044 16600 13050 16612
rect 13173 16609 13185 16612
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 4614 16572 4620 16584
rect 3191 16544 4620 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 8113 16575 8171 16581
rect 8113 16572 8125 16575
rect 7484 16544 8125 16572
rect 3510 16464 3516 16516
rect 3568 16504 3574 16516
rect 5166 16504 5172 16516
rect 3568 16476 5172 16504
rect 3568 16464 3574 16476
rect 5166 16464 5172 16476
rect 5224 16464 5230 16516
rect 1535 16439 1593 16445
rect 1535 16405 1547 16439
rect 1581 16436 1593 16439
rect 1670 16436 1676 16448
rect 1581 16408 1676 16436
rect 1581 16405 1593 16408
rect 1535 16399 1593 16405
rect 1670 16396 1676 16408
rect 1728 16396 1734 16448
rect 1946 16436 1952 16448
rect 1907 16408 1952 16436
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 4203 16439 4261 16445
rect 4203 16436 4215 16439
rect 2832 16408 4215 16436
rect 2832 16396 2838 16408
rect 4203 16405 4215 16408
rect 4249 16405 4261 16439
rect 4203 16399 4261 16405
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7484 16445 7512 16544
rect 8113 16541 8125 16544
rect 8159 16541 8171 16575
rect 9674 16572 9680 16584
rect 9635 16544 9680 16572
rect 8113 16535 8171 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 11974 16572 11980 16584
rect 11935 16544 11980 16572
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 13786 16572 13814 16748
rect 15381 16745 15393 16748
rect 15427 16745 15439 16779
rect 15381 16739 15439 16745
rect 13909 16711 13967 16717
rect 13909 16677 13921 16711
rect 13955 16708 13967 16711
rect 15654 16708 15660 16720
rect 13955 16680 15660 16708
rect 13955 16677 13967 16680
rect 13909 16671 13967 16677
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 15562 16640 15568 16652
rect 15523 16612 15568 16640
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15749 16643 15807 16649
rect 15749 16609 15761 16643
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 12584 16544 13814 16572
rect 12584 16532 12590 16544
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 15764 16572 15792 16603
rect 15344 16544 15792 16572
rect 15344 16532 15350 16544
rect 7469 16439 7527 16445
rect 7469 16436 7481 16439
rect 7156 16408 7481 16436
rect 7156 16396 7162 16408
rect 7469 16405 7481 16408
rect 7515 16405 7527 16439
rect 7469 16399 7527 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2958 16232 2964 16244
rect 2919 16204 2964 16232
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3602 16232 3608 16244
rect 3563 16204 3608 16232
rect 3602 16192 3608 16204
rect 3660 16192 3666 16244
rect 5350 16232 5356 16244
rect 5311 16204 5356 16232
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 9309 16235 9367 16241
rect 9309 16201 9321 16235
rect 9355 16232 9367 16235
rect 9674 16232 9680 16244
rect 9355 16204 9680 16232
rect 9355 16201 9367 16204
rect 9309 16195 9367 16201
rect 9674 16192 9680 16204
rect 9732 16232 9738 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 9732 16204 11345 16232
rect 9732 16192 9738 16204
rect 11333 16201 11345 16204
rect 11379 16201 11391 16235
rect 11333 16195 11391 16201
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 12621 16235 12679 16241
rect 12621 16232 12633 16235
rect 12032 16204 12633 16232
rect 12032 16192 12038 16204
rect 12621 16201 12633 16204
rect 12667 16232 12679 16235
rect 12667 16204 13814 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 9858 16124 9864 16176
rect 9916 16164 9922 16176
rect 11057 16167 11115 16173
rect 11057 16164 11069 16167
rect 9916 16136 11069 16164
rect 9916 16124 9922 16136
rect 11057 16133 11069 16136
rect 11103 16133 11115 16167
rect 11057 16127 11115 16133
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 7423 16068 8800 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 8772 16040 8800 16068
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 9677 16099 9735 16105
rect 9677 16096 9689 16099
rect 9640 16068 9689 16096
rect 9640 16056 9646 16068
rect 9677 16065 9689 16068
rect 9723 16096 9735 16099
rect 13265 16099 13323 16105
rect 9723 16068 9996 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 1946 16028 1952 16040
rect 1907 16000 1952 16028
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 4065 16031 4123 16037
rect 4065 15997 4077 16031
rect 4111 16028 4123 16031
rect 4246 16028 4252 16040
rect 4111 16000 4252 16028
rect 4111 15997 4123 16000
rect 4065 15991 4123 15997
rect 4246 15988 4252 16000
rect 4304 15988 4310 16040
rect 4890 16028 4896 16040
rect 4851 16000 4896 16028
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 15997 8263 16031
rect 8754 16028 8760 16040
rect 8715 16000 8760 16028
rect 8205 15991 8263 15997
rect 2222 15920 2228 15972
rect 2280 15960 2286 15972
rect 5721 15963 5779 15969
rect 5721 15960 5733 15963
rect 2280 15932 5733 15960
rect 2280 15920 2286 15932
rect 5721 15929 5733 15932
rect 5767 15929 5779 15963
rect 5721 15923 5779 15929
rect 7374 15920 7380 15972
rect 7432 15960 7438 15972
rect 8021 15963 8079 15969
rect 8021 15960 8033 15963
rect 7432 15932 8033 15960
rect 7432 15920 7438 15932
rect 8021 15929 8033 15932
rect 8067 15960 8079 15963
rect 8220 15960 8248 15991
rect 8754 15988 8760 16000
rect 8812 15988 8818 16040
rect 9033 16031 9091 16037
rect 9033 15997 9045 16031
rect 9079 16028 9091 16031
rect 9858 16028 9864 16040
rect 9079 16000 9864 16028
rect 9079 15997 9091 16000
rect 9033 15991 9091 15997
rect 8067 15932 8248 15960
rect 8067 15929 8079 15932
rect 8021 15923 8079 15929
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 2130 15892 2136 15904
rect 2091 15864 2136 15892
rect 2130 15852 2136 15864
rect 2188 15852 2194 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7745 15895 7803 15901
rect 7745 15861 7757 15895
rect 7791 15892 7803 15895
rect 9048 15892 9076 15991
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 9968 15960 9996 16068
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13538 16096 13544 16108
rect 13311 16068 13544 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 13786 16096 13814 16204
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 13786 16068 15485 16096
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 10134 16028 10140 16040
rect 10095 16000 10140 16028
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 16028 14887 16031
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14875 16000 14933 16028
rect 14875 15997 14887 16000
rect 14829 15991 14887 15997
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 10458 15963 10516 15969
rect 10458 15960 10470 15963
rect 9968 15932 10470 15960
rect 10458 15929 10470 15932
rect 10504 15960 10516 15963
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 10504 15932 11989 15960
rect 10504 15929 10516 15932
rect 10458 15923 10516 15929
rect 11977 15929 11989 15932
rect 12023 15960 12035 15963
rect 12158 15960 12164 15972
rect 12023 15932 12164 15960
rect 12023 15929 12035 15932
rect 11977 15923 12035 15929
rect 12158 15920 12164 15932
rect 12216 15960 12222 15972
rect 12894 15960 12900 15972
rect 12216 15932 12900 15960
rect 12216 15920 12222 15932
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 13449 15963 13507 15969
rect 13449 15929 13461 15963
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 7791 15864 9076 15892
rect 7791 15861 7803 15864
rect 7745 15855 7803 15861
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13464 15892 13492 15923
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 14090 15960 14096 15972
rect 13596 15932 13641 15960
rect 14051 15932 14096 15960
rect 13596 15920 13602 15932
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 14936 15960 14964 15991
rect 15286 15988 15292 16040
rect 15344 16028 15350 16040
rect 24670 16037 24676 16040
rect 15381 16031 15439 16037
rect 15381 16028 15393 16031
rect 15344 16000 15393 16028
rect 15344 15988 15350 16000
rect 15381 15997 15393 16000
rect 15427 15997 15439 16031
rect 24648 16031 24676 16037
rect 24648 16028 24660 16031
rect 24583 16000 24660 16028
rect 15381 15991 15439 15997
rect 24648 15997 24660 16000
rect 24728 16028 24734 16040
rect 25041 16031 25099 16037
rect 25041 16028 25053 16031
rect 24728 16000 25053 16028
rect 24648 15991 24676 15997
rect 24670 15988 24676 15991
rect 24728 15988 24734 16000
rect 25041 15997 25053 16000
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 15470 15960 15476 15972
rect 14936 15932 15476 15960
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 18414 15920 18420 15972
rect 18472 15960 18478 15972
rect 20714 15960 20720 15972
rect 18472 15932 20720 15960
rect 18472 15920 18478 15932
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 13412 15864 13492 15892
rect 13412 15852 13418 15864
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 14332 15864 14381 15892
rect 14332 15852 14338 15864
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 14369 15855 14427 15861
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 15933 15895 15991 15901
rect 15933 15892 15945 15895
rect 15620 15864 15945 15892
rect 15620 15852 15626 15864
rect 15933 15861 15945 15864
rect 15979 15861 15991 15895
rect 15933 15855 15991 15861
rect 18598 15852 18604 15904
rect 18656 15892 18662 15904
rect 24719 15895 24777 15901
rect 24719 15892 24731 15895
rect 18656 15864 24731 15892
rect 18656 15852 18662 15864
rect 24719 15861 24731 15864
rect 24765 15861 24777 15895
rect 24719 15855 24777 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1118 15648 1124 15700
rect 1176 15688 1182 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1176 15660 1777 15688
rect 1176 15648 1182 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 1765 15651 1823 15657
rect 1780 15484 1808 15651
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 4028 15660 4261 15688
rect 4028 15648 4034 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 4249 15651 4307 15657
rect 2130 15620 2136 15632
rect 2091 15592 2136 15620
rect 2130 15580 2136 15592
rect 2188 15580 2194 15632
rect 4264 15620 4292 15651
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 8757 15691 8815 15697
rect 8757 15657 8769 15691
rect 8803 15688 8815 15691
rect 10134 15688 10140 15700
rect 8803 15660 10140 15688
rect 8803 15657 8815 15660
rect 8757 15651 8815 15657
rect 10134 15648 10140 15660
rect 10192 15688 10198 15700
rect 10505 15691 10563 15697
rect 10505 15688 10517 15691
rect 10192 15660 10517 15688
rect 10192 15648 10198 15660
rect 10505 15657 10517 15660
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 13596 15660 15424 15688
rect 13596 15648 13602 15660
rect 4525 15623 4583 15629
rect 4525 15620 4537 15623
rect 4264 15592 4537 15620
rect 4525 15589 4537 15592
rect 4571 15589 4583 15623
rect 4525 15583 4583 15589
rect 4614 15580 4620 15632
rect 4672 15620 4678 15632
rect 4672 15592 4717 15620
rect 4672 15580 4678 15592
rect 4890 15580 4896 15632
rect 4948 15620 4954 15632
rect 4948 15592 8892 15620
rect 4948 15580 4954 15592
rect 6362 15552 6368 15564
rect 6323 15524 6368 15552
rect 6362 15512 6368 15524
rect 6420 15512 6426 15564
rect 7374 15512 7380 15564
rect 7432 15552 7438 15564
rect 7653 15555 7711 15561
rect 7653 15552 7665 15555
rect 7432 15524 7665 15552
rect 7432 15512 7438 15524
rect 7653 15521 7665 15524
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 7742 15512 7748 15564
rect 7800 15552 7806 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 7800 15524 8493 15552
rect 7800 15512 7806 15524
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 8481 15515 8539 15521
rect 8665 15555 8723 15561
rect 8665 15521 8677 15555
rect 8711 15552 8723 15555
rect 8754 15552 8760 15564
rect 8711 15524 8760 15552
rect 8711 15521 8723 15524
rect 8665 15515 8723 15521
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 8864 15552 8892 15592
rect 9122 15580 9128 15632
rect 9180 15620 9186 15632
rect 9309 15623 9367 15629
rect 9309 15620 9321 15623
rect 9180 15592 9321 15620
rect 9180 15580 9186 15592
rect 9309 15589 9321 15592
rect 9355 15589 9367 15623
rect 9309 15583 9367 15589
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 9640 15592 10241 15620
rect 9640 15580 9646 15592
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 10229 15583 10287 15589
rect 11333 15623 11391 15629
rect 11333 15589 11345 15623
rect 11379 15620 11391 15623
rect 11422 15620 11428 15632
rect 11379 15592 11428 15620
rect 11379 15589 11391 15592
rect 11333 15583 11391 15589
rect 11422 15580 11428 15592
rect 11480 15580 11486 15632
rect 13814 15580 13820 15632
rect 13872 15620 13878 15632
rect 15289 15623 15347 15629
rect 15289 15620 15301 15623
rect 13872 15592 15301 15620
rect 13872 15580 13878 15592
rect 15289 15589 15301 15592
rect 15335 15589 15347 15623
rect 15289 15583 15347 15589
rect 15396 15564 15424 15660
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 8864 15524 9689 15552
rect 9677 15521 9689 15524
rect 9723 15552 9735 15555
rect 10318 15552 10324 15564
rect 9723 15524 10324 15552
rect 9723 15521 9735 15524
rect 9677 15515 9735 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 15378 15552 15384 15564
rect 15291 15524 15384 15552
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1780 15456 2053 15484
rect 2041 15453 2053 15456
rect 2087 15453 2099 15487
rect 5166 15484 5172 15496
rect 5127 15456 5172 15484
rect 2041 15447 2099 15453
rect 5166 15444 5172 15456
rect 5224 15444 5230 15496
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5408 15456 6101 15484
rect 5408 15444 5414 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 11238 15484 11244 15496
rect 11199 15456 11244 15484
rect 6089 15447 6147 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 11514 15484 11520 15496
rect 11475 15456 11520 15484
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13722 15484 13728 15496
rect 13127 15456 13728 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14090 15484 14096 15496
rect 14051 15456 14096 15484
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 2590 15416 2596 15428
rect 2551 15388 2596 15416
rect 2590 15376 2596 15388
rect 2648 15376 2654 15428
rect 14274 15376 14280 15428
rect 14332 15416 14338 15428
rect 14921 15419 14979 15425
rect 14921 15416 14933 15419
rect 14332 15388 14933 15416
rect 14332 15376 14338 15388
rect 14921 15385 14933 15388
rect 14967 15416 14979 15419
rect 15286 15416 15292 15428
rect 14967 15388 15292 15416
rect 14967 15385 14979 15388
rect 14921 15379 14979 15385
rect 15286 15376 15292 15388
rect 15344 15376 15350 15428
rect 24762 15416 24768 15428
rect 24723 15388 24768 15416
rect 24762 15376 24768 15388
rect 24820 15376 24826 15428
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 7650 15348 7656 15360
rect 7515 15320 7656 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 9858 15348 9864 15360
rect 9819 15320 9864 15348
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 13354 15348 13360 15360
rect 13315 15320 13360 15348
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2130 15144 2136 15156
rect 1995 15116 2136 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2958 15104 2964 15156
rect 3016 15144 3022 15156
rect 3329 15147 3387 15153
rect 3329 15144 3341 15147
rect 3016 15116 3341 15144
rect 3016 15104 3022 15116
rect 3329 15113 3341 15116
rect 3375 15144 3387 15147
rect 3421 15147 3479 15153
rect 3421 15144 3433 15147
rect 3375 15116 3433 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3421 15113 3433 15116
rect 3467 15113 3479 15147
rect 4614 15144 4620 15156
rect 4575 15116 4620 15144
rect 3421 15107 3479 15113
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 4939 15116 6561 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 6549 15113 6561 15116
rect 6595 15144 6607 15147
rect 7742 15144 7748 15156
rect 6595 15116 7748 15144
rect 6595 15113 6607 15116
rect 6549 15107 6607 15113
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 9125 15147 9183 15153
rect 9125 15144 9137 15147
rect 8812 15116 9137 15144
rect 8812 15104 8818 15116
rect 9125 15113 9137 15116
rect 9171 15113 9183 15147
rect 10318 15144 10324 15156
rect 10279 15116 10324 15144
rect 9125 15107 9183 15113
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15144 13783 15147
rect 13814 15144 13820 15156
rect 13771 15116 13820 15144
rect 13771 15113 13783 15116
rect 13725 15107 13783 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 15378 15144 15384 15156
rect 15339 15116 15384 15144
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 23799 15147 23857 15153
rect 23799 15113 23811 15147
rect 23845 15144 23857 15147
rect 24670 15144 24676 15156
rect 23845 15116 24676 15144
rect 23845 15113 23857 15116
rect 23799 15107 23857 15113
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 3053 15079 3111 15085
rect 3053 15076 3065 15079
rect 2148 15048 3065 15076
rect 1670 14968 1676 15020
rect 1728 15008 1734 15020
rect 2148 15017 2176 15048
rect 3053 15045 3065 15048
rect 3099 15045 3111 15079
rect 3053 15039 3111 15045
rect 4249 15079 4307 15085
rect 4249 15045 4261 15079
rect 4295 15076 4307 15079
rect 5166 15076 5172 15088
rect 4295 15048 5172 15076
rect 4295 15045 4307 15048
rect 4249 15039 4307 15045
rect 5166 15036 5172 15048
rect 5224 15036 5230 15088
rect 8202 15076 8208 15088
rect 8163 15048 8208 15076
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 11514 15036 11520 15088
rect 11572 15076 11578 15088
rect 11572 15048 12848 15076
rect 11572 15036 11578 15048
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 1728 14980 2145 15008
rect 1728 14968 1734 14980
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2133 14971 2191 14977
rect 2590 14968 2596 14980
rect 2648 15008 2654 15020
rect 3694 15008 3700 15020
rect 2648 14980 3700 15008
rect 2648 14968 2654 14980
rect 3694 14968 3700 14980
rect 3752 14968 3758 15020
rect 4154 14968 4160 15020
rect 4212 15008 4218 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4212 14980 4905 15008
rect 4212 14968 4218 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 5258 15008 5264 15020
rect 5171 14980 5264 15008
rect 4893 14971 4951 14977
rect 5258 14968 5264 14980
rect 5316 15008 5322 15020
rect 6822 15008 6828 15020
rect 5316 14980 6828 15008
rect 5316 14968 5322 14980
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 7024 14980 9689 15008
rect 5905 14943 5963 14949
rect 5905 14909 5917 14943
rect 5951 14940 5963 14943
rect 5994 14940 6000 14952
rect 5951 14912 6000 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 5994 14900 6000 14912
rect 6052 14940 6058 14952
rect 7024 14940 7052 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11793 15011 11851 15017
rect 11793 15008 11805 15011
rect 11296 14980 11805 15008
rect 11296 14968 11302 14980
rect 11793 14977 11805 14980
rect 11839 15008 11851 15011
rect 12710 15008 12716 15020
rect 11839 14980 12716 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12820 15017 12848 15048
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 14977 12863 15011
rect 12805 14971 12863 14977
rect 7650 14940 7656 14952
rect 6052 14912 7052 14940
rect 7611 14912 7656 14940
rect 6052 14900 6058 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 8202 14940 8208 14952
rect 7800 14912 8208 14940
rect 7800 14900 7806 14912
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8386 14940 8392 14952
rect 8299 14912 8392 14940
rect 8386 14900 8392 14912
rect 8444 14940 8450 14952
rect 8754 14940 8760 14952
rect 8444 14912 8760 14940
rect 8444 14900 8450 14912
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15344 14912 15577 14940
rect 15344 14900 15350 14912
rect 15565 14909 15577 14912
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16577 14943 16635 14949
rect 16577 14940 16589 14943
rect 16255 14912 16589 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16577 14909 16589 14912
rect 16623 14909 16635 14943
rect 16577 14903 16635 14909
rect 23728 14943 23786 14949
rect 23728 14909 23740 14943
rect 23774 14940 23786 14943
rect 24118 14940 24124 14952
rect 23774 14912 24124 14940
rect 23774 14909 23786 14912
rect 23728 14903 23786 14909
rect 1946 14832 1952 14884
rect 2004 14872 2010 14884
rect 2225 14875 2283 14881
rect 2225 14872 2237 14875
rect 2004 14844 2237 14872
rect 2004 14832 2010 14844
rect 2225 14841 2237 14844
rect 2271 14841 2283 14875
rect 2225 14835 2283 14841
rect 3329 14875 3387 14881
rect 3329 14841 3341 14875
rect 3375 14872 3387 14875
rect 3786 14872 3792 14884
rect 3375 14844 3792 14872
rect 3375 14841 3387 14844
rect 3329 14835 3387 14841
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 6270 14872 6276 14884
rect 5408 14844 5453 14872
rect 6183 14844 6276 14872
rect 5408 14832 5414 14844
rect 6270 14832 6276 14844
rect 6328 14872 6334 14884
rect 8404 14872 8432 14900
rect 6328 14844 8432 14872
rect 6328 14832 6334 14844
rect 9122 14832 9128 14884
rect 9180 14872 9186 14884
rect 9401 14875 9459 14881
rect 9401 14872 9413 14875
rect 9180 14844 9413 14872
rect 9180 14832 9186 14844
rect 9401 14841 9413 14844
rect 9447 14841 9459 14875
rect 9401 14835 9459 14841
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 10873 14875 10931 14881
rect 9548 14844 9593 14872
rect 9548 14832 9554 14844
rect 10873 14841 10885 14875
rect 10919 14872 10931 14875
rect 12526 14872 12532 14884
rect 10919 14844 12532 14872
rect 10919 14841 10931 14844
rect 10873 14835 10931 14841
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 12621 14875 12679 14881
rect 12621 14841 12633 14875
rect 12667 14872 12679 14875
rect 12802 14872 12808 14884
rect 12667 14844 12808 14872
rect 12667 14841 12679 14844
rect 12621 14835 12679 14841
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5368 14804 5396 14832
rect 5123 14776 5396 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 6788 14776 7205 14804
rect 6788 14764 6794 14776
rect 7193 14773 7205 14776
rect 7239 14804 7251 14807
rect 7374 14804 7380 14816
rect 7239 14776 7380 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8757 14807 8815 14813
rect 8757 14804 8769 14807
rect 8260 14776 8769 14804
rect 8260 14764 8266 14776
rect 8757 14773 8769 14776
rect 8803 14804 8815 14807
rect 8938 14804 8944 14816
rect 8803 14776 8944 14804
rect 8803 14773 8815 14776
rect 8757 14767 8815 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 11422 14804 11428 14816
rect 11383 14776 11428 14804
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 12636 14804 12664 14835
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 14090 14872 14096 14884
rect 14051 14844 14096 14872
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 14185 14875 14243 14881
rect 14185 14841 14197 14875
rect 14231 14841 14243 14875
rect 14185 14835 14243 14841
rect 14737 14875 14795 14881
rect 14737 14841 14749 14875
rect 14783 14872 14795 14875
rect 14826 14872 14832 14884
rect 14783 14844 14832 14872
rect 14783 14841 14795 14844
rect 14737 14835 14795 14841
rect 12299 14776 12664 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 13998 14764 14004 14816
rect 14056 14804 14062 14816
rect 14200 14804 14228 14835
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 16224 14804 16252 14903
rect 24118 14900 24124 14912
rect 24176 14900 24182 14952
rect 14056 14776 16252 14804
rect 14056 14764 14062 14776
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 2004 14572 2053 14600
rect 2004 14560 2010 14572
rect 2041 14569 2053 14572
rect 2087 14600 2099 14603
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 2087 14572 3157 14600
rect 2087 14569 2099 14572
rect 2041 14563 2099 14569
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3694 14600 3700 14612
rect 3655 14572 3700 14600
rect 3145 14563 3203 14569
rect 3694 14560 3700 14572
rect 3752 14560 3758 14612
rect 3786 14560 3792 14612
rect 3844 14600 3850 14612
rect 4985 14603 5043 14609
rect 4985 14600 4997 14603
rect 3844 14572 4997 14600
rect 3844 14560 3850 14572
rect 4985 14569 4997 14572
rect 5031 14569 5043 14603
rect 5258 14600 5264 14612
rect 5219 14572 5264 14600
rect 4985 14563 5043 14569
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 6362 14600 6368 14612
rect 6323 14572 6368 14600
rect 6362 14560 6368 14572
rect 6420 14560 6426 14612
rect 6733 14603 6791 14609
rect 6733 14569 6745 14603
rect 6779 14600 6791 14603
rect 6822 14600 6828 14612
rect 6779 14572 6828 14600
rect 6779 14569 6791 14572
rect 6733 14563 6791 14569
rect 6822 14560 6828 14572
rect 6880 14600 6886 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 6880 14572 7297 14600
rect 6880 14560 6886 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 7285 14563 7343 14569
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14569 11207 14603
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 11149 14563 11207 14569
rect 1670 14532 1676 14544
rect 1583 14504 1676 14532
rect 1670 14492 1676 14504
rect 1728 14532 1734 14544
rect 2222 14532 2228 14544
rect 1728 14504 2228 14532
rect 1728 14492 1734 14504
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 2590 14541 2596 14544
rect 2587 14532 2596 14541
rect 2551 14504 2596 14532
rect 2587 14495 2596 14504
rect 2590 14492 2596 14495
rect 2648 14492 2654 14544
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4427 14535 4485 14541
rect 4427 14532 4439 14535
rect 4028 14504 4439 14532
rect 4028 14492 4034 14504
rect 4427 14501 4439 14504
rect 4473 14532 4485 14535
rect 6546 14532 6552 14544
rect 4473 14504 6552 14532
rect 4473 14501 4485 14504
rect 4427 14495 4485 14501
rect 6546 14492 6552 14504
rect 6604 14492 6610 14544
rect 7650 14532 7656 14544
rect 7484 14504 7656 14532
rect 5880 14467 5938 14473
rect 5880 14433 5892 14467
rect 5926 14464 5938 14467
rect 5994 14464 6000 14476
rect 5926 14436 6000 14464
rect 5926 14433 5938 14436
rect 5880 14427 5938 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 7484 14473 7512 14504
rect 7650 14492 7656 14504
rect 7708 14532 7714 14544
rect 8754 14532 8760 14544
rect 7708 14504 8760 14532
rect 7708 14492 7714 14504
rect 8754 14492 8760 14504
rect 8812 14492 8818 14544
rect 10591 14535 10649 14541
rect 10591 14501 10603 14535
rect 10637 14532 10649 14535
rect 10778 14532 10784 14544
rect 10637 14504 10784 14532
rect 10637 14501 10649 14504
rect 10591 14495 10649 14501
rect 10778 14492 10784 14504
rect 10836 14492 10842 14544
rect 11164 14532 11192 14563
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 12894 14560 12900 14612
rect 12952 14600 12958 14612
rect 12989 14603 13047 14609
rect 12989 14600 13001 14603
rect 12952 14572 13001 14600
rect 12952 14560 12958 14572
rect 12989 14569 13001 14572
rect 13035 14569 13047 14603
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 12989 14563 13047 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13998 14600 14004 14612
rect 13959 14572 14004 14600
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14090 14560 14096 14612
rect 14148 14600 14154 14612
rect 15013 14603 15071 14609
rect 15013 14600 15025 14603
rect 14148 14572 15025 14600
rect 14148 14560 14154 14572
rect 15013 14569 15025 14572
rect 15059 14569 15071 14603
rect 15013 14563 15071 14569
rect 11422 14532 11428 14544
rect 11164 14504 11428 14532
rect 11422 14492 11428 14504
rect 11480 14532 11486 14544
rect 11480 14504 12756 14532
rect 11480 14492 11486 14504
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14464 8263 14467
rect 8386 14464 8392 14476
rect 8251 14436 8392 14464
rect 8251 14433 8263 14436
rect 8205 14427 8263 14433
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4246 14356 4252 14408
rect 4304 14396 4310 14408
rect 7101 14399 7159 14405
rect 7101 14396 7113 14399
rect 4304 14368 7113 14396
rect 4304 14356 4310 14368
rect 7101 14365 7113 14368
rect 7147 14396 7159 14399
rect 8036 14396 8064 14427
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 10229 14467 10287 14473
rect 10229 14433 10241 14467
rect 10275 14464 10287 14467
rect 12066 14464 12072 14476
rect 10275 14436 12072 14464
rect 10275 14433 10287 14436
rect 10229 14427 10287 14433
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 9858 14396 9864 14408
rect 7147 14368 9864 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12084 14368 12633 14396
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5592 14232 5733 14260
rect 5592 14220 5598 14232
rect 5721 14229 5733 14232
rect 5767 14260 5779 14263
rect 5951 14263 6009 14269
rect 5951 14260 5963 14263
rect 5767 14232 5963 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 5951 14229 5963 14232
rect 5997 14229 6009 14263
rect 5951 14223 6009 14229
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 8754 14260 8760 14272
rect 8711 14232 8760 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9309 14263 9367 14269
rect 9309 14260 9321 14263
rect 9088 14232 9321 14260
rect 9088 14220 9094 14232
rect 9309 14229 9321 14232
rect 9355 14260 9367 14263
rect 9490 14260 9496 14272
rect 9355 14232 9496 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12084 14269 12112 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 12728 14328 12756 14504
rect 12802 14424 12808 14476
rect 12860 14464 12866 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 12860 14436 15301 14464
rect 12860 14424 12866 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15436 14436 15481 14464
rect 15436 14424 15442 14436
rect 14734 14396 14740 14408
rect 14647 14368 14740 14396
rect 14734 14356 14740 14368
rect 14792 14396 14798 14408
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 14792 14368 16865 14396
rect 14792 14356 14798 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 15378 14328 15384 14340
rect 12728 14300 15384 14328
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 11940 14232 12081 14260
rect 11940 14220 11946 14232
rect 12069 14229 12081 14232
rect 12115 14229 12127 14263
rect 12069 14223 12127 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2590 14056 2596 14068
rect 2372 14028 2596 14056
rect 2372 14016 2378 14028
rect 2590 14016 2596 14028
rect 2648 14056 2654 14068
rect 2685 14059 2743 14065
rect 2685 14056 2697 14059
rect 2648 14028 2697 14056
rect 2648 14016 2654 14028
rect 2685 14025 2697 14028
rect 2731 14056 2743 14059
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 2731 14028 3893 14056
rect 2731 14025 2743 14028
rect 2685 14019 2743 14025
rect 3881 14025 3893 14028
rect 3927 14056 3939 14059
rect 3970 14056 3976 14068
rect 3927 14028 3976 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 5445 14059 5503 14065
rect 5445 14025 5457 14059
rect 5491 14056 5503 14059
rect 5994 14056 6000 14068
rect 5491 14028 6000 14056
rect 5491 14025 5503 14028
rect 5445 14019 5503 14025
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6270 14056 6276 14068
rect 6231 14028 6276 14056
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 6420 14028 7757 14056
rect 6420 14016 6426 14028
rect 7745 14025 7757 14028
rect 7791 14056 7803 14059
rect 9030 14056 9036 14068
rect 7791 14028 9036 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 9030 14016 9036 14028
rect 9088 14016 9094 14068
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 13817 14059 13875 14065
rect 13817 14025 13829 14059
rect 13863 14056 13875 14059
rect 13998 14056 14004 14068
rect 13863 14028 14004 14056
rect 13863 14025 13875 14028
rect 13817 14019 13875 14025
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 14826 14056 14832 14068
rect 14608 14028 14832 14056
rect 14608 14016 14614 14028
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15378 14016 15384 14068
rect 15436 14056 15442 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 15436 14028 15669 14056
rect 15436 14016 15442 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 6546 13988 6552 14000
rect 6507 13960 6552 13988
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 8846 13988 8852 14000
rect 8807 13960 8852 13988
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 10321 13991 10379 13997
rect 10321 13957 10333 13991
rect 10367 13988 10379 13991
rect 10778 13988 10784 14000
rect 10367 13960 10784 13988
rect 10367 13957 10379 13960
rect 10321 13951 10379 13957
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 12250 13948 12256 14000
rect 12308 13988 12314 14000
rect 16025 13991 16083 13997
rect 16025 13988 16037 13991
rect 12308 13960 16037 13988
rect 12308 13948 12314 13960
rect 16025 13957 16037 13960
rect 16071 13957 16083 13991
rect 16025 13951 16083 13957
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 3559 13892 3924 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2682 13852 2688 13864
rect 2363 13824 2688 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2682 13812 2688 13824
rect 2740 13852 2746 13864
rect 3418 13852 3424 13864
rect 2740 13824 3424 13852
rect 2740 13812 2746 13824
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3896 13852 3924 13892
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 6822 13920 6828 13932
rect 4120 13892 4752 13920
rect 6783 13892 6828 13920
rect 4120 13880 4126 13892
rect 4246 13852 4252 13864
rect 3896 13824 4252 13852
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4522 13852 4528 13864
rect 4479 13824 4528 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 1765 13787 1823 13793
rect 1765 13784 1777 13787
rect 1728 13756 1777 13784
rect 1728 13744 1734 13756
rect 1765 13753 1777 13756
rect 1811 13784 1823 13787
rect 1854 13784 1860 13796
rect 1811 13756 1860 13784
rect 1811 13753 1823 13756
rect 1765 13747 1823 13753
rect 1854 13744 1860 13756
rect 1912 13744 1918 13796
rect 3145 13787 3203 13793
rect 3145 13753 3157 13787
rect 3191 13784 3203 13787
rect 4448 13784 4476 13815
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 4724 13861 4752 13892
rect 6822 13880 6828 13892
rect 6880 13880 6886 13932
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 8720 13923 8778 13929
rect 8720 13920 8732 13923
rect 8628 13892 8732 13920
rect 8628 13880 8634 13892
rect 8720 13889 8732 13892
rect 8766 13889 8778 13923
rect 8720 13883 8778 13889
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 4709 13855 4767 13861
rect 4709 13821 4721 13855
rect 4755 13852 4767 13855
rect 4985 13855 5043 13861
rect 4985 13852 4997 13855
rect 4755 13824 4997 13852
rect 4755 13821 4767 13824
rect 4709 13815 4767 13821
rect 4985 13821 4997 13824
rect 5031 13821 5043 13855
rect 5534 13852 5540 13864
rect 5495 13824 5540 13852
rect 4985 13815 5043 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8956 13852 8984 13883
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 9916 13892 10701 13920
rect 9916 13880 9922 13892
rect 10689 13889 10701 13892
rect 10735 13920 10747 13923
rect 14090 13920 14096 13932
rect 10735 13892 14096 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 11072 13861 11100 13892
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14734 13920 14740 13932
rect 14695 13892 14740 13920
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 14826 13880 14832 13932
rect 14884 13920 14890 13932
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14884 13892 15025 13920
rect 14884 13880 14890 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 8343 13824 8984 13852
rect 11057 13855 11115 13861
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 11057 13821 11069 13855
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 11241 13855 11299 13861
rect 11241 13821 11253 13855
rect 11287 13821 11299 13855
rect 11241 13815 11299 13821
rect 11517 13855 11575 13861
rect 11517 13821 11529 13855
rect 11563 13852 11575 13855
rect 11974 13852 11980 13864
rect 11563 13824 11980 13852
rect 11563 13821 11575 13824
rect 11517 13815 11575 13821
rect 3191 13756 4476 13784
rect 3191 13753 3203 13756
rect 3145 13747 3203 13753
rect 6546 13744 6552 13796
rect 6604 13784 6610 13796
rect 7146 13787 7204 13793
rect 7146 13784 7158 13787
rect 6604 13756 7158 13784
rect 6604 13744 6610 13756
rect 7146 13753 7158 13756
rect 7192 13784 7204 13787
rect 7374 13784 7380 13796
rect 7192 13756 7380 13784
rect 7192 13753 7204 13756
rect 7146 13747 7204 13753
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 8113 13787 8171 13793
rect 8113 13753 8125 13787
rect 8159 13784 8171 13787
rect 8573 13787 8631 13793
rect 8573 13784 8585 13787
rect 8159 13756 8585 13784
rect 8159 13753 8171 13756
rect 8113 13747 8171 13753
rect 8573 13753 8585 13756
rect 8619 13784 8631 13787
rect 8754 13784 8760 13796
rect 8619 13756 8760 13784
rect 8619 13753 8631 13756
rect 8573 13747 8631 13753
rect 8754 13744 8760 13756
rect 8812 13744 8818 13796
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 5721 13719 5779 13725
rect 5721 13716 5733 13719
rect 3936 13688 5733 13716
rect 3936 13676 3942 13688
rect 5721 13685 5733 13688
rect 5767 13685 5779 13719
rect 5721 13679 5779 13685
rect 8297 13719 8355 13725
rect 8297 13685 8309 13719
rect 8343 13716 8355 13719
rect 8386 13716 8392 13728
rect 8343 13688 8392 13716
rect 8343 13685 8355 13688
rect 8297 13679 8355 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 9858 13716 9864 13728
rect 9819 13688 9864 13716
rect 9858 13676 9864 13688
rect 9916 13716 9922 13728
rect 11256 13716 11284 13815
rect 11974 13812 11980 13824
rect 12032 13852 12038 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12032 13824 12909 13852
rect 12032 13812 12038 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 16040 13852 16068 13951
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 16040 13824 16313 13852
rect 12897 13815 12955 13821
rect 16301 13821 16313 13824
rect 16347 13821 16359 13855
rect 18230 13852 18236 13864
rect 18143 13824 18236 13852
rect 16301 13815 16359 13821
rect 18230 13812 18236 13824
rect 18288 13852 18294 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18288 13824 18797 13852
rect 18288 13812 18294 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 11698 13744 11704 13796
rect 11756 13784 11762 13796
rect 12161 13787 12219 13793
rect 12161 13784 12173 13787
rect 11756 13756 12173 13784
rect 11756 13744 11762 13756
rect 12161 13753 12173 13756
rect 12207 13784 12219 13787
rect 12713 13787 12771 13793
rect 12713 13784 12725 13787
rect 12207 13756 12725 13784
rect 12207 13753 12219 13756
rect 12161 13747 12219 13753
rect 12713 13753 12725 13756
rect 12759 13784 12771 13787
rect 13218 13787 13276 13793
rect 13218 13784 13230 13787
rect 12759 13756 13230 13784
rect 12759 13753 12771 13756
rect 12713 13747 12771 13753
rect 12912 13728 12940 13756
rect 13218 13753 13230 13756
rect 13264 13753 13276 13787
rect 13218 13747 13276 13753
rect 14553 13787 14611 13793
rect 14553 13753 14565 13787
rect 14599 13784 14611 13787
rect 14826 13784 14832 13796
rect 14599 13756 14832 13784
rect 14599 13753 14611 13756
rect 14553 13747 14611 13753
rect 14826 13744 14832 13756
rect 14884 13744 14890 13796
rect 16206 13784 16212 13796
rect 16167 13756 16212 13784
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 11790 13716 11796 13728
rect 9916 13688 11796 13716
rect 9916 13676 9922 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 11885 13719 11943 13725
rect 11885 13685 11897 13719
rect 11931 13716 11943 13719
rect 12066 13716 12072 13728
rect 11931 13688 12072 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 12066 13676 12072 13688
rect 12124 13676 12130 13728
rect 12894 13676 12900 13728
rect 12952 13676 12958 13728
rect 14185 13719 14243 13725
rect 14185 13685 14197 13719
rect 14231 13716 14243 13719
rect 14366 13716 14372 13728
rect 14231 13688 14372 13716
rect 14231 13685 14243 13688
rect 14185 13679 14243 13685
rect 14366 13676 14372 13688
rect 14424 13676 14430 13728
rect 18414 13716 18420 13728
rect 18375 13688 18420 13716
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1670 13512 1676 13524
rect 1631 13484 1676 13512
rect 1670 13472 1676 13484
rect 1728 13472 1734 13524
rect 2222 13472 2228 13524
rect 2280 13512 2286 13524
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 2280 13484 3249 13512
rect 2280 13472 2286 13484
rect 3237 13481 3249 13484
rect 3283 13512 3295 13515
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 3283 13484 4169 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4580 13484 4844 13512
rect 4580 13472 4586 13484
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 1946 13444 1952 13456
rect 1544 13416 1952 13444
rect 1544 13404 1550 13416
rect 1946 13404 1952 13416
rect 2004 13444 2010 13456
rect 2041 13447 2099 13453
rect 2041 13444 2053 13447
rect 2004 13416 2053 13444
rect 2004 13404 2010 13416
rect 2041 13413 2053 13416
rect 2087 13413 2099 13447
rect 2041 13407 2099 13413
rect 2593 13447 2651 13453
rect 2593 13413 2605 13447
rect 2639 13444 2651 13447
rect 2682 13444 2688 13456
rect 2639 13416 2688 13444
rect 2639 13413 2651 13416
rect 2593 13407 2651 13413
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 4212 13348 4257 13376
rect 4212 13336 4218 13348
rect 4522 13336 4528 13388
rect 4580 13376 4586 13388
rect 4580 13348 4625 13376
rect 4580 13336 4586 13348
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2130 13308 2136 13320
rect 1995 13280 2136 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2130 13268 2136 13280
rect 2188 13308 2194 13320
rect 3605 13311 3663 13317
rect 3605 13308 3617 13311
rect 2188 13280 3617 13308
rect 2188 13268 2194 13280
rect 3605 13277 3617 13280
rect 3651 13277 3663 13311
rect 4816 13308 4844 13484
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 10778 13512 10784 13524
rect 7432 13484 10784 13512
rect 7432 13472 7438 13484
rect 6086 13404 6092 13456
rect 6144 13444 6150 13456
rect 6730 13444 6736 13456
rect 6144 13416 6736 13444
rect 6144 13404 6150 13416
rect 6730 13404 6736 13416
rect 6788 13444 6794 13456
rect 10698 13453 10726 13484
rect 10778 13472 10784 13484
rect 10836 13512 10842 13524
rect 11698 13512 11704 13524
rect 10836 13484 11704 13512
rect 10836 13472 10842 13484
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 11974 13512 11980 13524
rect 11935 13484 11980 13512
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 15381 13515 15439 13521
rect 15381 13512 15393 13515
rect 12124 13484 15393 13512
rect 12124 13472 12130 13484
rect 15381 13481 15393 13484
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 16991 13515 17049 13521
rect 16991 13481 17003 13515
rect 17037 13512 17049 13515
rect 18230 13512 18236 13524
rect 17037 13484 18236 13512
rect 17037 13481 17049 13484
rect 16991 13475 17049 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 10683 13447 10741 13453
rect 10683 13444 10695 13447
rect 6788 13416 9674 13444
rect 10661 13416 10695 13444
rect 6788 13404 6794 13416
rect 9646 13388 9674 13416
rect 10683 13413 10695 13416
rect 10729 13413 10741 13447
rect 12250 13444 12256 13456
rect 10683 13407 10741 13413
rect 11256 13416 12256 13444
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 6270 13376 6276 13388
rect 5675 13348 6276 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 7101 13379 7159 13385
rect 7101 13376 7113 13379
rect 6696 13348 7113 13376
rect 6696 13336 6702 13348
rect 7101 13345 7113 13348
rect 7147 13345 7159 13379
rect 7101 13339 7159 13345
rect 7202 13348 7604 13376
rect 9646 13348 9680 13388
rect 7202 13308 7230 13348
rect 4816 13280 7230 13308
rect 3605 13271 3663 13277
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7576 13317 7604 13348
rect 9674 13336 9680 13348
rect 9732 13376 9738 13388
rect 11256 13385 11284 13416
rect 12250 13404 12256 13416
rect 12308 13444 12314 13456
rect 12618 13444 12624 13456
rect 12308 13416 12624 13444
rect 12308 13404 12314 13416
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 12802 13444 12808 13456
rect 12763 13416 12808 13444
rect 12802 13404 12808 13416
rect 12860 13404 12866 13456
rect 12986 13404 12992 13456
rect 13044 13444 13050 13456
rect 13081 13447 13139 13453
rect 13081 13444 13093 13447
rect 13044 13416 13093 13444
rect 13044 13404 13050 13416
rect 13081 13413 13093 13416
rect 13127 13444 13139 13447
rect 14369 13447 14427 13453
rect 13127 13416 13814 13444
rect 13127 13413 13139 13416
rect 13081 13407 13139 13413
rect 11241 13379 11299 13385
rect 9732 13348 9996 13376
rect 9732 13336 9738 13348
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7432 13280 7481 13308
rect 7432 13268 7438 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 2961 13243 3019 13249
rect 2961 13240 2973 13243
rect 2464 13212 2973 13240
rect 2464 13200 2470 13212
rect 2961 13209 2973 13212
rect 3007 13240 3019 13243
rect 4982 13240 4988 13252
rect 3007 13212 4988 13240
rect 3007 13209 3019 13212
rect 2961 13203 3019 13209
rect 4982 13200 4988 13212
rect 5040 13200 5046 13252
rect 7266 13243 7324 13249
rect 7266 13209 7278 13243
rect 7312 13240 7324 13243
rect 8018 13240 8024 13252
rect 7312 13212 8024 13240
rect 7312 13209 7324 13212
rect 7266 13203 7324 13209
rect 8018 13200 8024 13212
rect 8076 13200 8082 13252
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 8665 13243 8723 13249
rect 8665 13240 8677 13243
rect 8628 13212 8677 13240
rect 8628 13200 8634 13212
rect 8665 13209 8677 13212
rect 8711 13240 8723 13243
rect 9122 13240 9128 13252
rect 8711 13212 9128 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 9122 13200 9128 13212
rect 9180 13240 9186 13252
rect 9766 13240 9772 13252
rect 9180 13212 9772 13240
rect 9180 13200 9186 13212
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 9968 13249 9996 13348
rect 11241 13345 11253 13379
rect 11287 13345 11299 13379
rect 11241 13339 11299 13345
rect 11425 13379 11483 13385
rect 11425 13345 11437 13379
rect 11471 13376 11483 13379
rect 11471 13348 12020 13376
rect 11471 13345 11483 13348
rect 11425 13339 11483 13345
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10778 13308 10784 13320
rect 10367 13280 10784 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11992 13308 12020 13348
rect 13170 13336 13176 13388
rect 13228 13376 13234 13388
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13228 13348 13645 13376
rect 13228 13336 13234 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 11348 13280 11652 13308
rect 11992 13280 12173 13308
rect 9953 13243 10011 13249
rect 9953 13209 9965 13243
rect 9999 13240 10011 13243
rect 11348 13240 11376 13280
rect 9999 13212 11376 13240
rect 9999 13209 10011 13212
rect 9953 13203 10011 13209
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 3752 13144 5825 13172
rect 3752 13132 3758 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 6270 13172 6276 13184
rect 6231 13144 6276 13172
rect 5813 13135 5871 13141
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 7006 13172 7012 13184
rect 6967 13144 7012 13172
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7377 13175 7435 13181
rect 7377 13141 7389 13175
rect 7423 13172 7435 13175
rect 7742 13172 7748 13184
rect 7423 13144 7748 13172
rect 7423 13141 7435 13144
rect 7377 13135 7435 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 8205 13175 8263 13181
rect 8205 13141 8217 13175
rect 8251 13172 8263 13175
rect 8294 13172 8300 13184
rect 8251 13144 8300 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8294 13132 8300 13144
rect 8352 13132 8358 13184
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 9030 13172 9036 13184
rect 8904 13144 9036 13172
rect 8904 13132 8910 13144
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 11112 13144 11437 13172
rect 11112 13132 11118 13144
rect 11425 13141 11437 13144
rect 11471 13172 11483 13175
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11471 13144 11529 13172
rect 11471 13141 11483 13144
rect 11425 13135 11483 13141
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11624 13172 11652 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 13786 13308 13814 13416
rect 14369 13413 14381 13447
rect 14415 13444 14427 13447
rect 14415 13416 15792 13444
rect 14415 13413 14427 13416
rect 14369 13407 14427 13413
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 14642 13376 14648 13388
rect 14332 13348 14648 13376
rect 14332 13336 14338 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 14826 13336 14832 13388
rect 14884 13376 14890 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 14884 13348 15301 13376
rect 14884 13336 14890 13348
rect 15289 13345 15301 13348
rect 15335 13376 15347 13379
rect 15562 13376 15568 13388
rect 15335 13348 15568 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 15764 13385 15792 13416
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 16022 13376 16028 13388
rect 15795 13348 16028 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16920 13379 16978 13385
rect 16920 13345 16932 13379
rect 16966 13376 16978 13379
rect 17310 13376 17316 13388
rect 16966 13348 17316 13376
rect 16966 13345 16978 13348
rect 16920 13339 16978 13345
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 24581 13379 24639 13385
rect 24581 13345 24593 13379
rect 24627 13376 24639 13379
rect 24670 13376 24676 13388
rect 24627 13348 24676 13376
rect 24627 13345 24639 13348
rect 24581 13339 24639 13345
rect 24670 13336 24676 13348
rect 24728 13336 24734 13388
rect 14001 13311 14059 13317
rect 14001 13308 14013 13311
rect 13786 13280 14013 13308
rect 12161 13271 12219 13277
rect 14001 13277 14013 13280
rect 14047 13308 14059 13311
rect 14366 13308 14372 13320
rect 14047 13280 14372 13308
rect 14047 13277 14059 13280
rect 14001 13271 14059 13277
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 13538 13200 13544 13252
rect 13596 13240 13602 13252
rect 13798 13243 13856 13249
rect 13798 13240 13810 13243
rect 13596 13212 13810 13240
rect 13596 13200 13602 13212
rect 13798 13209 13810 13212
rect 13844 13240 13856 13243
rect 14182 13240 14188 13252
rect 13844 13212 14188 13240
rect 13844 13209 13856 13212
rect 13798 13203 13856 13209
rect 14182 13200 14188 13212
rect 14240 13240 14246 13252
rect 14645 13243 14703 13249
rect 14645 13240 14657 13243
rect 14240 13212 14657 13240
rect 14240 13200 14246 13212
rect 14645 13209 14657 13212
rect 14691 13209 14703 13243
rect 14645 13203 14703 13209
rect 13446 13172 13452 13184
rect 11624 13144 13452 13172
rect 11517 13135 11575 13141
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 13906 13172 13912 13184
rect 13867 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 24719 13175 24777 13181
rect 24719 13172 24731 13175
rect 15436 13144 24731 13172
rect 15436 13132 15442 13144
rect 24719 13141 24731 13144
rect 24765 13141 24777 13175
rect 24719 13135 24777 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 1857 12971 1915 12977
rect 1857 12968 1869 12971
rect 1820 12940 1869 12968
rect 1820 12928 1826 12940
rect 1857 12937 1869 12940
rect 1903 12937 1915 12971
rect 1857 12931 1915 12937
rect 1946 12928 1952 12980
rect 2004 12968 2010 12980
rect 3329 12971 3387 12977
rect 3329 12968 3341 12971
rect 2004 12940 3341 12968
rect 2004 12928 2010 12940
rect 3329 12937 3341 12940
rect 3375 12937 3387 12971
rect 3329 12931 3387 12937
rect 4065 12971 4123 12977
rect 4065 12937 4077 12971
rect 4111 12968 4123 12971
rect 4522 12968 4528 12980
rect 4111 12940 4528 12968
rect 4111 12937 4123 12940
rect 4065 12931 4123 12937
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 6420 12940 7205 12968
rect 6420 12928 6426 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 8110 12968 8116 12980
rect 7193 12931 7251 12937
rect 7392 12940 8116 12968
rect 7392 12912 7420 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8662 12968 8668 12980
rect 8623 12940 8668 12968
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 9950 12968 9956 12980
rect 8812 12940 9956 12968
rect 8812 12928 8818 12940
rect 9950 12928 9956 12940
rect 10008 12968 10014 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 10008 12940 11345 12968
rect 10008 12928 10014 12940
rect 11333 12937 11345 12940
rect 11379 12968 11391 12971
rect 13170 12968 13176 12980
rect 11379 12940 13176 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 14182 12977 14188 12980
rect 14166 12971 14188 12977
rect 14166 12937 14178 12971
rect 14166 12931 14188 12937
rect 14182 12928 14188 12931
rect 14240 12928 14246 12980
rect 14458 12968 14464 12980
rect 14419 12940 14464 12968
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 2314 12900 2320 12912
rect 2275 12872 2320 12900
rect 2314 12860 2320 12872
rect 2372 12860 2378 12912
rect 3697 12903 3755 12909
rect 3697 12869 3709 12903
rect 3743 12900 3755 12903
rect 4154 12900 4160 12912
rect 3743 12872 4160 12900
rect 3743 12869 3755 12872
rect 3697 12863 3755 12869
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 6273 12903 6331 12909
rect 6273 12869 6285 12903
rect 6319 12900 6331 12903
rect 7374 12900 7380 12912
rect 6319 12872 7380 12900
rect 6319 12869 6331 12872
rect 6273 12863 6331 12869
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 7466 12860 7472 12912
rect 7524 12900 7530 12912
rect 8294 12900 8300 12912
rect 7524 12872 8300 12900
rect 7524 12860 7530 12872
rect 8294 12860 8300 12872
rect 8352 12900 8358 12912
rect 9582 12900 9588 12912
rect 8352 12872 9588 12900
rect 8352 12860 8358 12872
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 9766 12909 9772 12912
rect 9750 12903 9772 12909
rect 9750 12869 9762 12903
rect 9750 12863 9772 12869
rect 9766 12860 9772 12863
rect 9824 12860 9830 12912
rect 9861 12903 9919 12909
rect 9861 12869 9873 12903
rect 9907 12900 9919 12903
rect 10965 12903 11023 12909
rect 10965 12900 10977 12903
rect 9907 12872 10977 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 10965 12869 10977 12872
rect 11011 12869 11023 12903
rect 10965 12863 11023 12869
rect 1535 12835 1593 12841
rect 1535 12801 1547 12835
rect 1581 12832 1593 12835
rect 2866 12832 2872 12844
rect 1581 12804 2872 12832
rect 1581 12801 1593 12804
rect 1535 12795 1593 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4479 12804 5488 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 5460 12776 5488 12804
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8168 12835 8226 12841
rect 8168 12832 8180 12835
rect 8076 12804 8180 12832
rect 8076 12792 8082 12804
rect 8168 12801 8180 12804
rect 8214 12801 8226 12835
rect 8386 12832 8392 12844
rect 8347 12804 8392 12832
rect 8168 12795 8226 12801
rect 8386 12792 8392 12804
rect 8444 12792 8450 12844
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 9030 12832 9036 12844
rect 8628 12804 9036 12832
rect 8628 12792 8634 12804
rect 9030 12792 9036 12804
rect 9088 12832 9094 12844
rect 9876 12832 9904 12863
rect 12802 12860 12808 12912
rect 12860 12900 12866 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12860 12872 13093 12900
rect 12860 12860 12866 12872
rect 13081 12869 13093 12872
rect 13127 12869 13139 12903
rect 13081 12863 13139 12869
rect 13725 12903 13783 12909
rect 13725 12869 13737 12903
rect 13771 12900 13783 12903
rect 13906 12900 13912 12912
rect 13771 12872 13912 12900
rect 13771 12869 13783 12872
rect 13725 12863 13783 12869
rect 13906 12860 13912 12872
rect 13964 12900 13970 12912
rect 14274 12900 14280 12912
rect 13964 12872 14280 12900
rect 13964 12860 13970 12872
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 15289 12903 15347 12909
rect 15289 12900 15301 12903
rect 14884 12872 15301 12900
rect 14884 12860 14890 12872
rect 15289 12869 15301 12872
rect 15335 12869 15347 12903
rect 15289 12863 15347 12869
rect 9088 12804 9904 12832
rect 9953 12835 10011 12841
rect 9088 12792 9094 12804
rect 9953 12801 9965 12835
rect 9999 12832 10011 12835
rect 10042 12832 10048 12844
rect 9999 12804 10048 12832
rect 9999 12801 10011 12804
rect 9953 12795 10011 12801
rect 10042 12792 10048 12804
rect 10100 12792 10106 12844
rect 10686 12832 10692 12844
rect 10647 12804 10692 12832
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 14366 12832 14372 12844
rect 12575 12804 14209 12832
rect 14327 12804 14372 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 1448 12767 1506 12773
rect 1448 12733 1460 12767
rect 1494 12764 1506 12767
rect 1762 12764 1768 12776
rect 1494 12736 1768 12764
rect 1494 12733 1506 12736
rect 1448 12727 1506 12733
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2406 12764 2412 12776
rect 2367 12736 2412 12764
rect 2406 12724 2412 12736
rect 2464 12724 2470 12776
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5166 12764 5172 12776
rect 4847 12736 5172 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5442 12724 5448 12776
rect 5500 12764 5506 12776
rect 7006 12764 7012 12776
rect 5500 12736 5593 12764
rect 6919 12736 7012 12764
rect 5500 12724 5506 12736
rect 7006 12724 7012 12736
rect 7064 12764 7070 12776
rect 8294 12764 8300 12776
rect 7064 12736 8300 12764
rect 7064 12724 7070 12736
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 8680 12736 11161 12764
rect 8680 12708 8708 12736
rect 11149 12733 11161 12736
rect 11195 12764 11207 12767
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11195 12736 11621 12764
rect 11195 12733 11207 12736
rect 11149 12727 11207 12733
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 13446 12724 13452 12776
rect 13504 12764 13510 12776
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13504 12736 14013 12764
rect 13504 12724 13510 12736
rect 14001 12733 14013 12736
rect 14047 12733 14059 12767
rect 14181 12764 14209 12804
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 14458 12792 14464 12844
rect 14516 12832 14522 12844
rect 16577 12835 16635 12841
rect 16577 12832 16589 12835
rect 14516 12804 16589 12832
rect 14516 12792 14522 12804
rect 15378 12764 15384 12776
rect 14181 12736 15384 12764
rect 14001 12727 14059 12733
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 15470 12724 15476 12776
rect 15528 12764 15534 12776
rect 15580 12773 15608 12804
rect 16577 12801 16589 12804
rect 16623 12801 16635 12835
rect 16577 12795 16635 12801
rect 15565 12767 15623 12773
rect 15565 12764 15577 12767
rect 15528 12736 15577 12764
rect 15528 12724 15534 12736
rect 15565 12733 15577 12736
rect 15611 12733 15623 12767
rect 16022 12764 16028 12776
rect 15983 12736 16028 12764
rect 15565 12727 15623 12733
rect 16022 12724 16028 12736
rect 16080 12764 16086 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16080 12736 16957 12764
rect 16080 12724 16086 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 2314 12656 2320 12708
rect 2372 12696 2378 12708
rect 2682 12696 2688 12708
rect 2372 12668 2688 12696
rect 2372 12656 2378 12668
rect 2682 12656 2688 12668
rect 2740 12705 2746 12708
rect 2740 12699 2788 12705
rect 2740 12665 2742 12699
rect 2776 12665 2788 12699
rect 2740 12659 2788 12665
rect 7469 12699 7527 12705
rect 7469 12665 7481 12699
rect 7515 12696 7527 12699
rect 7742 12696 7748 12708
rect 7515 12668 7748 12696
rect 7515 12665 7527 12668
rect 7469 12659 7527 12665
rect 2740 12656 2746 12659
rect 7742 12656 7748 12668
rect 7800 12656 7806 12708
rect 8021 12699 8079 12705
rect 8021 12665 8033 12699
rect 8067 12696 8079 12699
rect 8662 12696 8668 12708
rect 8067 12668 8668 12696
rect 8067 12665 8079 12668
rect 8021 12659 8079 12665
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 9585 12699 9643 12705
rect 8772 12668 9536 12696
rect 4982 12628 4988 12640
rect 4943 12600 4988 12628
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 7558 12588 7564 12640
rect 7616 12628 7622 12640
rect 7929 12631 7987 12637
rect 7929 12628 7941 12631
rect 7616 12600 7941 12628
rect 7616 12588 7622 12600
rect 7929 12597 7941 12600
rect 7975 12628 7987 12631
rect 8386 12628 8392 12640
rect 7975 12600 8392 12628
rect 7975 12597 7987 12600
rect 7929 12591 7987 12597
rect 8386 12588 8392 12600
rect 8444 12628 8450 12640
rect 8772 12628 8800 12668
rect 9122 12628 9128 12640
rect 8444 12600 8800 12628
rect 9083 12600 9128 12628
rect 8444 12588 8450 12600
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9508 12637 9536 12668
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 9674 12696 9680 12708
rect 9631 12668 9680 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10321 12699 10379 12705
rect 10321 12665 10333 12699
rect 10367 12696 10379 12699
rect 10870 12696 10876 12708
rect 10367 12668 10876 12696
rect 10367 12665 10379 12668
rect 10321 12659 10379 12665
rect 10870 12656 10876 12668
rect 10928 12656 10934 12708
rect 12253 12699 12311 12705
rect 12253 12665 12265 12699
rect 12299 12696 12311 12699
rect 12621 12699 12679 12705
rect 12621 12696 12633 12699
rect 12299 12668 12633 12696
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 12621 12665 12633 12668
rect 12667 12696 12679 12699
rect 16206 12696 16212 12708
rect 12667 12668 16212 12696
rect 12667 12665 12679 12668
rect 12621 12659 12679 12665
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 9493 12631 9551 12637
rect 9493 12597 9505 12631
rect 9539 12628 9551 12631
rect 9766 12628 9772 12640
rect 9539 12600 9772 12628
rect 9539 12597 9551 12600
rect 9493 12591 9551 12597
rect 9766 12588 9772 12600
rect 9824 12628 9830 12640
rect 10042 12628 10048 12640
rect 9824 12600 10048 12628
rect 9824 12588 9830 12600
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 15654 12628 15660 12640
rect 15615 12600 15660 12628
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 17310 12628 17316 12640
rect 17271 12600 17316 12628
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1673 12427 1731 12433
rect 1673 12424 1685 12427
rect 1636 12396 1685 12424
rect 1636 12384 1642 12396
rect 1673 12393 1685 12396
rect 1719 12424 1731 12427
rect 2038 12424 2044 12436
rect 1719 12396 2044 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 2038 12384 2044 12396
rect 2096 12384 2102 12436
rect 2774 12424 2780 12436
rect 2424 12396 2780 12424
rect 2424 12368 2452 12396
rect 2774 12384 2780 12396
rect 2832 12384 2838 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 6273 12427 6331 12433
rect 6273 12424 6285 12427
rect 5500 12396 6285 12424
rect 5500 12384 5506 12396
rect 6273 12393 6285 12396
rect 6319 12424 6331 12427
rect 6362 12424 6368 12436
rect 6319 12396 6368 12424
rect 6319 12393 6331 12396
rect 6273 12387 6331 12393
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 7834 12424 7840 12436
rect 7795 12396 7840 12424
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 10870 12424 10876 12436
rect 10831 12396 10876 12424
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 15654 12424 15660 12436
rect 12728 12396 15660 12424
rect 1946 12356 1952 12368
rect 1907 12328 1952 12356
rect 1946 12316 1952 12328
rect 2004 12316 2010 12368
rect 2406 12356 2412 12368
rect 2319 12328 2412 12356
rect 2406 12316 2412 12328
rect 2464 12316 2470 12368
rect 2501 12359 2559 12365
rect 2501 12325 2513 12359
rect 2547 12356 2559 12359
rect 2866 12356 2872 12368
rect 2547 12328 2872 12356
rect 2547 12325 2559 12328
rect 2501 12319 2559 12325
rect 2866 12316 2872 12328
rect 2924 12316 2930 12368
rect 5258 12316 5264 12368
rect 5316 12356 5322 12368
rect 8846 12356 8852 12368
rect 5316 12328 8852 12356
rect 5316 12316 5322 12328
rect 8846 12316 8852 12328
rect 8904 12316 8910 12368
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 8996 12328 10358 12356
rect 8996 12316 9002 12328
rect 4062 12288 4068 12300
rect 4023 12260 4068 12288
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4338 12248 4344 12300
rect 4396 12288 4402 12300
rect 4525 12291 4583 12297
rect 4525 12288 4537 12291
rect 4396 12260 4537 12288
rect 4396 12248 4402 12260
rect 4525 12257 4537 12260
rect 4571 12288 4583 12291
rect 5166 12288 5172 12300
rect 4571 12260 5172 12288
rect 4571 12257 4583 12260
rect 4525 12251 4583 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 5592 12260 5641 12288
rect 5592 12248 5598 12260
rect 5629 12257 5641 12260
rect 5675 12288 5687 12291
rect 6086 12288 6092 12300
rect 5675 12260 6092 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 6086 12248 6092 12260
rect 6144 12248 6150 12300
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 6696 12260 7205 12288
rect 6696 12248 6702 12260
rect 7193 12257 7205 12260
rect 7239 12288 7251 12291
rect 8202 12288 8208 12300
rect 7239 12260 8208 12288
rect 7239 12257 7251 12260
rect 7193 12251 7251 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 9950 12288 9956 12300
rect 9723 12260 9956 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10330 12288 10358 12328
rect 10778 12316 10784 12368
rect 10836 12356 10842 12368
rect 11241 12359 11299 12365
rect 11241 12356 11253 12359
rect 10836 12328 11253 12356
rect 10836 12316 10842 12328
rect 11241 12325 11253 12328
rect 11287 12356 11299 12359
rect 12728 12356 12756 12396
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 16080 12396 16313 12424
rect 16080 12384 16086 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 13170 12356 13176 12368
rect 11287 12328 12756 12356
rect 13131 12328 13176 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 13538 12356 13544 12368
rect 13499 12328 13544 12356
rect 13538 12316 13544 12328
rect 13596 12316 13602 12368
rect 13817 12359 13875 12365
rect 13817 12325 13829 12359
rect 13863 12356 13875 12359
rect 14366 12356 14372 12368
rect 13863 12328 14372 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 15105 12359 15163 12365
rect 15105 12325 15117 12359
rect 15151 12356 15163 12359
rect 15378 12356 15384 12368
rect 15151 12328 15384 12356
rect 15151 12325 15163 12328
rect 15105 12319 15163 12325
rect 15378 12316 15384 12328
rect 15436 12316 15442 12368
rect 15473 12359 15531 12365
rect 15473 12325 15485 12359
rect 15519 12356 15531 12359
rect 15562 12356 15568 12368
rect 15519 12328 15568 12356
rect 15519 12325 15531 12328
rect 15473 12319 15531 12325
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 11609 12291 11667 12297
rect 11609 12288 11621 12291
rect 10330 12260 11621 12288
rect 11609 12257 11621 12260
rect 11655 12288 11667 12291
rect 11698 12288 11704 12300
rect 11655 12260 11704 12288
rect 11655 12257 11667 12260
rect 11609 12251 11667 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11848 12260 12081 12288
rect 11848 12248 11854 12260
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12288 17923 12291
rect 18230 12288 18236 12300
rect 17911 12260 18236 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 18230 12248 18236 12260
rect 18288 12248 18294 12300
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 2556 12192 2697 12220
rect 2556 12180 2562 12192
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 4614 12220 4620 12232
rect 4575 12192 4620 12220
rect 2685 12183 2743 12189
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5994 12220 6000 12232
rect 5907 12192 6000 12220
rect 5994 12180 6000 12192
rect 6052 12220 6058 12232
rect 7558 12220 7564 12232
rect 6052 12192 7564 12220
rect 6052 12180 6058 12192
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9824 12192 10057 12220
rect 9824 12180 9830 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 13722 12220 13728 12232
rect 13683 12192 13728 12220
rect 10045 12183 10103 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 13998 12220 14004 12232
rect 13959 12192 14004 12220
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 14734 12180 14740 12232
rect 14792 12220 14798 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 14792 12192 15393 12220
rect 14792 12180 14798 12192
rect 15381 12189 15393 12192
rect 15427 12220 15439 12223
rect 16853 12223 16911 12229
rect 16853 12220 16865 12223
rect 15427 12192 16865 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 16853 12189 16865 12192
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 5794 12155 5852 12161
rect 5794 12121 5806 12155
rect 5840 12152 5852 12155
rect 6546 12152 6552 12164
rect 5840 12124 6552 12152
rect 5840 12121 5852 12124
rect 5794 12115 5852 12121
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 9953 12155 10011 12161
rect 9953 12152 9965 12155
rect 9640 12124 9965 12152
rect 9640 12112 9646 12124
rect 9953 12121 9965 12124
rect 9999 12152 10011 12155
rect 14274 12152 14280 12164
rect 9999 12124 14280 12152
rect 9999 12121 10011 12124
rect 9953 12115 10011 12121
rect 14274 12112 14280 12124
rect 14332 12152 14338 12164
rect 14645 12155 14703 12161
rect 14645 12152 14657 12155
rect 14332 12124 14657 12152
rect 14332 12112 14338 12124
rect 14645 12121 14657 12124
rect 14691 12152 14703 12155
rect 14691 12124 15332 12152
rect 14691 12121 14703 12124
rect 14645 12115 14703 12121
rect 3418 12084 3424 12096
rect 3331 12056 3424 12084
rect 3418 12044 3424 12056
rect 3476 12084 3482 12096
rect 4798 12084 4804 12096
rect 3476 12056 4804 12084
rect 3476 12044 3482 12056
rect 4798 12044 4804 12056
rect 4856 12044 4862 12096
rect 5166 12084 5172 12096
rect 5127 12056 5172 12084
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 5905 12087 5963 12093
rect 5905 12053 5917 12087
rect 5951 12084 5963 12087
rect 6178 12084 6184 12096
rect 5951 12056 6184 12084
rect 5951 12053 5963 12056
rect 5905 12047 5963 12053
rect 6178 12044 6184 12056
rect 6236 12044 6242 12096
rect 6638 12084 6644 12096
rect 6599 12056 6644 12084
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 7006 12084 7012 12096
rect 6967 12056 7012 12084
rect 7006 12044 7012 12056
rect 7064 12084 7070 12096
rect 7331 12087 7389 12093
rect 7331 12084 7343 12087
rect 7064 12056 7343 12084
rect 7064 12044 7070 12056
rect 7331 12053 7343 12056
rect 7377 12053 7389 12087
rect 7466 12084 7472 12096
rect 7427 12056 7472 12084
rect 7331 12047 7389 12053
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8662 12084 8668 12096
rect 8623 12056 8668 12084
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9033 12087 9091 12093
rect 9033 12053 9045 12087
rect 9079 12084 9091 12087
rect 9398 12084 9404 12096
rect 9079 12056 9404 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 9815 12087 9873 12093
rect 9815 12084 9827 12087
rect 9732 12056 9827 12084
rect 9732 12044 9738 12056
rect 9815 12053 9827 12056
rect 9861 12053 9873 12087
rect 10134 12084 10140 12096
rect 10095 12056 10140 12084
rect 9815 12047 9873 12053
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 15304 12084 15332 12124
rect 15470 12112 15476 12164
rect 15528 12152 15534 12164
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 15528 12124 15945 12152
rect 15528 12112 15534 12124
rect 15933 12121 15945 12124
rect 15979 12152 15991 12155
rect 17310 12152 17316 12164
rect 15979 12124 17316 12152
rect 15979 12121 15991 12124
rect 15933 12115 15991 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 18049 12087 18107 12093
rect 18049 12084 18061 12087
rect 15304 12056 18061 12084
rect 18049 12053 18061 12056
rect 18095 12053 18107 12087
rect 18049 12047 18107 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 2740 11852 2789 11880
rect 2740 11840 2746 11852
rect 2777 11849 2789 11852
rect 2823 11880 2835 11883
rect 3326 11880 3332 11892
rect 2823 11852 3332 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4157 11883 4215 11889
rect 4157 11880 4169 11883
rect 4120 11852 4169 11880
rect 4120 11840 4126 11852
rect 4157 11849 4169 11852
rect 4203 11849 4215 11883
rect 4157 11843 4215 11849
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4304 11852 4537 11880
rect 4304 11840 4310 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 4525 11843 4583 11849
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 5994 11880 6000 11892
rect 5859 11852 6000 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 2501 11815 2559 11821
rect 2501 11781 2513 11815
rect 2547 11812 2559 11815
rect 2866 11812 2872 11824
rect 2547 11784 2872 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2866 11772 2872 11784
rect 2924 11812 2930 11824
rect 3786 11812 3792 11824
rect 2924 11784 3792 11812
rect 2924 11772 2930 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1946 11744 1952 11756
rect 1535 11716 1952 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3418 11744 3424 11756
rect 3007 11716 3424 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 4540 11676 4568 11843
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6963 11883 7021 11889
rect 6963 11880 6975 11883
rect 6328 11852 6975 11880
rect 6328 11840 6334 11852
rect 6963 11849 6975 11852
rect 7009 11849 7021 11883
rect 6963 11843 7021 11849
rect 7377 11883 7435 11889
rect 7377 11849 7389 11883
rect 7423 11880 7435 11883
rect 7558 11880 7564 11892
rect 7423 11852 7564 11880
rect 7423 11849 7435 11852
rect 7377 11843 7435 11849
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8536 11852 8585 11880
rect 8536 11840 8542 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 8573 11843 8631 11849
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 9582 11880 9588 11892
rect 9543 11852 9588 11880
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 11790 11840 11796 11892
rect 11848 11880 11854 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 11848 11852 12173 11880
rect 11848 11840 11854 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12894 11880 12900 11892
rect 12855 11852 12900 11880
rect 12161 11843 12219 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 24719 11883 24777 11889
rect 24719 11880 24731 11883
rect 15344 11852 24731 11880
rect 15344 11840 15350 11852
rect 24719 11849 24731 11852
rect 24765 11849 24777 11883
rect 24719 11843 24777 11849
rect 6178 11812 6184 11824
rect 6091 11784 6184 11812
rect 6178 11772 6184 11784
rect 6236 11812 6242 11824
rect 7466 11812 7472 11824
rect 6236 11784 7472 11812
rect 6236 11772 6242 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 8386 11812 8392 11824
rect 8347 11784 8392 11812
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 8846 11772 8852 11824
rect 8904 11812 8910 11824
rect 10597 11815 10655 11821
rect 10597 11812 10609 11815
rect 8904 11784 10609 11812
rect 8904 11772 8910 11784
rect 10597 11781 10609 11784
rect 10643 11812 10655 11815
rect 14826 11812 14832 11824
rect 10643 11784 14832 11812
rect 10643 11781 10655 11784
rect 10597 11775 10655 11781
rect 6546 11744 6552 11756
rect 6507 11716 6552 11744
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7984 11716 8493 11744
rect 7984 11704 7990 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 4709 11679 4767 11685
rect 4709 11676 4721 11679
rect 3160 11648 4476 11676
rect 4540 11648 4721 11676
rect 3160 11620 3188 11648
rect 1578 11568 1584 11620
rect 1636 11608 1642 11620
rect 2133 11611 2191 11617
rect 1636 11580 1681 11608
rect 1636 11568 1642 11580
rect 2133 11577 2145 11611
rect 2179 11608 2191 11611
rect 3142 11608 3148 11620
rect 2179 11580 3148 11608
rect 2179 11577 2191 11580
rect 2133 11571 2191 11577
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3326 11617 3332 11620
rect 3323 11608 3332 11617
rect 3287 11580 3332 11608
rect 3323 11571 3332 11580
rect 3384 11608 3390 11620
rect 4246 11608 4252 11620
rect 3384 11580 4252 11608
rect 3326 11568 3332 11571
rect 3384 11568 3390 11580
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 4448 11608 4476 11648
rect 4709 11645 4721 11648
rect 4755 11645 4767 11679
rect 4709 11639 4767 11645
rect 5166 11636 5172 11688
rect 5224 11676 5230 11688
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 5224 11648 5273 11676
rect 5224 11636 5230 11648
rect 5261 11645 5273 11648
rect 5307 11676 5319 11679
rect 6454 11676 6460 11688
rect 5307 11648 6460 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 6860 11679 6918 11685
rect 6860 11645 6872 11679
rect 6906 11645 6918 11679
rect 6860 11639 6918 11645
rect 6638 11608 6644 11620
rect 4448 11580 6644 11608
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 6875 11608 6903 11639
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 8018 11676 8024 11688
rect 7064 11648 8024 11676
rect 7064 11636 7070 11648
rect 8018 11636 8024 11648
rect 8076 11676 8082 11688
rect 8260 11679 8318 11685
rect 8260 11676 8272 11679
rect 8076 11648 8272 11676
rect 8076 11636 8082 11648
rect 8260 11645 8272 11648
rect 8306 11676 8318 11679
rect 9398 11676 9404 11688
rect 8306 11648 9404 11676
rect 8306 11645 8318 11648
rect 8260 11639 8318 11645
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10042 11676 10048 11688
rect 9723 11648 10048 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10612 11676 10640 11775
rect 14826 11772 14832 11784
rect 14884 11772 14890 11824
rect 15470 11812 15476 11824
rect 15431 11784 15476 11812
rect 15470 11772 15476 11784
rect 15528 11772 15534 11824
rect 11698 11704 11704 11756
rect 11756 11744 11762 11756
rect 11793 11747 11851 11753
rect 11793 11744 11805 11747
rect 11756 11716 11805 11744
rect 11756 11704 11762 11716
rect 11793 11713 11805 11716
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 12894 11704 12900 11756
rect 12952 11744 12958 11756
rect 12952 11716 13445 11744
rect 12952 11704 12958 11716
rect 10686 11676 10692 11688
rect 10599 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11676 10750 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10744 11648 10793 11676
rect 10744 11636 10750 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11241 11679 11299 11685
rect 11241 11676 11253 11679
rect 10928 11648 11253 11676
rect 10928 11636 10934 11648
rect 11241 11645 11253 11648
rect 11287 11645 11299 11679
rect 11241 11639 11299 11645
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 11388 11648 13093 11676
rect 11388 11636 11394 11648
rect 13081 11645 13093 11648
rect 13127 11676 13139 11679
rect 13170 11676 13176 11688
rect 13127 11648 13176 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 6696 11580 6903 11608
rect 8113 11611 8171 11617
rect 6696 11568 6702 11580
rect 8113 11577 8125 11611
rect 8159 11608 8171 11611
rect 8386 11608 8392 11620
rect 8159 11580 8392 11608
rect 8159 11577 8171 11580
rect 8113 11571 8171 11577
rect 8220 11552 8248 11580
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 9766 11608 9772 11620
rect 9640 11580 9772 11608
rect 9640 11568 9646 11580
rect 9766 11568 9772 11580
rect 9824 11608 9830 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9824 11580 10149 11608
rect 9824 11568 9830 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 11514 11608 11520 11620
rect 11475 11580 11520 11608
rect 10137 11571 10195 11577
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 12986 11608 12992 11620
rect 12176 11580 12992 11608
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3016 11512 3893 11540
rect 3016 11500 3022 11512
rect 3881 11509 3893 11512
rect 3927 11509 3939 11543
rect 4798 11540 4804 11552
rect 4759 11512 4804 11540
rect 3881 11503 3939 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 7926 11540 7932 11552
rect 7887 11512 7932 11540
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8202 11500 8208 11552
rect 8260 11500 8266 11552
rect 9674 11500 9680 11552
rect 9732 11540 9738 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9732 11512 9873 11540
rect 9732 11500 9738 11512
rect 9861 11509 9873 11512
rect 9907 11540 9919 11543
rect 12176 11540 12204 11580
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 13417 11617 13445 11716
rect 14734 11704 14740 11756
rect 14792 11744 14798 11756
rect 14921 11747 14979 11753
rect 14921 11744 14933 11747
rect 14792 11716 14933 11744
rect 14792 11704 14798 11716
rect 14921 11713 14933 11716
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15620 11716 15945 11744
rect 15620 11704 15626 11716
rect 15933 11713 15945 11716
rect 15979 11744 15991 11747
rect 16393 11747 16451 11753
rect 16393 11744 16405 11747
rect 15979 11716 16405 11744
rect 15979 11713 15991 11716
rect 15933 11707 15991 11713
rect 16393 11713 16405 11716
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11676 16359 11679
rect 16485 11679 16543 11685
rect 16485 11676 16497 11679
rect 16347 11648 16497 11676
rect 16347 11645 16359 11648
rect 16301 11639 16359 11645
rect 16485 11645 16497 11648
rect 16531 11645 16543 11679
rect 16485 11639 16543 11645
rect 24648 11679 24706 11685
rect 24648 11645 24660 11679
rect 24694 11676 24706 11679
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24694 11648 25145 11676
rect 24694 11645 24706 11648
rect 24648 11639 24706 11645
rect 25133 11645 25145 11648
rect 25179 11676 25191 11679
rect 27614 11676 27620 11688
rect 25179 11648 27620 11676
rect 25179 11645 25191 11648
rect 25133 11639 25191 11645
rect 13402 11611 13460 11617
rect 13402 11577 13414 11611
rect 13448 11577 13460 11611
rect 14990 11611 15048 11617
rect 14990 11608 15002 11611
rect 13402 11571 13460 11577
rect 14200 11580 15002 11608
rect 14200 11552 14228 11580
rect 14990 11577 15002 11580
rect 15036 11577 15048 11611
rect 14990 11571 15048 11577
rect 15194 11568 15200 11620
rect 15252 11608 15258 11620
rect 16316 11608 16344 11639
rect 27614 11636 27620 11648
rect 27672 11636 27678 11688
rect 15252 11580 16344 11608
rect 15252 11568 15258 11580
rect 9907 11512 12204 11540
rect 14001 11543 14059 11549
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 14182 11540 14188 11552
rect 14047 11512 14188 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14366 11540 14372 11552
rect 14327 11512 14372 11540
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 18230 11540 18236 11552
rect 18191 11512 18236 11540
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2406 11336 2412 11348
rect 2363 11308 2412 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2516 11308 3433 11336
rect 2516 11280 2544 11308
rect 3421 11305 3433 11308
rect 3467 11336 3479 11339
rect 3602 11336 3608 11348
rect 3467 11308 3608 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 7285 11339 7343 11345
rect 4126 11308 5856 11336
rect 2498 11268 2504 11280
rect 2459 11240 2504 11268
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 2593 11271 2651 11277
rect 2593 11237 2605 11271
rect 2639 11268 2651 11271
rect 2958 11268 2964 11280
rect 2639 11240 2964 11268
rect 2639 11237 2651 11240
rect 2593 11231 2651 11237
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 3142 11268 3148 11280
rect 3103 11240 3148 11268
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 3970 11228 3976 11280
rect 4028 11268 4034 11280
rect 4126 11268 4154 11308
rect 4028 11240 4154 11268
rect 4028 11228 4034 11240
rect 4246 11228 4252 11280
rect 4304 11268 4310 11280
rect 4386 11271 4444 11277
rect 4386 11268 4398 11271
rect 4304 11240 4398 11268
rect 4304 11228 4310 11240
rect 4386 11237 4398 11240
rect 4432 11237 4444 11271
rect 4386 11231 4444 11237
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 5629 11271 5687 11277
rect 5629 11268 5641 11271
rect 5592 11240 5641 11268
rect 5592 11228 5598 11240
rect 5629 11237 5641 11240
rect 5675 11237 5687 11271
rect 5629 11231 5687 11237
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 2314 11200 2320 11212
rect 1510 11172 2320 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4614 11200 4620 11212
rect 4111 11172 4620 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5828 11209 5856 11308
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7466 11336 7472 11348
rect 7331 11308 7472 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7466 11296 7472 11308
rect 7524 11296 7530 11348
rect 9950 11336 9956 11348
rect 9911 11308 9956 11336
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 13722 11336 13728 11348
rect 13683 11308 13728 11336
rect 13722 11296 13728 11308
rect 13780 11336 13786 11348
rect 13909 11339 13967 11345
rect 13909 11336 13921 11339
rect 13780 11308 13921 11336
rect 13780 11296 13786 11308
rect 13909 11305 13921 11308
rect 13955 11305 13967 11339
rect 13909 11299 13967 11305
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14240 11308 14933 11336
rect 14240 11296 14246 11308
rect 14921 11305 14933 11308
rect 14967 11336 14979 11339
rect 15194 11336 15200 11348
rect 14967 11308 15200 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 15378 11336 15384 11348
rect 15339 11308 15384 11336
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 8573 11271 8631 11277
rect 8573 11237 8585 11271
rect 8619 11268 8631 11271
rect 9858 11268 9864 11280
rect 8619 11240 9864 11268
rect 8619 11237 8631 11240
rect 8573 11231 8631 11237
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 11330 11268 11336 11280
rect 10192 11240 11100 11268
rect 11291 11240 11336 11268
rect 10192 11228 10198 11240
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 6086 11200 6092 11212
rect 5859 11172 6092 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 6086 11160 6092 11172
rect 6144 11160 6150 11212
rect 6362 11200 6368 11212
rect 6323 11172 6368 11200
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6917 11203 6975 11209
rect 6917 11169 6929 11203
rect 6963 11200 6975 11203
rect 7006 11200 7012 11212
rect 6963 11172 7012 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7616 11172 7849 11200
rect 7616 11160 7622 11172
rect 7837 11169 7849 11172
rect 7883 11200 7895 11203
rect 8662 11200 8668 11212
rect 7883 11172 8668 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8662 11160 8668 11172
rect 8720 11160 8726 11212
rect 10686 11200 10692 11212
rect 10647 11172 10692 11200
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11072 11209 11100 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 12523 11271 12581 11277
rect 12523 11268 12535 11271
rect 12400 11240 12535 11268
rect 12400 11228 12406 11240
rect 12523 11237 12535 11240
rect 12569 11268 12581 11271
rect 12894 11268 12900 11280
rect 12569 11240 12900 11268
rect 12569 11237 12581 11240
rect 12523 11231 12581 11237
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 16853 11271 16911 11277
rect 16853 11268 16865 11271
rect 14424 11240 16865 11268
rect 14424 11228 14430 11240
rect 16853 11237 16865 11240
rect 16899 11237 16911 11271
rect 16853 11231 16911 11237
rect 11057 11203 11115 11209
rect 11057 11169 11069 11203
rect 11103 11200 11115 11203
rect 11238 11200 11244 11212
rect 11103 11172 11244 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11572 11172 12173 11200
rect 11572 11160 11578 11172
rect 12161 11169 12173 11172
rect 12207 11200 12219 11203
rect 12250 11200 12256 11212
rect 12207 11172 12256 11200
rect 12207 11169 12219 11172
rect 12161 11163 12219 11169
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11169 15347 11203
rect 15746 11200 15752 11212
rect 15707 11172 15752 11200
rect 15289 11163 15347 11169
rect 3881 11135 3939 11141
rect 2745 11104 3188 11132
rect 1535 11067 1593 11073
rect 1535 11033 1547 11067
rect 1581 11064 1593 11067
rect 2745 11064 2773 11104
rect 1581 11036 2773 11064
rect 3160 11064 3188 11104
rect 3881 11101 3893 11135
rect 3927 11132 3939 11135
rect 4338 11132 4344 11144
rect 3927 11104 4344 11132
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 6273 11135 6331 11141
rect 6273 11132 6285 11135
rect 4488 11104 6285 11132
rect 4488 11092 4494 11104
rect 6273 11101 6285 11104
rect 6319 11101 6331 11135
rect 7024 11132 7052 11160
rect 7984 11135 8042 11141
rect 7984 11132 7996 11135
rect 7024 11104 7996 11132
rect 6273 11095 6331 11101
rect 7984 11101 7996 11104
rect 8030 11101 8042 11135
rect 7984 11095 8042 11101
rect 8110 11092 8116 11144
rect 8168 11132 8174 11144
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 8168 11104 8217 11132
rect 8168 11092 8174 11104
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 11698 11092 11704 11144
rect 11756 11132 11762 11144
rect 15304 11132 15332 11163
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 16942 11200 16948 11212
rect 16903 11172 16948 11200
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 15838 11132 15844 11144
rect 11756 11104 15844 11132
rect 11756 11092 11762 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 6178 11064 6184 11076
rect 3160 11036 6184 11064
rect 1581 11033 1593 11036
rect 1535 11027 1593 11033
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 7653 11067 7711 11073
rect 7653 11033 7665 11067
rect 7699 11064 7711 11067
rect 8386 11064 8392 11076
rect 7699 11036 8392 11064
rect 7699 11033 7711 11036
rect 7653 11027 7711 11033
rect 8386 11024 8392 11036
rect 8444 11024 8450 11076
rect 1946 10996 1952 11008
rect 1859 10968 1952 10996
rect 1946 10956 1952 10968
rect 2004 10996 2010 11008
rect 3694 10996 3700 11008
rect 2004 10968 3700 10996
rect 2004 10956 2010 10968
rect 3694 10956 3700 10968
rect 3752 10956 3758 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4985 10999 5043 11005
rect 4985 10996 4997 10999
rect 3844 10968 4997 10996
rect 3844 10956 3850 10968
rect 4985 10965 4997 10968
rect 5031 10965 5043 10999
rect 4985 10959 5043 10965
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 5261 10999 5319 11005
rect 5261 10996 5273 10999
rect 5224 10968 5273 10996
rect 5224 10956 5230 10968
rect 5261 10965 5273 10968
rect 5307 10965 5319 10999
rect 5261 10959 5319 10965
rect 7834 10956 7840 11008
rect 7892 10996 7898 11008
rect 8113 10999 8171 11005
rect 8113 10996 8125 10999
rect 7892 10968 8125 10996
rect 7892 10956 7898 10968
rect 8113 10965 8125 10968
rect 8159 10965 8171 10999
rect 8113 10959 8171 10965
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 8849 10999 8907 11005
rect 8849 10996 8861 10999
rect 8536 10968 8861 10996
rect 8536 10956 8542 10968
rect 8849 10965 8861 10968
rect 8895 10965 8907 10999
rect 8849 10959 8907 10965
rect 9493 10999 9551 11005
rect 9493 10965 9505 10999
rect 9539 10996 9551 10999
rect 9766 10996 9772 11008
rect 9539 10968 9772 10996
rect 9539 10965 9551 10968
rect 9493 10959 9551 10965
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 10042 10956 10048 11008
rect 10100 10996 10106 11008
rect 10229 10999 10287 11005
rect 10229 10996 10241 10999
rect 10100 10968 10241 10996
rect 10100 10956 10106 10968
rect 10229 10965 10241 10968
rect 10275 10965 10287 10999
rect 13078 10996 13084 11008
rect 13039 10968 13084 10996
rect 10229 10959 10287 10965
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14461 10999 14519 11005
rect 14461 10996 14473 10999
rect 13780 10968 14473 10996
rect 13780 10956 13786 10968
rect 14461 10965 14473 10968
rect 14507 10996 14519 10999
rect 14734 10996 14740 11008
rect 14507 10968 14740 10996
rect 14507 10965 14519 10968
rect 14461 10959 14519 10965
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4157 10795 4215 10801
rect 4157 10792 4169 10795
rect 4120 10764 4169 10792
rect 4120 10752 4126 10764
rect 4157 10761 4169 10764
rect 4203 10792 4215 10795
rect 4246 10792 4252 10804
rect 4203 10764 4252 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4522 10792 4528 10804
rect 4483 10764 4528 10792
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6362 10792 6368 10804
rect 5951 10764 6368 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 7006 10792 7012 10804
rect 6687 10764 7012 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9456 10764 9965 10792
rect 9456 10752 9462 10764
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 10192 10764 10241 10792
rect 10192 10752 10198 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10686 10792 10692 10804
rect 10647 10764 10692 10792
rect 10229 10755 10287 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 12342 10792 12348 10804
rect 12299 10764 12348 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 13078 10792 13084 10804
rect 12851 10764 13084 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 13078 10752 13084 10764
rect 13136 10792 13142 10804
rect 13446 10792 13452 10804
rect 13136 10764 13452 10792
rect 13136 10752 13142 10764
rect 13446 10752 13452 10764
rect 13504 10792 13510 10804
rect 13504 10764 13814 10792
rect 13504 10752 13510 10764
rect 3602 10724 3608 10736
rect 3563 10696 3608 10724
rect 3602 10684 3608 10696
rect 3660 10684 3666 10736
rect 3694 10684 3700 10736
rect 3752 10724 3758 10736
rect 3752 10696 6868 10724
rect 3752 10684 3758 10696
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3418 10656 3424 10668
rect 3099 10628 3424 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 6086 10616 6092 10668
rect 6144 10656 6150 10668
rect 6840 10665 6868 10696
rect 7190 10684 7196 10736
rect 7248 10724 7254 10736
rect 7561 10727 7619 10733
rect 7561 10724 7573 10727
rect 7248 10696 7573 10724
rect 7248 10684 7254 10696
rect 7561 10693 7573 10696
rect 7607 10724 7619 10727
rect 8343 10727 8401 10733
rect 8343 10724 8355 10727
rect 7607 10696 8355 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 8343 10693 8355 10696
rect 8389 10693 8401 10727
rect 8478 10724 8484 10736
rect 8439 10696 8484 10724
rect 8343 10687 8401 10693
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 9674 10724 9680 10736
rect 9048 10696 9680 10724
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 6144 10628 6193 10656
rect 6144 10616 6150 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10557 2099 10591
rect 2041 10551 2099 10557
rect 2056 10464 2084 10551
rect 4522 10548 4528 10600
rect 4580 10588 4586 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4580 10560 4629 10588
rect 4580 10548 4586 10560
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 5166 10588 5172 10600
rect 5127 10560 5172 10588
rect 4617 10551 4675 10557
rect 3145 10523 3203 10529
rect 3145 10489 3157 10523
rect 3191 10489 3203 10523
rect 4632 10520 4660 10551
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 6196 10588 6224 10619
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 8110 10656 8116 10668
rect 7524 10628 8116 10656
rect 7524 10616 7530 10628
rect 8110 10616 8116 10628
rect 8168 10656 8174 10668
rect 8570 10656 8576 10668
rect 8168 10628 8576 10656
rect 8168 10616 8174 10628
rect 8570 10616 8576 10628
rect 8628 10656 8634 10668
rect 9048 10656 9076 10696
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 13170 10724 13176 10736
rect 13131 10696 13176 10724
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 13786 10724 13814 10764
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14553 10795 14611 10801
rect 14553 10792 14565 10795
rect 14148 10764 14565 10792
rect 14148 10752 14154 10764
rect 14553 10761 14565 10764
rect 14599 10792 14611 10795
rect 14645 10795 14703 10801
rect 14645 10792 14657 10795
rect 14599 10764 14657 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14645 10761 14657 10764
rect 14691 10761 14703 10795
rect 15838 10792 15844 10804
rect 15799 10764 15844 10792
rect 14645 10755 14703 10761
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 16531 10795 16589 10801
rect 16531 10761 16543 10795
rect 16577 10792 16589 10795
rect 19334 10792 19340 10804
rect 16577 10764 19340 10792
rect 16577 10761 16589 10764
rect 16531 10755 16589 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 16853 10727 16911 10733
rect 16853 10724 16865 10727
rect 13786 10696 16865 10724
rect 16853 10693 16865 10696
rect 16899 10724 16911 10727
rect 16942 10724 16948 10736
rect 16899 10696 16948 10724
rect 16899 10693 16911 10696
rect 16853 10687 16911 10693
rect 16942 10684 16948 10696
rect 17000 10684 17006 10736
rect 8628 10628 9076 10656
rect 9309 10659 9367 10665
rect 8628 10616 8634 10628
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9950 10656 9956 10668
rect 9355 10628 9956 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 8205 10591 8263 10597
rect 6196 10560 8156 10588
rect 6546 10520 6552 10532
rect 4632 10492 6552 10520
rect 3145 10483 3203 10489
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 2409 10455 2467 10461
rect 2409 10452 2421 10455
rect 2096 10424 2421 10452
rect 2096 10412 2102 10424
rect 2409 10421 2421 10424
rect 2455 10421 2467 10455
rect 2409 10415 2467 10421
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 3050 10452 3056 10464
rect 2915 10424 3056 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 3050 10412 3056 10424
rect 3108 10452 3114 10464
rect 3160 10452 3188 10483
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 3108 10424 3188 10452
rect 3108 10412 3114 10424
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 4580 10424 4721 10452
rect 4580 10412 4586 10424
rect 4709 10421 4721 10424
rect 4755 10421 4767 10455
rect 4709 10415 4767 10421
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 7834 10452 7840 10464
rect 7708 10424 7840 10452
rect 7708 10412 7714 10424
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 8128 10452 8156 10560
rect 8205 10557 8217 10591
rect 8251 10588 8263 10591
rect 9324 10588 9352 10619
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 13412 10628 14289 10656
rect 13412 10616 13418 10628
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 8251 10560 9352 10588
rect 9769 10591 9827 10597
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 9769 10557 9781 10591
rect 9815 10588 9827 10591
rect 9858 10588 9864 10600
rect 9815 10560 9864 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10962 10588 10968 10600
rect 10923 10560 10968 10588
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11238 10588 11244 10600
rect 11199 10560 11244 10588
rect 11238 10548 11244 10560
rect 11296 10588 11302 10600
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11296 10560 11805 10588
rect 11296 10548 11302 10560
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14553 10591 14611 10597
rect 14056 10560 14101 10588
rect 14056 10548 14062 10560
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 14829 10591 14887 10597
rect 14829 10588 14841 10591
rect 14599 10560 14841 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 14829 10557 14841 10560
rect 14875 10557 14887 10591
rect 15286 10588 15292 10600
rect 15247 10560 15292 10588
rect 14829 10551 14887 10557
rect 15286 10548 15292 10560
rect 15344 10588 15350 10600
rect 15746 10588 15752 10600
rect 15344 10560 15752 10588
rect 15344 10548 15350 10560
rect 15746 10548 15752 10560
rect 15804 10588 15810 10600
rect 23750 10597 23756 10600
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 15804 10560 16221 10588
rect 15804 10548 15810 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16428 10591 16486 10597
rect 16428 10557 16440 10591
rect 16474 10588 16486 10591
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 16474 10560 17233 10588
rect 16474 10557 16486 10560
rect 16428 10551 16486 10557
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 23728 10591 23756 10597
rect 23728 10588 23740 10591
rect 23663 10560 23740 10588
rect 17221 10551 17279 10557
rect 23728 10557 23740 10560
rect 23808 10588 23814 10600
rect 24121 10591 24179 10597
rect 24121 10588 24133 10591
rect 23808 10560 24133 10588
rect 23728 10551 23756 10557
rect 8938 10520 8944 10532
rect 8899 10492 8944 10520
rect 8938 10480 8944 10492
rect 8996 10480 9002 10532
rect 11514 10520 11520 10532
rect 9508 10492 9674 10520
rect 11475 10492 11520 10520
rect 9508 10452 9536 10492
rect 8128 10424 9536 10452
rect 9646 10452 9674 10492
rect 11514 10480 11520 10492
rect 11572 10480 11578 10532
rect 13354 10520 13360 10532
rect 13315 10492 13360 10520
rect 13354 10480 13360 10492
rect 13412 10480 13418 10532
rect 13446 10480 13452 10532
rect 13504 10520 13510 10532
rect 14016 10520 14044 10548
rect 16443 10520 16471 10551
rect 23750 10548 23756 10551
rect 23808 10548 23814 10560
rect 24121 10557 24133 10560
rect 24167 10557 24179 10591
rect 24121 10551 24179 10557
rect 13504 10492 13549 10520
rect 14016 10492 16471 10520
rect 13504 10480 13510 10492
rect 10962 10452 10968 10464
rect 9646 10424 10968 10452
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14792 10424 14933 10452
rect 14792 10412 14798 10424
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 23799 10455 23857 10461
rect 23799 10452 23811 10455
rect 18196 10424 23811 10452
rect 18196 10412 18202 10424
rect 23799 10421 23811 10424
rect 23845 10421 23857 10455
rect 23799 10415 23857 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 2280 10220 4721 10248
rect 2280 10208 2286 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 4709 10211 4767 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 6512 10220 7880 10248
rect 6512 10208 6518 10220
rect 1670 10140 1676 10192
rect 1728 10180 1734 10192
rect 1765 10183 1823 10189
rect 1765 10180 1777 10183
rect 1728 10152 1777 10180
rect 1728 10140 1734 10152
rect 1765 10149 1777 10152
rect 1811 10149 1823 10183
rect 2958 10180 2964 10192
rect 2919 10152 2964 10180
rect 1765 10143 1823 10149
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 7006 10180 7012 10192
rect 6967 10152 7012 10180
rect 7006 10140 7012 10152
rect 7064 10180 7070 10192
rect 7852 10180 7880 10220
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8570 10248 8576 10260
rect 8168 10220 8576 10248
rect 8168 10208 8174 10220
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8938 10208 8944 10260
rect 8996 10248 9002 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 8996 10220 9321 10248
rect 8996 10208 9002 10220
rect 9309 10217 9321 10220
rect 9355 10248 9367 10251
rect 9490 10248 9496 10260
rect 9355 10220 9496 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 12250 10248 12256 10260
rect 12211 10220 12256 10248
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12400 10220 12909 10248
rect 12400 10208 12406 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 12897 10211 12955 10217
rect 10413 10183 10471 10189
rect 10413 10180 10425 10183
rect 7064 10152 7751 10180
rect 7852 10152 10425 10180
rect 7064 10140 7070 10152
rect 2682 10112 2688 10124
rect 2595 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10112 2746 10124
rect 4522 10112 4528 10124
rect 2740 10084 4528 10112
rect 2740 10072 2746 10084
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 4893 10115 4951 10121
rect 4893 10081 4905 10115
rect 4939 10081 4951 10115
rect 5166 10112 5172 10124
rect 5127 10084 5172 10112
rect 4893 10075 4951 10081
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 1762 10044 1768 10056
rect 1719 10016 1768 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 1762 10004 1768 10016
rect 1820 10004 1826 10056
rect 2314 10004 2320 10056
rect 2372 10044 2378 10056
rect 3694 10044 3700 10056
rect 2372 10016 3700 10044
rect 2372 10004 2378 10016
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 4798 10004 4804 10056
rect 4856 10044 4862 10056
rect 4908 10044 4936 10075
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 6178 10112 6184 10124
rect 6139 10084 6184 10112
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 7723 10121 7751 10152
rect 10413 10149 10425 10152
rect 10459 10149 10471 10183
rect 10413 10143 10471 10149
rect 10873 10183 10931 10189
rect 10873 10149 10885 10183
rect 10919 10180 10931 10183
rect 10962 10180 10968 10192
rect 10919 10152 10968 10180
rect 10919 10149 10931 10152
rect 10873 10143 10931 10149
rect 10962 10140 10968 10152
rect 11020 10180 11026 10192
rect 14458 10180 14464 10192
rect 11020 10152 12848 10180
rect 11020 10140 11026 10152
rect 12820 10124 12848 10152
rect 13096 10152 14464 10180
rect 7708 10115 7766 10121
rect 7708 10081 7720 10115
rect 7754 10081 7766 10115
rect 7708 10075 7766 10081
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 8444 10084 9689 10112
rect 8444 10072 8450 10084
rect 9677 10081 9689 10084
rect 9723 10112 9735 10115
rect 10134 10112 10140 10124
rect 9723 10084 10140 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 11330 10112 11336 10124
rect 11291 10084 11336 10112
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 12802 10072 12808 10124
rect 12860 10112 12866 10124
rect 13096 10121 13124 10152
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 12860 10084 13093 10112
rect 12860 10072 12866 10084
rect 13081 10081 13093 10084
rect 13127 10081 13139 10115
rect 13262 10112 13268 10124
rect 13223 10084 13268 10112
rect 13081 10075 13139 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 15930 10112 15936 10124
rect 15891 10084 15936 10112
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 7282 10044 7288 10056
rect 4856 10016 7288 10044
rect 4856 10004 4862 10016
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 7926 10044 7932 10056
rect 7887 10016 7932 10044
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 10042 10044 10048 10056
rect 10003 10016 10048 10044
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 10330 10016 11253 10044
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 2590 9976 2596 9988
rect 2271 9948 2596 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 2590 9936 2596 9948
rect 2648 9936 2654 9988
rect 4341 9979 4399 9985
rect 4341 9945 4353 9979
rect 4387 9976 4399 9979
rect 4614 9976 4620 9988
rect 4387 9948 4620 9976
rect 4387 9945 4399 9948
rect 4341 9939 4399 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 8478 9976 8484 9988
rect 7852 9948 8484 9976
rect 7852 9920 7880 9948
rect 8478 9936 8484 9948
rect 8536 9976 8542 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8536 9948 8953 9976
rect 8536 9936 8542 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 9732 9948 9965 9976
rect 9732 9936 9738 9948
rect 9953 9945 9965 9948
rect 9999 9976 10011 9979
rect 10330 9976 10358 10016
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 11348 10044 11376 10072
rect 18230 10044 18236 10056
rect 11348 10016 18236 10044
rect 11241 10007 11299 10013
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 9999 9948 10358 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 3418 9908 3424 9920
rect 3379 9880 3424 9908
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8018 9908 8024 9920
rect 7979 9880 8024 9908
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9858 9917 9864 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8444 9880 8585 9908
rect 8444 9868 8450 9880
rect 8573 9877 8585 9880
rect 8619 9877 8631 9911
rect 8573 9871 8631 9877
rect 9842 9911 9864 9917
rect 9842 9877 9854 9911
rect 9842 9871 9864 9877
rect 9858 9868 9864 9871
rect 9916 9868 9922 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 11204 9880 14841 9908
rect 11204 9868 11210 9880
rect 14829 9877 14841 9880
rect 14875 9908 14887 9911
rect 15286 9908 15292 9920
rect 14875 9880 15292 9908
rect 14875 9877 14887 9880
rect 14829 9871 14887 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1670 9704 1676 9716
rect 1631 9676 1676 9704
rect 1670 9664 1676 9676
rect 1728 9664 1734 9716
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 3789 9707 3847 9713
rect 3789 9704 3801 9707
rect 3292 9676 3801 9704
rect 3292 9664 3298 9676
rect 3789 9673 3801 9676
rect 3835 9704 3847 9707
rect 5905 9707 5963 9713
rect 3835 9676 4154 9704
rect 3835 9673 3847 9676
rect 3789 9667 3847 9673
rect 2133 9571 2191 9577
rect 2133 9537 2145 9571
rect 2179 9568 2191 9571
rect 2682 9568 2688 9580
rect 2179 9540 2688 9568
rect 2179 9537 2191 9540
rect 2133 9531 2191 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 4126 9568 4154 9676
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6178 9704 6184 9716
rect 5951 9676 6184 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 6546 9704 6552 9716
rect 6507 9676 6552 9704
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8386 9704 8392 9716
rect 7616 9676 8392 9704
rect 7616 9664 7622 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 10870 9664 10876 9716
rect 10928 9704 10934 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 10928 9676 12173 9704
rect 10928 9664 10934 9676
rect 12161 9673 12173 9676
rect 12207 9704 12219 9707
rect 13262 9704 13268 9716
rect 12207 9676 13268 9704
rect 12207 9673 12219 9676
rect 12161 9667 12219 9673
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 14369 9707 14427 9713
rect 14369 9704 14381 9707
rect 13786 9676 14381 9704
rect 4249 9639 4307 9645
rect 4249 9605 4261 9639
rect 4295 9636 4307 9639
rect 5166 9636 5172 9648
rect 4295 9608 5172 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 11330 9636 11336 9648
rect 7800 9608 11336 9636
rect 7800 9596 7806 9608
rect 11330 9596 11336 9608
rect 11388 9636 11394 9648
rect 11609 9639 11667 9645
rect 11609 9636 11621 9639
rect 11388 9608 11621 9636
rect 11388 9596 11394 9608
rect 11609 9605 11621 9608
rect 11655 9605 11667 9639
rect 12894 9636 12900 9648
rect 12855 9608 12900 9636
rect 11609 9599 11667 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 4126 9540 4813 9568
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6273 9571 6331 9577
rect 6273 9568 6285 9571
rect 6144 9540 6285 9568
rect 6144 9528 6150 9540
rect 6273 9537 6285 9540
rect 6319 9568 6331 9571
rect 9030 9568 9036 9580
rect 6319 9540 7420 9568
rect 8943 9540 9036 9568
rect 6319 9537 6331 9540
rect 6273 9531 6331 9537
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 7392 9509 7420 9540
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6604 9472 6837 9500
rect 6604 9460 6610 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 8018 9500 8024 9512
rect 7423 9472 8024 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 1949 9435 2007 9441
rect 1949 9432 1961 9435
rect 1912 9404 1961 9432
rect 1912 9392 1918 9404
rect 1949 9401 1961 9404
rect 1995 9432 2007 9435
rect 2454 9435 2512 9441
rect 2454 9432 2466 9435
rect 1995 9404 2466 9432
rect 1995 9401 2007 9404
rect 1949 9395 2007 9401
rect 2454 9401 2466 9404
rect 2500 9401 2512 9435
rect 2454 9395 2512 9401
rect 4617 9435 4675 9441
rect 4617 9401 4629 9435
rect 4663 9432 4675 9435
rect 4890 9432 4896 9444
rect 4663 9404 4896 9432
rect 4663 9401 4675 9404
rect 4617 9395 4675 9401
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 5445 9435 5503 9441
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 6730 9432 6736 9444
rect 5491 9404 6736 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6840 9432 6868 9463
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8956 9432 8984 9540
rect 9030 9528 9036 9540
rect 9088 9568 9094 9580
rect 10689 9571 10747 9577
rect 9088 9540 9168 9568
rect 9088 9528 9094 9540
rect 9140 9509 9168 9540
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 10778 9568 10784 9580
rect 10735 9540 10784 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 13081 9571 13139 9577
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13786 9568 13814 9676
rect 14369 9673 14381 9676
rect 14415 9704 14427 9707
rect 15378 9704 15384 9716
rect 14415 9676 15384 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16117 9707 16175 9713
rect 16117 9704 16129 9707
rect 15988 9676 16129 9704
rect 15988 9664 15994 9676
rect 16117 9673 16129 9676
rect 16163 9673 16175 9707
rect 16117 9667 16175 9673
rect 16485 9639 16543 9645
rect 16485 9636 16497 9639
rect 15212 9608 16497 9636
rect 13127 9540 13814 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 15212 9577 15240 9608
rect 16485 9605 16497 9608
rect 16531 9605 16543 9639
rect 16485 9599 16543 9605
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14700 9540 15209 9568
rect 14700 9528 14706 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15654 9568 15660 9580
rect 15615 9540 15660 9568
rect 15197 9531 15255 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9490 9500 9496 9512
rect 9451 9472 9496 9500
rect 9125 9463 9183 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 14047 9472 14933 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 9766 9432 9772 9444
rect 6840 9404 8984 9432
rect 9727 9404 9772 9432
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 10781 9435 10839 9441
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 10870 9432 10876 9444
rect 10827 9404 10876 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 3053 9367 3111 9373
rect 3053 9364 3065 9367
rect 2096 9336 3065 9364
rect 2096 9324 2102 9336
rect 3053 9333 3065 9336
rect 3099 9333 3111 9367
rect 6914 9364 6920 9376
rect 6875 9336 6920 9364
rect 3053 9327 3111 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7708 9336 7849 9364
rect 7708 9324 7714 9336
rect 7837 9333 7849 9336
rect 7883 9364 7895 9367
rect 7926 9364 7932 9376
rect 7883 9336 7932 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8297 9367 8355 9373
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8386 9364 8392 9376
rect 8343 9336 8392 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8941 9367 8999 9373
rect 8941 9333 8953 9367
rect 8987 9364 8999 9367
rect 9674 9364 9680 9376
rect 8987 9336 9680 9364
rect 8987 9333 8999 9336
rect 8941 9327 8999 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10505 9367 10563 9373
rect 10505 9333 10517 9367
rect 10551 9364 10563 9367
rect 10796 9364 10824 9395
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 11333 9435 11391 9441
rect 11333 9401 11345 9435
rect 11379 9432 11391 9435
rect 11882 9432 11888 9444
rect 11379 9404 11888 9432
rect 11379 9401 11391 9404
rect 11333 9395 11391 9401
rect 11882 9392 11888 9404
rect 11940 9392 11946 9444
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 13402 9435 13460 9441
rect 13402 9432 13414 9435
rect 12952 9404 13414 9432
rect 12952 9392 12958 9404
rect 13402 9401 13414 9404
rect 13448 9401 13460 9435
rect 13402 9395 13460 9401
rect 10551 9336 10824 9364
rect 14936 9364 14964 9463
rect 15289 9435 15347 9441
rect 15289 9401 15301 9435
rect 15335 9432 15347 9435
rect 16942 9432 16948 9444
rect 15335 9404 16948 9432
rect 15335 9401 15347 9404
rect 15289 9395 15347 9401
rect 15304 9364 15332 9395
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 14936 9336 15332 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 4709 9163 4767 9169
rect 4709 9160 4721 9163
rect 4580 9132 4721 9160
rect 4580 9120 4586 9132
rect 4709 9129 4721 9132
rect 4755 9160 4767 9163
rect 4798 9160 4804 9172
rect 4755 9132 4804 9160
rect 4755 9129 4767 9132
rect 4709 9123 4767 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 5258 9160 5264 9172
rect 5219 9132 5264 9160
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 9030 9160 9036 9172
rect 8991 9132 9036 9160
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 12434 9160 12440 9172
rect 11572 9132 12440 9160
rect 11572 9120 11578 9132
rect 12434 9120 12440 9132
rect 12492 9120 12498 9172
rect 12802 9160 12808 9172
rect 12763 9132 12808 9160
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 14001 9163 14059 9169
rect 14001 9129 14013 9163
rect 14047 9160 14059 9163
rect 15286 9160 15292 9172
rect 14047 9132 15292 9160
rect 14047 9129 14059 9132
rect 14001 9123 14059 9129
rect 15286 9120 15292 9132
rect 15344 9160 15350 9172
rect 15930 9160 15936 9172
rect 15344 9132 15936 9160
rect 15344 9120 15350 9132
rect 2038 9092 2044 9104
rect 1999 9064 2044 9092
rect 2038 9052 2044 9064
rect 2096 9052 2102 9104
rect 2590 9092 2596 9104
rect 2551 9064 2596 9092
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 7190 9092 7196 9104
rect 7151 9064 7196 9092
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 11330 9092 11336 9104
rect 11291 9064 11336 9092
rect 11330 9052 11336 9064
rect 11388 9052 11394 9104
rect 12894 9052 12900 9104
rect 12952 9092 12958 9104
rect 15488 9101 15516 9132
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 13402 9095 13460 9101
rect 13402 9092 13414 9095
rect 12952 9064 13414 9092
rect 12952 9052 12958 9064
rect 13402 9061 13414 9064
rect 13448 9061 13460 9095
rect 13402 9055 13460 9061
rect 15473 9095 15531 9101
rect 15473 9061 15485 9095
rect 15519 9061 15531 9095
rect 15473 9055 15531 9061
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 6641 9027 6699 9033
rect 6641 9024 6653 9027
rect 6328 8996 6653 9024
rect 6328 8984 6334 8996
rect 6641 8993 6653 8996
rect 6687 8993 6699 9027
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6641 8987 6699 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 7926 9024 7932 9036
rect 7340 8996 7932 9024
rect 7340 8984 7346 8996
rect 7926 8984 7932 8996
rect 7984 9024 7990 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7984 8996 8033 9024
rect 7984 8984 7990 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 9024 8631 9027
rect 8938 9024 8944 9036
rect 8619 8996 8944 9024
rect 8619 8993 8631 8996
rect 8573 8987 8631 8993
rect 8938 8984 8944 8996
rect 8996 9024 9002 9036
rect 9490 9024 9496 9036
rect 8996 8996 9496 9024
rect 8996 8984 9002 8996
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 16942 9024 16948 9036
rect 16903 8996 16948 9024
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4672 8928 4905 8956
rect 4672 8916 4678 8928
rect 4893 8925 4905 8928
rect 4939 8956 4951 8959
rect 6914 8956 6920 8968
rect 4939 8928 6920 8956
rect 4939 8925 4951 8928
rect 4893 8919 4951 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9950 8956 9956 8968
rect 8803 8928 9956 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11606 8956 11612 8968
rect 11287 8928 11612 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 11882 8956 11888 8968
rect 11843 8928 11888 8956
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 13078 8956 13084 8968
rect 13039 8928 13084 8956
rect 13078 8916 13084 8928
rect 13136 8956 13142 8968
rect 14734 8956 14740 8968
rect 13136 8928 14740 8956
rect 13136 8916 13142 8928
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 15105 8959 15163 8965
rect 15105 8925 15117 8959
rect 15151 8956 15163 8959
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15151 8928 15393 8956
rect 15151 8925 15163 8928
rect 15105 8919 15163 8925
rect 15381 8925 15393 8928
rect 15427 8956 15439 8959
rect 15654 8956 15660 8968
rect 15427 8928 15660 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16114 8956 16120 8968
rect 16071 8928 16120 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16264 8928 16865 8956
rect 16264 8916 16270 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 10042 8888 10048 8900
rect 8720 8860 10048 8888
rect 8720 8848 8726 8860
rect 10042 8848 10048 8860
rect 10100 8888 10106 8900
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 10100 8860 10149 8888
rect 10100 8848 10106 8860
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 1762 8820 1768 8832
rect 1719 8792 1768 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 1762 8780 1768 8792
rect 1820 8820 1826 8832
rect 3970 8820 3976 8832
rect 1820 8792 3976 8820
rect 1820 8780 1826 8792
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5592 8792 5825 8820
rect 5592 8780 5598 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 7834 8820 7840 8832
rect 7699 8792 7840 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 7834 8780 7840 8792
rect 7892 8820 7898 8832
rect 8018 8820 8024 8832
rect 7892 8792 8024 8820
rect 7892 8780 7898 8792
rect 8018 8780 8024 8792
rect 8076 8820 8082 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 8076 8792 9873 8820
rect 8076 8780 8082 8792
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 10502 8820 10508 8832
rect 10463 8792 10508 8820
rect 9861 8783 9919 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 10873 8823 10931 8829
rect 10873 8820 10885 8823
rect 10836 8792 10885 8820
rect 10836 8780 10842 8792
rect 10873 8789 10885 8792
rect 10919 8789 10931 8823
rect 14274 8820 14280 8832
rect 14235 8792 14280 8820
rect 10873 8783 10931 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4893 8619 4951 8625
rect 4893 8616 4905 8619
rect 4571 8588 4905 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4893 8585 4905 8588
rect 4939 8616 4951 8619
rect 5258 8616 5264 8628
rect 4939 8588 5264 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 2314 8508 2320 8560
rect 2372 8548 2378 8560
rect 4430 8548 4436 8560
rect 2372 8520 4436 8548
rect 2372 8508 2378 8520
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 2004 8452 3433 8480
rect 2004 8440 2010 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3970 8480 3976 8492
rect 3931 8452 3976 8480
rect 3421 8443 3479 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 2222 8412 2228 8424
rect 1811 8384 2228 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 2133 8347 2191 8353
rect 2133 8344 2145 8347
rect 1912 8316 2145 8344
rect 1912 8304 1918 8316
rect 2133 8313 2145 8316
rect 2179 8344 2191 8347
rect 2587 8347 2645 8353
rect 2587 8344 2599 8347
rect 2179 8316 2599 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 2587 8313 2599 8316
rect 2633 8344 2645 8347
rect 2958 8344 2964 8356
rect 2633 8316 2964 8344
rect 2633 8313 2645 8316
rect 2587 8307 2645 8313
rect 2958 8304 2964 8316
rect 3016 8344 3022 8356
rect 4062 8344 4068 8356
rect 3016 8316 4068 8344
rect 3016 8304 3022 8316
rect 4062 8304 4068 8316
rect 4120 8344 4126 8356
rect 4540 8344 4568 8579
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 7800 8588 8493 8616
rect 7800 8576 7806 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9674 8616 9680 8628
rect 9539 8588 9680 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 6641 8551 6699 8557
rect 6641 8517 6653 8551
rect 6687 8548 6699 8551
rect 6822 8548 6828 8560
rect 6687 8520 6828 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 6822 8508 6828 8520
rect 6880 8548 6886 8560
rect 8202 8548 8208 8560
rect 6880 8520 8208 8548
rect 6880 8508 6886 8520
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 8496 8548 8524 8579
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8616 9827 8619
rect 10042 8616 10048 8628
rect 9815 8588 10048 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 10042 8576 10048 8588
rect 10100 8616 10106 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 10100 8588 12173 8616
rect 10100 8576 10106 8588
rect 12161 8585 12173 8588
rect 12207 8616 12219 8619
rect 12894 8616 12900 8628
rect 12207 8588 12900 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 12894 8576 12900 8588
rect 12952 8616 12958 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 12952 8588 13645 8616
rect 12952 8576 12958 8588
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 15562 8616 15568 8628
rect 15523 8588 15568 8616
rect 13633 8579 13691 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 25130 8616 25136 8628
rect 25091 8588 25136 8616
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 9858 8548 9864 8560
rect 8496 8520 9864 8548
rect 9858 8508 9864 8520
rect 9916 8548 9922 8560
rect 10502 8548 10508 8560
rect 9916 8520 10508 8548
rect 9916 8508 9922 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 5500 8452 7205 8480
rect 5500 8440 5506 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7926 8480 7932 8492
rect 7887 8452 7932 8480
rect 7193 8443 7251 8449
rect 7926 8440 7932 8452
rect 7984 8440 7990 8492
rect 9950 8480 9956 8492
rect 9911 8452 9956 8480
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 12434 8480 12440 8492
rect 12395 8452 12440 8480
rect 12434 8440 12440 8452
rect 12492 8440 12498 8492
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 14366 8480 14372 8492
rect 13780 8452 14372 8480
rect 13780 8440 13786 8452
rect 14366 8440 14372 8452
rect 14424 8480 14430 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14424 8452 14565 8480
rect 14424 8440 14430 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 16114 8480 16120 8492
rect 16075 8452 16120 8480
rect 14553 8443 14611 8449
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 4982 8412 4988 8424
rect 4943 8384 4988 8412
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 7892 8384 8401 8412
rect 7892 8372 7898 8384
rect 8389 8381 8401 8384
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 8941 8415 8999 8421
rect 8941 8381 8953 8415
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 24648 8415 24706 8421
rect 13403 8384 13814 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 4120 8316 4568 8344
rect 4120 8304 4126 8316
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5592 8316 6684 8344
rect 5592 8304 5598 8316
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 5353 8279 5411 8285
rect 5353 8276 5365 8279
rect 5316 8248 5365 8276
rect 5316 8236 5322 8248
rect 5353 8245 5365 8248
rect 5399 8245 5411 8279
rect 5902 8276 5908 8288
rect 5863 8248 5908 8276
rect 5353 8239 5411 8245
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 6270 8276 6276 8288
rect 6231 8248 6276 8276
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 6656 8276 6684 8316
rect 6730 8304 6736 8356
rect 6788 8344 6794 8356
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 6788 8316 6929 8344
rect 6788 8304 6794 8316
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 6917 8307 6975 8313
rect 7009 8347 7067 8353
rect 7009 8313 7021 8347
rect 7055 8313 7067 8347
rect 7009 8307 7067 8313
rect 7024 8276 7052 8307
rect 7282 8276 7288 8288
rect 6656 8248 7288 8276
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 8202 8276 8208 8288
rect 8163 8248 8208 8276
rect 8202 8236 8208 8248
rect 8260 8276 8266 8288
rect 8956 8276 8984 8375
rect 10042 8304 10048 8356
rect 10100 8344 10106 8356
rect 10274 8347 10332 8353
rect 10274 8344 10286 8347
rect 10100 8316 10286 8344
rect 10100 8304 10106 8316
rect 10274 8313 10286 8316
rect 10320 8313 10332 8347
rect 10274 8307 10332 8313
rect 12799 8347 12857 8353
rect 12799 8313 12811 8347
rect 12845 8344 12857 8347
rect 12894 8344 12900 8356
rect 12845 8316 12900 8344
rect 12845 8313 12857 8316
rect 12799 8307 12857 8313
rect 12894 8304 12900 8316
rect 12952 8304 12958 8356
rect 8260 8248 8984 8276
rect 8260 8236 8266 8248
rect 10686 8236 10692 8288
rect 10744 8276 10750 8288
rect 10873 8279 10931 8285
rect 10873 8276 10885 8279
rect 10744 8248 10885 8276
rect 10744 8236 10750 8248
rect 10873 8245 10885 8248
rect 10919 8276 10931 8279
rect 11149 8279 11207 8285
rect 11149 8276 11161 8279
rect 10919 8248 11161 8276
rect 10919 8245 10931 8248
rect 10873 8239 10931 8245
rect 11149 8245 11161 8248
rect 11195 8276 11207 8279
rect 11330 8276 11336 8288
rect 11195 8248 11336 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11606 8276 11612 8288
rect 11567 8248 11612 8276
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 13786 8276 13814 8384
rect 24648 8381 24660 8415
rect 24694 8412 24706 8415
rect 25130 8412 25136 8424
rect 24694 8384 25136 8412
rect 24694 8381 24706 8384
rect 24648 8375 24706 8381
rect 25130 8372 25136 8384
rect 25188 8372 25194 8424
rect 14274 8344 14280 8356
rect 14235 8316 14280 8344
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 15289 8347 15347 8353
rect 15289 8313 15301 8347
rect 15335 8344 15347 8347
rect 15838 8344 15844 8356
rect 15335 8316 15844 8344
rect 15335 8313 15347 8316
rect 15289 8307 15347 8313
rect 14090 8276 14096 8288
rect 13786 8248 14096 8276
rect 14090 8236 14096 8248
rect 14148 8276 14154 8288
rect 14384 8276 14412 8307
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 15933 8347 15991 8353
rect 15933 8313 15945 8347
rect 15979 8313 15991 8347
rect 15933 8307 15991 8313
rect 14148 8248 14412 8276
rect 14148 8236 14154 8248
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 15948 8276 15976 8307
rect 15620 8248 15976 8276
rect 15620 8236 15626 8248
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 24719 8279 24777 8285
rect 24719 8276 24731 8279
rect 18656 8248 24731 8276
rect 18656 8236 18662 8248
rect 24719 8245 24731 8248
rect 24765 8245 24777 8279
rect 24719 8239 24777 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 2096 8044 2605 8072
rect 2096 8032 2102 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 4614 8072 4620 8084
rect 4575 8044 4620 8072
rect 2593 8035 2651 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5721 8075 5779 8081
rect 5721 8072 5733 8075
rect 5040 8044 5733 8072
rect 5040 8032 5046 8044
rect 5721 8041 5733 8044
rect 5767 8041 5779 8075
rect 7282 8072 7288 8084
rect 7243 8044 7288 8072
rect 5721 8035 5779 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9950 8072 9956 8084
rect 9911 8044 9956 8072
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 13078 8072 13084 8084
rect 13039 8044 13084 8072
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8072 15163 8075
rect 15286 8072 15292 8084
rect 15151 8044 15292 8072
rect 15151 8041 15163 8044
rect 15105 8035 15163 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 15838 8032 15844 8084
rect 15896 8072 15902 8084
rect 16853 8075 16911 8081
rect 16853 8072 16865 8075
rect 15896 8044 16865 8072
rect 15896 8032 15902 8044
rect 16853 8041 16865 8044
rect 16899 8041 16911 8075
rect 16853 8035 16911 8041
rect 1762 8004 1768 8016
rect 1723 7976 1768 8004
rect 1762 7964 1768 7976
rect 1820 7964 1826 8016
rect 4798 7964 4804 8016
rect 4856 8004 4862 8016
rect 4893 8007 4951 8013
rect 4893 8004 4905 8007
rect 4856 7976 4905 8004
rect 4856 7964 4862 7976
rect 4893 7973 4905 7976
rect 4939 7973 4951 8007
rect 5442 8004 5448 8016
rect 5403 7976 5448 8004
rect 4893 7967 4951 7973
rect 5442 7964 5448 7976
rect 5500 7964 5506 8016
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 6362 8004 6368 8016
rect 5960 7976 6368 8004
rect 5960 7964 5966 7976
rect 6362 7964 6368 7976
rect 6420 8004 6426 8016
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 6420 7976 6469 8004
rect 6420 7964 6426 7976
rect 6457 7973 6469 7976
rect 6503 7973 6515 8007
rect 6457 7967 6515 7973
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 10642 8007 10700 8013
rect 10642 8004 10654 8007
rect 10100 7976 10654 8004
rect 10100 7964 10106 7976
rect 10642 7973 10654 7976
rect 10688 7973 10700 8007
rect 12250 8004 12256 8016
rect 10642 7967 10700 7973
rect 11256 7976 12256 8004
rect 8481 7939 8539 7945
rect 8481 7905 8493 7939
rect 8527 7936 8539 7939
rect 8570 7936 8576 7948
rect 8527 7908 8576 7936
rect 8527 7905 8539 7908
rect 8481 7899 8539 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 9824 7908 10333 7936
rect 9824 7896 9830 7908
rect 10321 7905 10333 7908
rect 10367 7936 10379 7939
rect 10962 7936 10968 7948
rect 10367 7908 10968 7936
rect 10367 7905 10379 7908
rect 10321 7899 10379 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11256 7945 11284 7976
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 13814 7964 13820 8016
rect 13872 8004 13878 8016
rect 14366 8004 14372 8016
rect 13872 7976 13917 8004
rect 14327 7976 14372 8004
rect 13872 7964 13878 7976
rect 14366 7964 14372 7976
rect 14424 7964 14430 8016
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 15473 8007 15531 8013
rect 15473 8004 15485 8007
rect 15436 7976 15485 8004
rect 15436 7964 15442 7976
rect 15473 7973 15485 7976
rect 15519 8004 15531 8007
rect 16206 8004 16212 8016
rect 15519 7976 16212 8004
rect 15519 7973 15531 7976
rect 15473 7967 15531 7973
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7905 11299 7939
rect 11241 7899 11299 7905
rect 24648 7939 24706 7945
rect 24648 7905 24660 7939
rect 24694 7936 24706 7939
rect 25498 7936 25504 7948
rect 24694 7908 25504 7936
rect 24694 7905 24706 7908
rect 24648 7899 24706 7905
rect 25498 7896 25504 7908
rect 25556 7896 25562 7948
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1673 7831 1731 7837
rect 1578 7760 1584 7812
rect 1636 7800 1642 7812
rect 1688 7800 1716 7831
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 5074 7868 5080 7880
rect 4847 7840 5080 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 6454 7868 6460 7880
rect 6411 7840 6460 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 6730 7868 6736 7880
rect 6691 7840 6736 7868
rect 6730 7828 6736 7840
rect 6788 7868 6794 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 6788 7840 7665 7868
rect 6788 7828 6794 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7834 7868 7840 7880
rect 7795 7840 7840 7868
rect 7653 7831 7711 7837
rect 7834 7828 7840 7840
rect 7892 7868 7898 7880
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 7892 7840 9229 7868
rect 7892 7828 7898 7840
rect 9217 7837 9229 7840
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11940 7840 12173 7868
rect 11940 7828 11946 7840
rect 12161 7837 12173 7840
rect 12207 7868 12219 7871
rect 12618 7868 12624 7880
rect 12207 7840 12624 7868
rect 12207 7837 12219 7840
rect 12161 7831 12219 7837
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7837 15439 7871
rect 15654 7868 15660 7880
rect 15615 7840 15660 7868
rect 15381 7831 15439 7837
rect 1636 7772 1716 7800
rect 1636 7760 1642 7772
rect 1688 7732 1716 7772
rect 1854 7760 1860 7812
rect 1912 7800 1918 7812
rect 2590 7800 2596 7812
rect 1912 7772 2596 7800
rect 1912 7760 1918 7772
rect 2590 7760 2596 7772
rect 2648 7800 2654 7812
rect 2961 7803 3019 7809
rect 2961 7800 2973 7803
rect 2648 7772 2973 7800
rect 2648 7760 2654 7772
rect 2961 7769 2973 7772
rect 3007 7769 3019 7803
rect 2961 7763 3019 7769
rect 3694 7760 3700 7812
rect 3752 7800 3758 7812
rect 5442 7800 5448 7812
rect 3752 7772 5448 7800
rect 3752 7760 3758 7772
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 3329 7735 3387 7741
rect 3329 7732 3341 7735
rect 1688 7704 3341 7732
rect 3329 7701 3341 7704
rect 3375 7701 3387 7735
rect 15396 7732 15424 7831
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 16206 7732 16212 7744
rect 15396 7704 16212 7732
rect 3329 7695 3387 7701
rect 16206 7692 16212 7704
rect 16264 7732 16270 7744
rect 24719 7735 24777 7741
rect 24719 7732 24731 7735
rect 16264 7704 24731 7732
rect 16264 7692 16270 7704
rect 24719 7701 24731 7704
rect 24765 7701 24777 7735
rect 24719 7695 24777 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 3142 7528 3148 7540
rect 2823 7500 3148 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 6086 7528 6092 7540
rect 6047 7500 6092 7528
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 6362 7528 6368 7540
rect 6323 7500 6368 7528
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9180 7500 9597 7528
rect 9180 7488 9186 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9585 7491 9643 7497
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10100 7500 10333 7528
rect 10100 7488 10106 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 10870 7528 10876 7540
rect 10831 7500 10876 7528
rect 10321 7491 10379 7497
rect 6270 7420 6276 7472
rect 6328 7460 6334 7472
rect 7377 7463 7435 7469
rect 7377 7460 7389 7463
rect 6328 7432 7389 7460
rect 6328 7420 6334 7432
rect 7377 7429 7389 7432
rect 7423 7460 7435 7463
rect 8570 7460 8576 7472
rect 7423 7432 8576 7460
rect 7423 7429 7435 7432
rect 7377 7423 7435 7429
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 1854 7392 1860 7404
rect 1811 7364 1860 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 2004 7364 2053 7392
rect 2004 7352 2010 7364
rect 2041 7361 2053 7364
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 7190 7352 7196 7404
rect 7248 7392 7254 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 7248 7364 9873 7392
rect 7248 7352 7254 7364
rect 3142 7284 3148 7336
rect 3200 7324 3206 7336
rect 3329 7327 3387 7333
rect 3329 7324 3341 7327
rect 3200 7296 3341 7324
rect 3200 7284 3206 7296
rect 3329 7293 3341 7296
rect 3375 7293 3387 7327
rect 3329 7287 3387 7293
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7324 4491 7327
rect 4522 7324 4528 7336
rect 4479 7296 4528 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 4522 7284 4528 7296
rect 4580 7324 4586 7336
rect 4985 7327 5043 7333
rect 4985 7324 4997 7327
rect 4580 7296 4997 7324
rect 4580 7284 4586 7296
rect 4985 7293 4997 7296
rect 5031 7293 5043 7327
rect 4985 7287 5043 7293
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 6086 7324 6092 7336
rect 5583 7296 6092 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 7650 7284 7656 7336
rect 7708 7324 7714 7336
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7708 7296 7757 7324
rect 7708 7284 7714 7296
rect 7745 7293 7757 7296
rect 7791 7324 7803 7327
rect 7926 7324 7932 7336
rect 7791 7296 7932 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 9416 7333 9444 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 10336 7392 10364 7491
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12250 7528 12256 7540
rect 11931 7500 12256 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 15378 7528 15384 7540
rect 15339 7500 15384 7528
rect 15378 7488 15384 7500
rect 15436 7488 15442 7540
rect 16117 7531 16175 7537
rect 16117 7497 16129 7531
rect 16163 7528 16175 7531
rect 16206 7528 16212 7540
rect 16163 7500 16212 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 24719 7463 24777 7469
rect 24719 7429 24731 7463
rect 24765 7429 24777 7463
rect 24719 7423 24777 7429
rect 10870 7392 10876 7404
rect 10336 7364 10876 7392
rect 9861 7355 9919 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 12802 7392 12808 7404
rect 12763 7364 12808 7392
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 13814 7392 13820 7404
rect 13771 7364 13820 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 13814 7352 13820 7364
rect 13872 7392 13878 7404
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13872 7364 14013 7392
rect 13872 7352 13878 7364
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 14001 7355 14059 7361
rect 24118 7352 24124 7404
rect 24176 7392 24182 7404
rect 24734 7392 24762 7423
rect 24176 7364 24762 7392
rect 24176 7352 24182 7364
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 10686 7324 10692 7336
rect 10647 7296 10692 7324
rect 9401 7287 9459 7293
rect 10686 7284 10692 7296
rect 10744 7284 10750 7336
rect 14090 7324 14096 7336
rect 14051 7296 14096 7324
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 15632 7327 15690 7333
rect 15632 7293 15644 7327
rect 15678 7324 15690 7327
rect 16114 7324 16120 7336
rect 15678 7296 16120 7324
rect 15678 7293 15690 7296
rect 15632 7287 15690 7293
rect 16114 7284 16120 7296
rect 16172 7324 16178 7336
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 16172 7296 16405 7324
rect 16172 7284 16178 7296
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 24648 7327 24706 7333
rect 24648 7293 24660 7327
rect 24694 7324 24706 7327
rect 25133 7327 25191 7333
rect 25133 7324 25145 7327
rect 24694 7296 25145 7324
rect 24694 7293 24706 7296
rect 24648 7287 24706 7293
rect 25133 7293 25145 7296
rect 25179 7324 25191 7327
rect 27614 7324 27620 7336
rect 25179 7296 27620 7324
rect 25179 7293 25191 7296
rect 25133 7287 25191 7293
rect 27614 7284 27620 7296
rect 27672 7284 27678 7336
rect 1857 7259 1915 7265
rect 1857 7225 1869 7259
rect 1903 7225 1915 7259
rect 1857 7219 1915 7225
rect 1872 7188 1900 7219
rect 3160 7188 3188 7284
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 8573 7259 8631 7265
rect 3292 7228 3337 7256
rect 3292 7216 3298 7228
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8662 7256 8668 7268
rect 8619 7228 8668 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 12526 7256 12532 7268
rect 12487 7228 12532 7256
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 12621 7259 12679 7265
rect 12621 7225 12633 7259
rect 12667 7225 12679 7259
rect 12621 7219 12679 7225
rect 4798 7188 4804 7200
rect 1872 7160 3188 7188
rect 4759 7160 4804 7188
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 5040 7160 5089 7188
rect 5040 7148 5046 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 5077 7151 5135 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 12158 7188 12164 7200
rect 12119 7160 12164 7188
rect 12158 7148 12164 7160
rect 12216 7188 12222 7200
rect 12636 7188 12664 7219
rect 12216 7160 12664 7188
rect 15703 7191 15761 7197
rect 12216 7148 12222 7160
rect 15703 7157 15715 7191
rect 15749 7188 15761 7191
rect 15838 7188 15844 7200
rect 15749 7160 15844 7188
rect 15749 7157 15761 7160
rect 15703 7151 15761 7157
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 25498 7188 25504 7200
rect 25411 7160 25504 7188
rect 25498 7148 25504 7160
rect 25556 7188 25562 7200
rect 26510 7188 26516 7200
rect 25556 7160 26516 7188
rect 25556 7148 25562 7160
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 1820 6956 2145 6984
rect 1820 6944 1826 6956
rect 2133 6953 2145 6956
rect 2179 6984 2191 6987
rect 3234 6984 3240 6996
rect 2179 6956 3240 6984
rect 2179 6953 2191 6956
rect 2133 6947 2191 6953
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 4801 6987 4859 6993
rect 4801 6953 4813 6987
rect 4847 6984 4859 6987
rect 5074 6984 5080 6996
rect 4847 6956 5080 6984
rect 4847 6953 4859 6956
rect 4801 6947 4859 6953
rect 5074 6944 5080 6956
rect 5132 6984 5138 6996
rect 6822 6984 6828 6996
rect 5132 6956 6828 6984
rect 5132 6944 5138 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 8665 6987 8723 6993
rect 8665 6984 8677 6987
rect 8168 6956 8677 6984
rect 8168 6944 8174 6956
rect 8665 6953 8677 6956
rect 8711 6984 8723 6987
rect 9674 6984 9680 6996
rect 8711 6956 9680 6984
rect 8711 6953 8723 6956
rect 8665 6947 8723 6953
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9861 6987 9919 6993
rect 9861 6984 9873 6987
rect 9784 6956 9873 6984
rect 2587 6919 2645 6925
rect 2587 6885 2599 6919
rect 2633 6916 2645 6919
rect 2958 6916 2964 6928
rect 2633 6888 2964 6916
rect 2633 6885 2645 6888
rect 2587 6879 2645 6885
rect 2958 6876 2964 6888
rect 3016 6876 3022 6928
rect 4890 6876 4896 6928
rect 4948 6916 4954 6928
rect 4985 6919 5043 6925
rect 4985 6916 4997 6919
rect 4948 6888 4997 6916
rect 4948 6876 4954 6888
rect 4985 6885 4997 6888
rect 5031 6885 5043 6919
rect 4985 6879 5043 6885
rect 5166 6876 5172 6928
rect 5224 6916 5230 6928
rect 8297 6919 8355 6925
rect 8297 6916 8309 6919
rect 5224 6888 8309 6916
rect 5224 6876 5230 6888
rect 8297 6885 8309 6888
rect 8343 6885 8355 6919
rect 8297 6879 8355 6885
rect 9582 6876 9588 6928
rect 9640 6916 9646 6928
rect 9784 6916 9812 6956
rect 9861 6953 9873 6956
rect 9907 6953 9919 6987
rect 10686 6984 10692 6996
rect 10647 6956 10692 6984
rect 9861 6947 9919 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 10962 6984 10968 6996
rect 10923 6956 10968 6984
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 12526 6984 12532 6996
rect 12487 6956 12532 6984
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12676 6956 12817 6984
rect 12676 6944 12682 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 14090 6984 14096 6996
rect 14051 6956 14096 6984
rect 12805 6947 12863 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 12158 6916 12164 6928
rect 9640 6888 9812 6916
rect 12119 6888 12164 6916
rect 9640 6876 9646 6888
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2314 6848 2320 6860
rect 2271 6820 2320 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6848 5687 6851
rect 6362 6848 6368 6860
rect 5675 6820 6368 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 6638 6848 6644 6860
rect 6595 6820 6644 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 6788 6820 7573 6848
rect 6788 6808 6794 6820
rect 7561 6817 7573 6820
rect 7607 6817 7619 6851
rect 7561 6811 7619 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9766 6848 9772 6860
rect 9723 6820 9772 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 12069 6851 12127 6857
rect 12069 6817 12081 6851
rect 12115 6848 12127 6851
rect 12250 6848 12256 6860
rect 12115 6820 12256 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12802 6808 12808 6860
rect 12860 6848 12866 6860
rect 13024 6851 13082 6857
rect 13024 6848 13036 6851
rect 12860 6820 13036 6848
rect 12860 6808 12866 6820
rect 13024 6817 13036 6820
rect 13070 6817 13082 6851
rect 15838 6848 15844 6860
rect 15799 6820 15844 6848
rect 13024 6811 13082 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17034 6848 17040 6860
rect 16991 6820 17040 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7708 6783 7766 6789
rect 7708 6780 7720 6783
rect 7248 6752 7720 6780
rect 7248 6740 7254 6752
rect 7708 6749 7720 6752
rect 7754 6749 7766 6783
rect 7708 6743 7766 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8478 6780 8484 6792
rect 7975 6752 8484 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 13633 6783 13691 6789
rect 13633 6780 13645 6783
rect 13320 6752 13645 6780
rect 13320 6740 13326 6752
rect 13633 6749 13645 6752
rect 13679 6780 13691 6783
rect 13722 6780 13728 6792
rect 13679 6752 13728 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 6365 6715 6423 6721
rect 6365 6681 6377 6715
rect 6411 6712 6423 6715
rect 6454 6712 6460 6724
rect 6411 6684 6460 6712
rect 6411 6681 6423 6684
rect 6365 6675 6423 6681
rect 6454 6672 6460 6684
rect 6512 6712 6518 6724
rect 17083 6715 17141 6721
rect 17083 6712 17095 6715
rect 6512 6684 17095 6712
rect 6512 6672 6518 6684
rect 17083 6681 17095 6684
rect 17129 6681 17141 6715
rect 17083 6675 17141 6681
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 1854 6644 1860 6656
rect 1811 6616 1860 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 3142 6644 3148 6656
rect 3103 6616 3148 6644
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 6730 6644 6736 6656
rect 5408 6616 6736 6644
rect 5408 6604 5414 6616
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 7742 6644 7748 6656
rect 7515 6616 7748 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 7837 6647 7895 6653
rect 7837 6613 7849 6647
rect 7883 6644 7895 6647
rect 8018 6644 8024 6656
rect 7883 6616 8024 6644
rect 7883 6613 7895 6616
rect 7837 6607 7895 6613
rect 8018 6604 8024 6616
rect 8076 6644 8082 6656
rect 9214 6644 9220 6656
rect 8076 6616 9220 6644
rect 8076 6604 8082 6616
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 13127 6647 13185 6653
rect 13127 6613 13139 6647
rect 13173 6644 13185 6647
rect 13446 6644 13452 6656
rect 13173 6616 13452 6644
rect 13173 6613 13185 6616
rect 13127 6607 13185 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 16025 6647 16083 6653
rect 16025 6613 16037 6647
rect 16071 6644 16083 6647
rect 16666 6644 16672 6656
rect 16071 6616 16672 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 6362 6440 6368 6452
rect 5951 6412 6368 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 7248 6412 7665 6440
rect 7248 6400 7254 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 7742 6400 7748 6452
rect 7800 6440 7806 6452
rect 7975 6443 8033 6449
rect 7975 6440 7987 6443
rect 7800 6412 7987 6440
rect 7800 6400 7806 6412
rect 7975 6409 7987 6412
rect 8021 6409 8033 6443
rect 8110 6440 8116 6452
rect 8071 6412 8116 6440
rect 7975 6403 8033 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8481 6443 8539 6449
rect 8481 6409 8493 6443
rect 8527 6440 8539 6443
rect 11146 6440 11152 6452
rect 8527 6412 11152 6440
rect 8527 6409 8539 6412
rect 8481 6403 8539 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 12250 6440 12256 6452
rect 11563 6412 12256 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12802 6400 12808 6452
rect 12860 6440 12866 6452
rect 12989 6443 13047 6449
rect 12989 6440 13001 6443
rect 12860 6412 13001 6440
rect 12860 6400 12866 6412
rect 12989 6409 13001 6412
rect 13035 6409 13047 6443
rect 15838 6440 15844 6452
rect 15799 6412 15844 6440
rect 12989 6403 13047 6409
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 9214 6372 9220 6384
rect 9175 6344 9220 6372
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 20993 6375 21051 6381
rect 20993 6341 21005 6375
rect 21039 6372 21051 6375
rect 22922 6372 22928 6384
rect 21039 6344 22928 6372
rect 21039 6341 21051 6344
rect 20993 6335 21051 6341
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 2130 6304 2136 6316
rect 2091 6276 2136 6304
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 2222 6264 2228 6316
rect 2280 6304 2286 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2280 6276 3065 6304
rect 2280 6264 2286 6276
rect 3053 6273 3065 6276
rect 3099 6304 3111 6307
rect 3142 6304 3148 6316
rect 3099 6276 3148 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3142 6264 3148 6276
rect 3200 6304 3206 6316
rect 4798 6304 4804 6316
rect 3200 6276 3372 6304
rect 4759 6276 4804 6304
rect 3200 6264 3206 6276
rect 3344 6245 3372 6276
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6788 6276 7205 6304
rect 6788 6264 6794 6276
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8662 6304 8668 6316
rect 8251 6276 8668 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12526 6304 12532 6316
rect 12483 6276 12532 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12526 6264 12532 6276
rect 12584 6264 12590 6316
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6205 3387 6239
rect 3329 6199 3387 6205
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4755 6208 4905 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4893 6205 4905 6208
rect 4939 6236 4951 6239
rect 5534 6236 5540 6248
rect 4939 6208 5540 6236
rect 4939 6205 4951 6208
rect 4893 6199 4951 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 20806 6236 20812 6248
rect 20767 6208 20812 6236
rect 20806 6196 20812 6208
rect 20864 6236 20870 6248
rect 21361 6239 21419 6245
rect 21361 6236 21373 6239
rect 20864 6208 21373 6236
rect 20864 6196 20870 6208
rect 21361 6205 21373 6208
rect 21407 6205 21419 6239
rect 21361 6199 21419 6205
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 3237 6171 3295 6177
rect 3237 6168 3249 6171
rect 1912 6140 2005 6168
rect 2602 6140 3249 6168
rect 1912 6128 1918 6140
rect 1872 6100 1900 6128
rect 2602 6100 2630 6140
rect 3237 6137 3249 6140
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 7650 6128 7656 6180
rect 7708 6168 7714 6180
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7708 6140 7849 6168
rect 7708 6128 7714 6140
rect 7837 6137 7849 6140
rect 7883 6168 7895 6171
rect 8386 6168 8392 6180
rect 7883 6140 8392 6168
rect 7883 6137 7895 6140
rect 7837 6131 7895 6137
rect 8386 6128 8392 6140
rect 8444 6168 8450 6180
rect 8849 6171 8907 6177
rect 8849 6168 8861 6171
rect 8444 6140 8861 6168
rect 8444 6128 8450 6140
rect 8849 6137 8861 6140
rect 8895 6137 8907 6171
rect 8849 6131 8907 6137
rect 1872 6072 2630 6100
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 2958 6100 2964 6112
rect 2823 6072 2964 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 6638 6100 6644 6112
rect 6599 6072 6644 6100
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 17034 6100 17040 6112
rect 16947 6072 17040 6100
rect 17034 6060 17040 6072
rect 17092 6100 17098 6112
rect 18598 6100 18604 6112
rect 17092 6072 18604 6100
rect 17092 6060 17098 6072
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 1820 5868 3065 5896
rect 1820 5856 1826 5868
rect 3053 5865 3065 5868
rect 3099 5896 3111 5899
rect 4203 5899 4261 5905
rect 4203 5896 4215 5899
rect 3099 5868 4215 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 4203 5865 4215 5868
rect 4249 5865 4261 5899
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 4203 5859 4261 5865
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8662 5896 8668 5908
rect 8623 5868 8668 5896
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 2222 5828 2228 5840
rect 1903 5800 2228 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 2685 5831 2743 5837
rect 2685 5828 2697 5831
rect 2464 5800 2697 5828
rect 2464 5788 2470 5800
rect 2685 5797 2697 5800
rect 2731 5797 2743 5831
rect 2685 5791 2743 5797
rect 7561 5831 7619 5837
rect 7561 5797 7573 5831
rect 7607 5828 7619 5831
rect 8478 5828 8484 5840
rect 7607 5800 8484 5828
rect 7607 5797 7619 5800
rect 7561 5791 7619 5797
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 3973 5763 4031 5769
rect 3973 5729 3985 5763
rect 4019 5760 4031 5763
rect 4062 5760 4068 5772
rect 4019 5732 4068 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 7248 5732 7665 5760
rect 7248 5720 7254 5732
rect 7653 5729 7665 5732
rect 7699 5760 7711 5763
rect 7834 5760 7840 5772
rect 7699 5732 7840 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 7818 5627 7876 5633
rect 7818 5593 7830 5627
rect 7864 5624 7876 5627
rect 8294 5624 8300 5636
rect 7864 5596 8300 5624
rect 7864 5593 7876 5596
rect 7818 5587 7876 5593
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 7926 5556 7932 5568
rect 7616 5528 7932 5556
rect 7616 5516 7622 5528
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 3050 5352 3056 5364
rect 3011 5324 3056 5352
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 6696 5324 8769 5352
rect 6696 5312 6702 5324
rect 8757 5321 8769 5324
rect 8803 5352 8815 5355
rect 10134 5352 10140 5364
rect 8803 5324 10140 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 4062 5284 4068 5296
rect 4023 5256 4068 5284
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 8018 5244 8024 5296
rect 8076 5284 8082 5296
rect 8389 5287 8447 5293
rect 8389 5284 8401 5287
rect 8076 5256 8401 5284
rect 8076 5244 8082 5256
rect 8389 5253 8401 5256
rect 8435 5284 8447 5287
rect 9766 5284 9772 5296
rect 8435 5256 9772 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 1535 5219 1593 5225
rect 1535 5185 1547 5219
rect 1581 5216 1593 5219
rect 3050 5216 3056 5228
rect 1581 5188 3056 5216
rect 1581 5185 1593 5188
rect 1535 5179 1593 5185
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 1448 5151 1506 5157
rect 1448 5117 1460 5151
rect 1494 5148 1506 5151
rect 1670 5148 1676 5160
rect 1494 5120 1676 5148
rect 1494 5117 1506 5120
rect 1448 5111 1506 5117
rect 1670 5108 1676 5120
rect 1728 5148 1734 5160
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1728 5120 1869 5148
rect 1728 5108 1734 5120
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2731 5120 2881 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 2869 5117 2881 5120
rect 2915 5148 2927 5151
rect 3786 5148 3792 5160
rect 2915 5120 3792 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 7009 5151 7067 5157
rect 7009 5117 7021 5151
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 8665 5151 8723 5157
rect 8665 5117 8677 5151
rect 8711 5148 8723 5151
rect 8711 5120 9444 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 1210 5040 1216 5092
rect 1268 5080 1274 5092
rect 6549 5083 6607 5089
rect 6549 5080 6561 5083
rect 1268 5052 6561 5080
rect 1268 5040 1274 5052
rect 6549 5049 6561 5052
rect 6595 5080 6607 5083
rect 7024 5080 7052 5111
rect 7282 5080 7288 5092
rect 6595 5052 7288 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 7282 5040 7288 5052
rect 7340 5040 7346 5092
rect 7653 5083 7711 5089
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 8478 5080 8484 5092
rect 7699 5052 8484 5080
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 9416 5024 9444 5120
rect 5166 4972 5172 5024
rect 5224 5012 5230 5024
rect 7926 5012 7932 5024
rect 5224 4984 7932 5012
rect 5224 4972 5230 4984
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 9398 5012 9404 5024
rect 9359 4984 9404 5012
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1857 4811 1915 4817
rect 1857 4808 1869 4811
rect 1820 4780 1869 4808
rect 1820 4768 1826 4780
rect 1857 4777 1869 4780
rect 1903 4777 1915 4811
rect 2590 4808 2596 4820
rect 2551 4780 2596 4808
rect 1857 4771 1915 4777
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 7190 4808 7196 4820
rect 7151 4780 7196 4808
rect 7190 4768 7196 4780
rect 7248 4768 7254 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 8665 4811 8723 4817
rect 8665 4808 8677 4811
rect 8536 4780 8677 4808
rect 8536 4768 8542 4780
rect 8665 4777 8677 4780
rect 8711 4777 8723 4811
rect 8665 4771 8723 4777
rect 1535 4743 1593 4749
rect 1535 4709 1547 4743
rect 1581 4740 1593 4743
rect 10778 4740 10784 4752
rect 1581 4712 10784 4740
rect 1581 4709 1593 4712
rect 1535 4703 1593 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 2406 4672 2412 4684
rect 2367 4644 2412 4672
rect 2406 4632 2412 4644
rect 2464 4632 2470 4684
rect 7282 4672 7288 4684
rect 7243 4644 7288 4672
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7466 4632 7472 4684
rect 7524 4672 7530 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7524 4644 8033 4672
rect 7524 4632 7530 4644
rect 8021 4641 8033 4644
rect 8067 4672 8079 4675
rect 9398 4672 9404 4684
rect 8067 4644 9404 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 7650 4604 7656 4616
rect 7611 4576 7656 4604
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8294 4468 8300 4480
rect 8255 4440 8300 4468
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 106 4224 112 4276
rect 164 4264 170 4276
rect 2406 4264 2412 4276
rect 164 4236 2412 4264
rect 164 4224 170 4236
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 7653 4267 7711 4273
rect 7653 4264 7665 4267
rect 7432 4236 7665 4264
rect 7432 4224 7438 4236
rect 7653 4233 7665 4236
rect 7699 4233 7711 4267
rect 7653 4227 7711 4233
rect 1535 4199 1593 4205
rect 1535 4165 1547 4199
rect 1581 4196 1593 4199
rect 1670 4196 1676 4208
rect 1581 4168 1676 4196
rect 1581 4165 1593 4168
rect 1535 4159 1593 4165
rect 1670 4156 1676 4168
rect 1728 4156 1734 4208
rect 7285 4199 7343 4205
rect 7285 4165 7297 4199
rect 7331 4196 7343 4199
rect 7466 4196 7472 4208
rect 7331 4168 7472 4196
rect 7331 4165 7343 4168
rect 7285 4159 7343 4165
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10686 4128 10692 4140
rect 10643 4100 10692 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 10686 4088 10692 4100
rect 10744 4128 10750 4140
rect 12342 4128 12348 4140
rect 10744 4100 12348 4128
rect 10744 4088 10750 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 1302 4020 1308 4072
rect 1360 4060 1366 4072
rect 1432 4063 1490 4069
rect 1432 4060 1444 4063
rect 1360 4032 1444 4060
rect 1360 4020 1366 4032
rect 1432 4029 1444 4032
rect 1478 4060 1490 4063
rect 1857 4063 1915 4069
rect 1857 4060 1869 4063
rect 1478 4032 1869 4060
rect 1478 4029 1490 4032
rect 1432 4023 1490 4029
rect 1857 4029 1869 4032
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 10505 3995 10563 4001
rect 10505 3961 10517 3995
rect 10551 3992 10563 3995
rect 10778 3992 10784 4004
rect 10551 3964 10784 3992
rect 10551 3961 10563 3964
rect 10505 3955 10563 3961
rect 10778 3952 10784 3964
rect 10836 3992 10842 4004
rect 10918 3995 10976 4001
rect 10918 3992 10930 3995
rect 10836 3964 10930 3992
rect 10836 3952 10842 3964
rect 10918 3961 10930 3964
rect 10964 3961 10976 3995
rect 10918 3955 10976 3961
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11480 3896 11529 3924
rect 11480 3884 11486 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1486 3680 1492 3732
rect 1544 3720 1550 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 1544 3692 1593 3720
rect 1544 3680 1550 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 10686 3720 10692 3732
rect 10647 3692 10692 3720
rect 1581 3683 1639 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11532 3692 13492 3720
rect 11422 3612 11428 3664
rect 11480 3652 11486 3664
rect 11532 3661 11560 3692
rect 11517 3655 11575 3661
rect 11517 3652 11529 3655
rect 11480 3624 11529 3652
rect 11480 3612 11486 3624
rect 11517 3621 11529 3624
rect 11563 3621 11575 3655
rect 11517 3615 11575 3621
rect 12069 3655 12127 3661
rect 12069 3621 12081 3655
rect 12115 3652 12127 3655
rect 13354 3652 13360 3664
rect 12115 3624 13360 3652
rect 12115 3621 12127 3624
rect 12069 3615 12127 3621
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 13464 3596 13492 3692
rect 13446 3584 13452 3596
rect 13407 3556 13452 3584
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 11514 3516 11520 3528
rect 11471 3488 11520 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 12894 3516 12900 3528
rect 12855 3488 12900 3516
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 12526 3380 12532 3392
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1535 3179 1593 3185
rect 1535 3145 1547 3179
rect 1581 3176 1593 3179
rect 3418 3176 3424 3188
rect 1581 3148 3424 3176
rect 1581 3145 1593 3148
rect 1535 3139 1593 3145
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 10367 3179 10425 3185
rect 10367 3145 10379 3179
rect 10413 3176 10425 3179
rect 10870 3176 10876 3188
rect 10413 3148 10876 3176
rect 10413 3145 10425 3148
rect 10367 3139 10425 3145
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 12526 3040 12532 3052
rect 12487 3012 12532 3040
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3040 13231 3043
rect 13354 3040 13360 3052
rect 13219 3012 13360 3040
rect 13219 3009 13231 3012
rect 13173 3003 13231 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 106 2932 112 2984
rect 164 2972 170 2984
rect 1432 2975 1490 2981
rect 1432 2972 1444 2975
rect 164 2944 1444 2972
rect 164 2932 170 2944
rect 1432 2941 1444 2944
rect 1478 2972 1490 2975
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1478 2944 1869 2972
rect 1478 2941 1490 2944
rect 1432 2935 1490 2941
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 10296 2975 10354 2981
rect 10296 2941 10308 2975
rect 10342 2972 10354 2975
rect 14068 2975 14126 2981
rect 10342 2944 10824 2972
rect 10342 2941 10354 2944
rect 10296 2935 10354 2941
rect 10796 2848 10824 2944
rect 14068 2941 14080 2975
rect 14114 2972 14126 2975
rect 14458 2972 14464 2984
rect 14114 2944 14464 2972
rect 14114 2941 14126 2944
rect 14068 2935 14126 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 12894 2904 12900 2916
rect 12667 2876 12900 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 10778 2836 10784 2848
rect 10739 2808 10784 2836
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 11701 2839 11759 2845
rect 11701 2836 11713 2839
rect 11572 2808 11713 2836
rect 11572 2796 11578 2808
rect 11701 2805 11713 2808
rect 11747 2805 11759 2839
rect 11701 2799 11759 2805
rect 12253 2839 12311 2845
rect 12253 2805 12265 2839
rect 12299 2836 12311 2839
rect 12636 2836 12664 2867
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 12299 2808 12664 2836
rect 12299 2805 12311 2808
rect 12253 2799 12311 2805
rect 13998 2796 14004 2848
rect 14056 2836 14062 2848
rect 14139 2839 14197 2845
rect 14139 2836 14151 2839
rect 14056 2808 14151 2836
rect 14056 2796 14062 2808
rect 14139 2805 14151 2808
rect 14185 2805 14197 2839
rect 14139 2799 14197 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 1762 2632 1768 2644
rect 1581 2604 1768 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 1762 2592 1768 2604
rect 1820 2592 1826 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5859 2635 5917 2641
rect 5859 2632 5871 2635
rect 4764 2604 5871 2632
rect 4764 2592 4770 2604
rect 5859 2601 5871 2604
rect 5905 2601 5917 2635
rect 5859 2595 5917 2601
rect 9907 2635 9965 2641
rect 9907 2601 9919 2635
rect 9953 2632 9965 2635
rect 11514 2632 11520 2644
rect 9953 2604 11520 2632
rect 9953 2601 9965 2604
rect 9907 2595 9965 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 11655 2635 11713 2641
rect 11655 2601 11667 2635
rect 11701 2632 11713 2635
rect 12526 2632 12532 2644
rect 11701 2604 12532 2632
rect 11701 2601 11713 2604
rect 11655 2595 11713 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2465 1522 2499
rect 1464 2459 1522 2465
rect 5788 2499 5846 2505
rect 5788 2465 5800 2499
rect 5834 2496 5846 2499
rect 5834 2468 6316 2496
rect 5834 2465 5846 2468
rect 5788 2459 5846 2465
rect 750 2388 756 2440
rect 808 2428 814 2440
rect 1479 2428 1507 2459
rect 1857 2431 1915 2437
rect 1857 2428 1869 2431
rect 808 2400 1869 2428
rect 808 2388 814 2400
rect 1857 2397 1869 2400
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 6288 2301 6316 2468
rect 9122 2456 9128 2508
rect 9180 2496 9186 2508
rect 9804 2499 9862 2505
rect 9804 2496 9816 2499
rect 9180 2468 9816 2496
rect 9180 2456 9186 2468
rect 9804 2465 9816 2468
rect 9850 2496 9862 2499
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9850 2468 10241 2496
rect 9850 2465 9862 2468
rect 9804 2459 9862 2465
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 11584 2499 11642 2505
rect 11584 2465 11596 2499
rect 11630 2496 11642 2499
rect 11630 2468 12112 2496
rect 11630 2465 11642 2468
rect 11584 2459 11642 2465
rect 6273 2295 6331 2301
rect 6273 2261 6285 2295
rect 6319 2292 6331 2295
rect 6638 2292 6644 2304
rect 6319 2264 6644 2292
rect 6319 2261 6331 2264
rect 6273 2255 6331 2261
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 12084 2301 12112 2468
rect 13998 2456 14004 2508
rect 14056 2496 14062 2508
rect 14093 2499 14151 2505
rect 14093 2496 14105 2499
rect 14056 2468 14105 2496
rect 14056 2456 14062 2468
rect 14093 2465 14105 2468
rect 14139 2496 14151 2499
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14139 2468 14657 2496
rect 14139 2465 14151 2468
rect 14093 2459 14151 2465
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 19036 2499 19094 2505
rect 19036 2465 19048 2499
rect 19082 2496 19094 2499
rect 19082 2468 19564 2496
rect 19082 2465 19094 2468
rect 19036 2459 19094 2465
rect 12069 2295 12127 2301
rect 12069 2261 12081 2295
rect 12115 2292 12127 2295
rect 12526 2292 12532 2304
rect 12115 2264 12532 2292
rect 12115 2261 12127 2264
rect 12069 2255 12127 2261
rect 12526 2252 12532 2264
rect 12584 2252 12590 2304
rect 14277 2295 14335 2301
rect 14277 2261 14289 2295
rect 14323 2292 14335 2295
rect 14550 2292 14556 2304
rect 14323 2264 14556 2292
rect 14323 2261 14335 2264
rect 14277 2255 14335 2261
rect 14550 2252 14556 2264
rect 14608 2252 14614 2304
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 19536 2301 19564 2468
rect 19107 2295 19165 2301
rect 19107 2292 19119 2295
rect 16080 2264 19119 2292
rect 16080 2252 16086 2264
rect 19107 2261 19119 2264
rect 19153 2261 19165 2295
rect 19107 2255 19165 2261
rect 19521 2295 19579 2301
rect 19521 2261 19533 2295
rect 19567 2292 19579 2295
rect 20622 2292 20628 2304
rect 19567 2264 20628 2292
rect 19567 2261 19579 2264
rect 19521 2255 19579 2261
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 23750 76 23756 128
rect 23808 116 23814 128
rect 24854 116 24860 128
rect 23808 88 24860 116
rect 23808 76 23814 88
rect 24854 76 24860 88
rect 24912 76 24918 128
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 10140 24148 10192 24200
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1308 23672 1360 23724
rect 6920 23808 6972 23860
rect 10876 23808 10928 23860
rect 1124 23468 1176 23520
rect 5448 23468 5500 23520
rect 11060 23604 11112 23656
rect 14832 23808 14884 23860
rect 16856 23808 16908 23860
rect 22836 23808 22888 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 19340 23604 19392 23656
rect 25136 23604 25188 23656
rect 21180 23536 21232 23588
rect 12532 23468 12584 23520
rect 14372 23468 14424 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 24860 23264 24912 23316
rect 10876 23239 10928 23248
rect 10876 23205 10885 23239
rect 10885 23205 10919 23239
rect 10919 23205 10928 23239
rect 10876 23196 10928 23205
rect 12440 23239 12492 23248
rect 12440 23205 12449 23239
rect 12449 23205 12483 23239
rect 12483 23205 12492 23239
rect 12440 23196 12492 23205
rect 112 23128 164 23180
rect 4068 23171 4120 23180
rect 4068 23137 4112 23171
rect 4112 23137 4120 23171
rect 4068 23128 4120 23137
rect 8300 23128 8352 23180
rect 9864 23128 9916 23180
rect 22836 23171 22888 23180
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 10784 23103 10836 23112
rect 10784 23069 10793 23103
rect 10793 23069 10827 23103
rect 10827 23069 10836 23103
rect 10784 23060 10836 23069
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 13452 23060 13504 23112
rect 12808 22992 12860 23044
rect 3240 22924 3292 22976
rect 9220 22924 9272 22976
rect 9312 22924 9364 22976
rect 10140 22924 10192 22976
rect 10416 22967 10468 22976
rect 10416 22933 10425 22967
rect 10425 22933 10459 22967
rect 10459 22933 10468 22967
rect 10416 22924 10468 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 4068 22763 4120 22772
rect 4068 22729 4077 22763
rect 4077 22729 4111 22763
rect 4111 22729 4120 22763
rect 4068 22720 4120 22729
rect 8852 22763 8904 22772
rect 8852 22729 8861 22763
rect 8861 22729 8895 22763
rect 8895 22729 8904 22763
rect 8852 22720 8904 22729
rect 9312 22763 9364 22772
rect 9312 22729 9321 22763
rect 9321 22729 9355 22763
rect 9355 22729 9364 22763
rect 9312 22720 9364 22729
rect 9864 22720 9916 22772
rect 12440 22720 12492 22772
rect 13452 22763 13504 22772
rect 13452 22729 13461 22763
rect 13461 22729 13495 22763
rect 13495 22729 13504 22763
rect 13452 22720 13504 22729
rect 10416 22627 10468 22636
rect 10416 22593 10425 22627
rect 10425 22593 10459 22627
rect 10459 22593 10468 22627
rect 10416 22584 10468 22593
rect 11060 22627 11112 22636
rect 11060 22593 11069 22627
rect 11069 22593 11103 22627
rect 11103 22593 11112 22627
rect 11060 22584 11112 22593
rect 12532 22627 12584 22636
rect 12532 22593 12541 22627
rect 12541 22593 12575 22627
rect 12575 22593 12584 22627
rect 12532 22584 12584 22593
rect 12808 22627 12860 22636
rect 12808 22593 12817 22627
rect 12817 22593 12851 22627
rect 12851 22593 12860 22627
rect 12808 22584 12860 22593
rect 7748 22516 7800 22568
rect 9312 22516 9364 22568
rect 7472 22423 7524 22432
rect 7472 22389 7481 22423
rect 7481 22389 7515 22423
rect 7515 22389 7524 22423
rect 7472 22380 7524 22389
rect 8300 22423 8352 22432
rect 8300 22389 8309 22423
rect 8309 22389 8343 22423
rect 8343 22389 8352 22423
rect 8300 22380 8352 22389
rect 10140 22423 10192 22432
rect 10140 22389 10149 22423
rect 10149 22389 10183 22423
rect 10183 22389 10192 22423
rect 10140 22380 10192 22389
rect 10876 22380 10928 22432
rect 12348 22380 12400 22432
rect 22836 22423 22888 22432
rect 22836 22389 22845 22423
rect 22845 22389 22879 22423
rect 22879 22389 22888 22423
rect 22836 22380 22888 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 10784 22176 10836 22228
rect 12624 22176 12676 22228
rect 1216 22108 1268 22160
rect 7472 22108 7524 22160
rect 10140 22108 10192 22160
rect 12440 22108 12492 22160
rect 4528 22083 4580 22092
rect 4528 22049 4546 22083
rect 4546 22049 4580 22083
rect 4528 22040 4580 22049
rect 4896 22040 4948 22092
rect 10876 22083 10928 22092
rect 10876 22049 10885 22083
rect 10885 22049 10919 22083
rect 10919 22049 10928 22083
rect 10876 22040 10928 22049
rect 12348 22083 12400 22092
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 17040 22083 17092 22092
rect 17040 22049 17058 22083
rect 17058 22049 17092 22083
rect 17040 22040 17092 22049
rect 18880 22040 18932 22092
rect 8208 21972 8260 22024
rect 6920 21904 6972 21956
rect 7564 21904 7616 21956
rect 8300 21904 8352 21956
rect 8484 21947 8536 21956
rect 8484 21913 8493 21947
rect 8493 21913 8527 21947
rect 8527 21913 8536 21947
rect 8484 21904 8536 21913
rect 5264 21836 5316 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1216 21632 1268 21684
rect 4528 21675 4580 21684
rect 4528 21641 4537 21675
rect 4537 21641 4571 21675
rect 4571 21641 4580 21675
rect 4528 21632 4580 21641
rect 7472 21632 7524 21684
rect 8208 21675 8260 21684
rect 8208 21641 8217 21675
rect 8217 21641 8251 21675
rect 8251 21641 8260 21675
rect 8208 21632 8260 21641
rect 10876 21632 10928 21684
rect 17040 21675 17092 21684
rect 17040 21641 17049 21675
rect 17049 21641 17083 21675
rect 17083 21641 17092 21675
rect 17040 21632 17092 21641
rect 5264 21539 5316 21548
rect 5264 21505 5273 21539
rect 5273 21505 5307 21539
rect 5307 21505 5316 21539
rect 5264 21496 5316 21505
rect 5540 21539 5592 21548
rect 5540 21505 5549 21539
rect 5549 21505 5583 21539
rect 5583 21505 5592 21539
rect 5540 21496 5592 21505
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 8484 21539 8536 21548
rect 8484 21505 8493 21539
rect 8493 21505 8527 21539
rect 8527 21505 8536 21539
rect 8484 21496 8536 21505
rect 9128 21496 9180 21548
rect 9864 21496 9916 21548
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 4988 21335 5040 21344
rect 4988 21301 4997 21335
rect 4997 21301 5031 21335
rect 5031 21301 5040 21335
rect 7012 21403 7064 21412
rect 7012 21369 7021 21403
rect 7021 21369 7055 21403
rect 7055 21369 7064 21403
rect 8576 21403 8628 21412
rect 7012 21360 7064 21369
rect 8576 21369 8585 21403
rect 8585 21369 8619 21403
rect 8619 21369 8628 21403
rect 8576 21360 8628 21369
rect 10692 21403 10744 21412
rect 10692 21369 10701 21403
rect 10701 21369 10735 21403
rect 10735 21369 10744 21403
rect 10692 21360 10744 21369
rect 4988 21292 5040 21301
rect 11980 21360 12032 21412
rect 12348 21292 12400 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 6920 21131 6972 21140
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 6276 21020 6328 21072
rect 7012 21063 7064 21072
rect 7012 21029 7021 21063
rect 7021 21029 7055 21063
rect 7055 21029 7064 21063
rect 7012 21020 7064 21029
rect 7564 20952 7616 21004
rect 8300 20952 8352 21004
rect 8576 21088 8628 21140
rect 11980 20995 12032 21004
rect 11980 20961 11989 20995
rect 11989 20961 12023 20995
rect 12023 20961 12032 20995
rect 11980 20952 12032 20961
rect 25228 20952 25280 21004
rect 3976 20884 4028 20936
rect 5540 20927 5592 20936
rect 5540 20893 5549 20927
rect 5549 20893 5583 20927
rect 5583 20893 5592 20927
rect 5540 20884 5592 20893
rect 11244 20884 11296 20936
rect 11336 20884 11388 20936
rect 10968 20859 11020 20868
rect 10968 20825 10977 20859
rect 10977 20825 11011 20859
rect 11011 20825 11020 20859
rect 10968 20816 11020 20825
rect 5172 20791 5224 20800
rect 5172 20757 5181 20791
rect 5181 20757 5215 20791
rect 5215 20757 5224 20791
rect 5172 20748 5224 20757
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 18604 20748 18656 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 5540 20544 5592 20596
rect 6276 20587 6328 20596
rect 4712 20476 4764 20528
rect 5172 20476 5224 20528
rect 6276 20553 6285 20587
rect 6285 20553 6319 20587
rect 6319 20553 6328 20587
rect 7748 20587 7800 20596
rect 6276 20544 6328 20553
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 11336 20544 11388 20596
rect 24768 20587 24820 20596
rect 24768 20553 24777 20587
rect 24777 20553 24811 20587
rect 24811 20553 24820 20587
rect 24768 20544 24820 20553
rect 25228 20587 25280 20596
rect 25228 20553 25237 20587
rect 25237 20553 25271 20587
rect 25271 20553 25280 20587
rect 25228 20544 25280 20553
rect 26884 20544 26936 20596
rect 4988 20408 5040 20460
rect 10876 20476 10928 20528
rect 11244 20519 11296 20528
rect 11244 20485 11253 20519
rect 11253 20485 11287 20519
rect 11287 20485 11296 20519
rect 11244 20476 11296 20485
rect 11980 20519 12032 20528
rect 11980 20485 11989 20519
rect 11989 20485 12023 20519
rect 12023 20485 12032 20519
rect 11980 20476 12032 20485
rect 10784 20408 10836 20460
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 1676 20340 1728 20392
rect 6736 20340 6788 20392
rect 7748 20340 7800 20392
rect 10692 20340 10744 20392
rect 5356 20315 5408 20324
rect 5356 20281 5365 20315
rect 5365 20281 5399 20315
rect 5399 20281 5408 20315
rect 5356 20272 5408 20281
rect 6276 20204 6328 20256
rect 9864 20272 9916 20324
rect 12992 20315 13044 20324
rect 12992 20281 13001 20315
rect 13001 20281 13035 20315
rect 13035 20281 13044 20315
rect 12992 20272 13044 20281
rect 9404 20204 9456 20256
rect 18604 20204 18656 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1952 20000 2004 20052
rect 5356 20000 5408 20052
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 11980 20000 12032 20052
rect 12348 20043 12400 20052
rect 12348 20009 12357 20043
rect 12357 20009 12391 20043
rect 12391 20009 12400 20043
rect 12348 20000 12400 20009
rect 6276 19932 6328 19984
rect 7656 19975 7708 19984
rect 7656 19941 7665 19975
rect 7665 19941 7699 19975
rect 7699 19941 7708 19975
rect 7656 19932 7708 19941
rect 9864 19932 9916 19984
rect 11428 19932 11480 19984
rect 12992 19932 13044 19984
rect 1952 19864 2004 19916
rect 3424 19864 3476 19916
rect 4620 19864 4672 19916
rect 13728 19907 13780 19916
rect 13728 19873 13737 19907
rect 13737 19873 13771 19907
rect 13771 19873 13780 19907
rect 13728 19864 13780 19873
rect 5448 19839 5500 19848
rect 5448 19805 5457 19839
rect 5457 19805 5491 19839
rect 5491 19805 5500 19839
rect 5448 19796 5500 19805
rect 8208 19796 8260 19848
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 11704 19796 11756 19848
rect 2044 19660 2096 19712
rect 3884 19660 3936 19712
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 6736 19660 6788 19712
rect 12808 19703 12860 19712
rect 12808 19669 12817 19703
rect 12817 19669 12851 19703
rect 12851 19669 12860 19703
rect 12808 19660 12860 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1676 19499 1728 19508
rect 1676 19465 1685 19499
rect 1685 19465 1719 19499
rect 1719 19465 1728 19499
rect 1676 19456 1728 19465
rect 2872 19456 2924 19508
rect 6276 19456 6328 19508
rect 7656 19456 7708 19508
rect 9864 19499 9916 19508
rect 9864 19465 9873 19499
rect 9873 19465 9907 19499
rect 9907 19465 9916 19499
rect 11428 19499 11480 19508
rect 9864 19456 9916 19465
rect 11428 19465 11437 19499
rect 11437 19465 11471 19499
rect 11471 19465 11480 19499
rect 11428 19456 11480 19465
rect 13728 19499 13780 19508
rect 13728 19465 13737 19499
rect 13737 19465 13771 19499
rect 13771 19465 13780 19499
rect 13728 19456 13780 19465
rect 5172 19388 5224 19440
rect 940 19320 992 19372
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 2872 19252 2924 19304
rect 4068 19294 4120 19346
rect 4344 19320 4396 19372
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 4436 19252 4488 19304
rect 5172 19295 5224 19304
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 6736 19320 6788 19372
rect 8024 19320 8076 19372
rect 7288 19295 7340 19304
rect 2412 19116 2464 19168
rect 2964 19116 3016 19168
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 4068 19116 4120 19168
rect 5356 19184 5408 19236
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 9680 19320 9732 19372
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 10876 19295 10928 19304
rect 10876 19261 10885 19295
rect 10885 19261 10919 19295
rect 10919 19261 10928 19295
rect 10876 19252 10928 19261
rect 12808 19227 12860 19236
rect 12808 19193 12817 19227
rect 12817 19193 12851 19227
rect 12851 19193 12860 19227
rect 12808 19184 12860 19193
rect 12900 19227 12952 19236
rect 12900 19193 12909 19227
rect 12909 19193 12943 19227
rect 12943 19193 12952 19227
rect 12900 19184 12952 19193
rect 13728 19184 13780 19236
rect 4436 19116 4488 19168
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 4804 19116 4856 19168
rect 6276 19159 6328 19168
rect 6276 19125 6285 19159
rect 6285 19125 6319 19159
rect 6319 19125 6328 19159
rect 6276 19116 6328 19125
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 8208 19159 8260 19168
rect 8208 19125 8217 19159
rect 8217 19125 8251 19159
rect 8251 19125 8260 19159
rect 8208 19116 8260 19125
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 10692 19116 10744 19125
rect 11704 19116 11756 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 5356 18955 5408 18964
rect 5356 18921 5365 18955
rect 5365 18921 5399 18955
rect 5399 18921 5408 18955
rect 5356 18912 5408 18921
rect 5448 18912 5500 18964
rect 6920 18912 6972 18964
rect 9680 18912 9732 18964
rect 12900 18912 12952 18964
rect 24768 18955 24820 18964
rect 24768 18921 24777 18955
rect 24777 18921 24811 18955
rect 24811 18921 24820 18955
rect 24768 18912 24820 18921
rect 6000 18887 6052 18896
rect 6000 18853 6009 18887
rect 6009 18853 6043 18887
rect 6043 18853 6052 18887
rect 6000 18844 6052 18853
rect 7564 18887 7616 18896
rect 7564 18853 7573 18887
rect 7573 18853 7607 18887
rect 7607 18853 7616 18887
rect 7564 18844 7616 18853
rect 8484 18844 8536 18896
rect 10876 18844 10928 18896
rect 11428 18844 11480 18896
rect 1768 18776 1820 18828
rect 2320 18776 2372 18828
rect 3056 18776 3108 18828
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 8116 18776 8168 18828
rect 9864 18776 9916 18828
rect 13176 18819 13228 18828
rect 5540 18708 5592 18760
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 7472 18751 7524 18760
rect 7472 18717 7481 18751
rect 7481 18717 7515 18751
rect 7515 18717 7524 18751
rect 7472 18708 7524 18717
rect 7748 18751 7800 18760
rect 7748 18717 7757 18751
rect 7757 18717 7791 18751
rect 7791 18717 7800 18751
rect 7748 18708 7800 18717
rect 5080 18572 5132 18624
rect 7288 18572 7340 18624
rect 7840 18572 7892 18624
rect 8668 18572 8720 18624
rect 9312 18708 9364 18760
rect 13176 18785 13185 18819
rect 13185 18785 13219 18819
rect 13219 18785 13228 18819
rect 13176 18776 13228 18785
rect 15660 18776 15712 18828
rect 24584 18819 24636 18828
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 25412 18776 25464 18828
rect 11796 18708 11848 18760
rect 13820 18751 13872 18760
rect 13820 18717 13829 18751
rect 13829 18717 13863 18751
rect 13863 18717 13872 18751
rect 13820 18708 13872 18717
rect 10508 18640 10560 18692
rect 18236 18640 18288 18692
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 2044 18411 2096 18420
rect 2044 18377 2053 18411
rect 2053 18377 2087 18411
rect 2087 18377 2096 18411
rect 2044 18368 2096 18377
rect 2320 18411 2372 18420
rect 2320 18377 2329 18411
rect 2329 18377 2363 18411
rect 2363 18377 2372 18411
rect 2320 18368 2372 18377
rect 3056 18368 3108 18420
rect 4160 18368 4212 18420
rect 4804 18368 4856 18420
rect 4896 18368 4948 18420
rect 6000 18368 6052 18420
rect 9864 18411 9916 18420
rect 4344 18343 4396 18352
rect 4344 18309 4353 18343
rect 4353 18309 4387 18343
rect 4387 18309 4396 18343
rect 4344 18300 4396 18309
rect 7564 18300 7616 18352
rect 6184 18232 6236 18284
rect 7748 18232 7800 18284
rect 2044 18164 2096 18216
rect 2504 18164 2556 18216
rect 4252 18164 4304 18216
rect 4896 18164 4948 18216
rect 6644 18164 6696 18216
rect 7104 18139 7156 18148
rect 7104 18105 7113 18139
rect 7113 18105 7147 18139
rect 7147 18105 7156 18139
rect 9864 18377 9873 18411
rect 9873 18377 9907 18411
rect 9907 18377 9916 18411
rect 9864 18368 9916 18377
rect 11428 18411 11480 18420
rect 11428 18377 11437 18411
rect 11437 18377 11471 18411
rect 11471 18377 11480 18411
rect 11428 18368 11480 18377
rect 11796 18411 11848 18420
rect 11796 18377 11805 18411
rect 11805 18377 11839 18411
rect 11839 18377 11848 18411
rect 11796 18368 11848 18377
rect 13176 18411 13228 18420
rect 13176 18377 13185 18411
rect 13185 18377 13219 18411
rect 13219 18377 13228 18411
rect 13176 18368 13228 18377
rect 25412 18411 25464 18420
rect 25412 18377 25421 18411
rect 25421 18377 25455 18411
rect 25455 18377 25464 18411
rect 25412 18368 25464 18377
rect 24584 18300 24636 18352
rect 8760 18232 8812 18284
rect 7104 18096 7156 18105
rect 4252 18028 4304 18080
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 6644 18071 6696 18080
rect 6644 18037 6653 18071
rect 6653 18037 6687 18071
rect 6687 18037 6696 18071
rect 6644 18028 6696 18037
rect 9220 18096 9272 18148
rect 10048 18096 10100 18148
rect 10508 18139 10560 18148
rect 10508 18105 10517 18139
rect 10517 18105 10551 18139
rect 10551 18105 10560 18139
rect 10508 18096 10560 18105
rect 11152 18139 11204 18148
rect 10140 18028 10192 18080
rect 11152 18105 11161 18139
rect 11161 18105 11195 18139
rect 11195 18105 11204 18139
rect 11152 18096 11204 18105
rect 14004 18139 14056 18148
rect 14004 18105 14013 18139
rect 14013 18105 14047 18139
rect 14047 18105 14056 18139
rect 14004 18096 14056 18105
rect 11888 18028 11940 18080
rect 13452 18028 13504 18080
rect 27620 18232 27672 18284
rect 15476 18139 15528 18148
rect 15476 18105 15485 18139
rect 15485 18105 15519 18139
rect 15519 18105 15528 18139
rect 15476 18096 15528 18105
rect 15660 18028 15712 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 4896 17867 4948 17876
rect 4896 17833 4905 17867
rect 4905 17833 4939 17867
rect 4939 17833 4948 17867
rect 4896 17824 4948 17833
rect 5540 17824 5592 17876
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 12716 17824 12768 17876
rect 4988 17756 5040 17808
rect 6000 17756 6052 17808
rect 6184 17799 6236 17808
rect 6184 17765 6193 17799
rect 6193 17765 6227 17799
rect 6227 17765 6236 17799
rect 6184 17756 6236 17765
rect 10048 17756 10100 17808
rect 10140 17756 10192 17808
rect 12992 17799 13044 17808
rect 12992 17765 13001 17799
rect 13001 17765 13035 17799
rect 13035 17765 13044 17799
rect 12992 17756 13044 17765
rect 13176 17756 13228 17808
rect 15476 17799 15528 17808
rect 15476 17765 15485 17799
rect 15485 17765 15519 17799
rect 15519 17765 15528 17799
rect 15476 17756 15528 17765
rect 2872 17688 2924 17740
rect 4252 17688 4304 17740
rect 8024 17731 8076 17740
rect 8024 17697 8033 17731
rect 8033 17697 8067 17731
rect 8067 17697 8076 17731
rect 8024 17688 8076 17697
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 10324 17731 10376 17740
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 11888 17688 11940 17740
rect 5172 17620 5224 17672
rect 11704 17620 11756 17672
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 1492 17484 1544 17536
rect 2044 17484 2096 17536
rect 4160 17484 4212 17536
rect 5264 17527 5316 17536
rect 5264 17493 5273 17527
rect 5273 17493 5307 17527
rect 5307 17493 5316 17527
rect 5264 17484 5316 17493
rect 8668 17484 8720 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 15568 17552 15620 17604
rect 14004 17527 14056 17536
rect 14004 17493 14013 17527
rect 14013 17493 14047 17527
rect 14047 17493 14056 17527
rect 14004 17484 14056 17493
rect 14648 17484 14700 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 6000 17280 6052 17332
rect 6276 17280 6328 17332
rect 6644 17280 6696 17332
rect 7104 17280 7156 17332
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 10968 17280 11020 17332
rect 11888 17323 11940 17332
rect 11888 17289 11897 17323
rect 11897 17289 11931 17323
rect 11931 17289 11940 17323
rect 11888 17280 11940 17289
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 13820 17280 13872 17332
rect 14464 17280 14516 17332
rect 15476 17280 15528 17332
rect 13176 17212 13228 17264
rect 9220 17187 9272 17196
rect 1492 17076 1544 17128
rect 3700 17076 3752 17128
rect 3884 17008 3936 17060
rect 4344 17051 4396 17060
rect 4344 17017 4353 17051
rect 4353 17017 4387 17051
rect 4387 17017 4396 17051
rect 4344 17008 4396 17017
rect 5264 17076 5316 17128
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 6092 17008 6144 17060
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 11152 17187 11204 17196
rect 11152 17153 11161 17187
rect 11161 17153 11195 17187
rect 11195 17153 11204 17187
rect 11152 17144 11204 17153
rect 14004 17144 14056 17196
rect 8300 17076 8352 17128
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 9864 17076 9916 17085
rect 12532 17119 12584 17128
rect 12532 17085 12541 17119
rect 12541 17085 12575 17119
rect 12575 17085 12584 17119
rect 12532 17076 12584 17085
rect 8760 17008 8812 17060
rect 10876 17051 10928 17060
rect 10876 17017 10885 17051
rect 10885 17017 10919 17051
rect 10919 17017 10928 17051
rect 10876 17008 10928 17017
rect 10968 17051 11020 17060
rect 10968 17017 10977 17051
rect 10977 17017 11011 17051
rect 11011 17017 11020 17051
rect 10968 17008 11020 17017
rect 1860 16983 1912 16992
rect 1860 16949 1869 16983
rect 1869 16949 1903 16983
rect 1903 16949 1912 16983
rect 1860 16940 1912 16949
rect 2872 16940 2924 16992
rect 4252 16940 4304 16992
rect 5080 16983 5132 16992
rect 5080 16949 5089 16983
rect 5089 16949 5123 16983
rect 5123 16949 5132 16983
rect 5080 16940 5132 16949
rect 7288 16940 7340 16992
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 12164 16983 12216 16992
rect 12164 16949 12173 16983
rect 12173 16949 12207 16983
rect 12207 16949 12216 16983
rect 12164 16940 12216 16949
rect 14464 17051 14516 17060
rect 14464 17017 14473 17051
rect 14473 17017 14507 17051
rect 14507 17017 14516 17051
rect 14464 17008 14516 17017
rect 14648 16940 14700 16992
rect 15660 16983 15712 16992
rect 15660 16949 15669 16983
rect 15669 16949 15703 16983
rect 15703 16949 15712 16983
rect 15660 16940 15712 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3700 16779 3752 16788
rect 3700 16745 3709 16779
rect 3709 16745 3743 16779
rect 3743 16745 3752 16779
rect 3700 16736 3752 16745
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 6000 16736 6052 16788
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7472 16736 7524 16788
rect 10968 16736 11020 16788
rect 13176 16736 13228 16788
rect 5356 16668 5408 16720
rect 6276 16668 6328 16720
rect 6552 16668 6604 16720
rect 8300 16668 8352 16720
rect 8760 16711 8812 16720
rect 8760 16677 8769 16711
rect 8769 16677 8803 16711
rect 8803 16677 8812 16711
rect 8760 16668 8812 16677
rect 9588 16668 9640 16720
rect 10876 16711 10928 16720
rect 10876 16677 10885 16711
rect 10885 16677 10919 16711
rect 10919 16677 10928 16711
rect 10876 16668 10928 16677
rect 12164 16668 12216 16720
rect 1584 16600 1636 16652
rect 2964 16643 3016 16652
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 3608 16600 3660 16652
rect 4344 16600 4396 16652
rect 5448 16600 5500 16652
rect 12992 16600 13044 16652
rect 4620 16532 4672 16584
rect 3516 16464 3568 16516
rect 5172 16464 5224 16516
rect 1676 16396 1728 16448
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 2780 16396 2832 16448
rect 7104 16396 7156 16448
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 9680 16532 9732 16541
rect 11980 16575 12032 16584
rect 11980 16541 11989 16575
rect 11989 16541 12023 16575
rect 12023 16541 12032 16575
rect 11980 16532 12032 16541
rect 12532 16532 12584 16584
rect 15660 16668 15712 16720
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 15292 16532 15344 16584
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 3608 16235 3660 16244
rect 3608 16201 3617 16235
rect 3617 16201 3651 16235
rect 3651 16201 3660 16235
rect 3608 16192 3660 16201
rect 5356 16235 5408 16244
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 9680 16192 9732 16244
rect 11980 16192 12032 16244
rect 9864 16124 9916 16176
rect 9588 16056 9640 16108
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 4252 16031 4304 16040
rect 4252 15997 4261 16031
rect 4261 15997 4295 16031
rect 4295 15997 4304 16031
rect 4252 15988 4304 15997
rect 4896 16031 4948 16040
rect 4896 15997 4905 16031
rect 4905 15997 4939 16031
rect 4939 15997 4948 16031
rect 4896 15988 4948 15997
rect 8760 16031 8812 16040
rect 2228 15920 2280 15972
rect 7380 15920 7432 15972
rect 8760 15997 8769 16031
rect 8769 15997 8803 16031
rect 8803 15997 8812 16031
rect 8760 15988 8812 15997
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 2136 15895 2188 15904
rect 2136 15861 2145 15895
rect 2145 15861 2179 15895
rect 2179 15861 2188 15895
rect 2136 15852 2188 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 9864 15988 9916 16040
rect 13544 16056 13596 16108
rect 10140 16031 10192 16040
rect 10140 15997 10149 16031
rect 10149 15997 10183 16031
rect 10183 15997 10192 16031
rect 10140 15988 10192 15997
rect 12164 15920 12216 15972
rect 12900 15920 12952 15972
rect 13360 15852 13412 15904
rect 13544 15963 13596 15972
rect 13544 15929 13553 15963
rect 13553 15929 13587 15963
rect 13587 15929 13596 15963
rect 14096 15963 14148 15972
rect 13544 15920 13596 15929
rect 14096 15929 14105 15963
rect 14105 15929 14139 15963
rect 14139 15929 14148 15963
rect 14096 15920 14148 15929
rect 15292 15988 15344 16040
rect 24676 16031 24728 16040
rect 24676 15997 24694 16031
rect 24694 15997 24728 16031
rect 24676 15988 24728 15997
rect 15476 15920 15528 15972
rect 18420 15920 18472 15972
rect 20720 15920 20772 15972
rect 14280 15852 14332 15904
rect 15568 15852 15620 15904
rect 18604 15852 18656 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1124 15648 1176 15700
rect 3976 15648 4028 15700
rect 5448 15691 5500 15700
rect 2136 15623 2188 15632
rect 2136 15589 2145 15623
rect 2145 15589 2179 15623
rect 2179 15589 2188 15623
rect 2136 15580 2188 15589
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 10140 15648 10192 15700
rect 13544 15648 13596 15700
rect 4620 15623 4672 15632
rect 4620 15589 4629 15623
rect 4629 15589 4663 15623
rect 4663 15589 4672 15623
rect 4620 15580 4672 15589
rect 4896 15580 4948 15632
rect 6368 15555 6420 15564
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 7380 15512 7432 15564
rect 7748 15512 7800 15564
rect 8760 15512 8812 15564
rect 9128 15580 9180 15632
rect 9588 15580 9640 15632
rect 11428 15580 11480 15632
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 13820 15580 13872 15589
rect 10324 15512 10376 15564
rect 15384 15555 15436 15564
rect 15384 15521 15393 15555
rect 15393 15521 15427 15555
rect 15427 15521 15436 15555
rect 15384 15512 15436 15521
rect 24676 15512 24728 15564
rect 5172 15487 5224 15496
rect 5172 15453 5181 15487
rect 5181 15453 5215 15487
rect 5215 15453 5224 15487
rect 5172 15444 5224 15453
rect 5356 15444 5408 15496
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 11244 15444 11296 15453
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 2596 15419 2648 15428
rect 2596 15385 2605 15419
rect 2605 15385 2639 15419
rect 2639 15385 2648 15419
rect 2596 15376 2648 15385
rect 14280 15376 14332 15428
rect 15292 15376 15344 15428
rect 24768 15419 24820 15428
rect 24768 15385 24777 15419
rect 24777 15385 24811 15419
rect 24811 15385 24820 15419
rect 24768 15376 24820 15385
rect 7656 15308 7708 15360
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2136 15104 2188 15156
rect 2964 15104 3016 15156
rect 4620 15147 4672 15156
rect 4620 15113 4629 15147
rect 4629 15113 4663 15147
rect 4663 15113 4672 15147
rect 4620 15104 4672 15113
rect 7748 15104 7800 15156
rect 8760 15104 8812 15156
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 13820 15104 13872 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 1676 14968 1728 15020
rect 5172 15036 5224 15088
rect 8208 15079 8260 15088
rect 8208 15045 8217 15079
rect 8217 15045 8251 15079
rect 8251 15045 8260 15079
rect 8208 15036 8260 15045
rect 11520 15036 11572 15088
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 3700 15011 3752 15020
rect 2596 14968 2648 14977
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 3700 14968 3752 14977
rect 4160 14968 4212 15020
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 6828 14968 6880 15020
rect 6000 14900 6052 14952
rect 11244 14968 11296 15020
rect 12716 14968 12768 15020
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 7748 14900 7800 14952
rect 8208 14943 8260 14952
rect 8208 14909 8217 14943
rect 8217 14909 8251 14943
rect 8251 14909 8260 14943
rect 8208 14900 8260 14909
rect 8392 14943 8444 14952
rect 8392 14909 8401 14943
rect 8401 14909 8435 14943
rect 8435 14909 8444 14943
rect 8392 14900 8444 14909
rect 8760 14900 8812 14952
rect 15292 14900 15344 14952
rect 24124 14943 24176 14952
rect 1952 14832 2004 14884
rect 3792 14875 3844 14884
rect 3792 14841 3801 14875
rect 3801 14841 3835 14875
rect 3835 14841 3844 14875
rect 3792 14832 3844 14841
rect 5356 14875 5408 14884
rect 5356 14841 5365 14875
rect 5365 14841 5399 14875
rect 5399 14841 5408 14875
rect 6276 14875 6328 14884
rect 5356 14832 5408 14841
rect 6276 14841 6285 14875
rect 6285 14841 6319 14875
rect 6319 14841 6328 14875
rect 6276 14832 6328 14841
rect 9128 14832 9180 14884
rect 9496 14875 9548 14884
rect 9496 14841 9505 14875
rect 9505 14841 9539 14875
rect 9539 14841 9548 14875
rect 9496 14832 9548 14841
rect 12532 14875 12584 14884
rect 12532 14841 12541 14875
rect 12541 14841 12575 14875
rect 12575 14841 12584 14875
rect 12532 14832 12584 14841
rect 6736 14764 6788 14816
rect 7380 14764 7432 14816
rect 8208 14764 8260 14816
rect 8944 14764 8996 14816
rect 11428 14807 11480 14816
rect 11428 14773 11437 14807
rect 11437 14773 11471 14807
rect 11471 14773 11480 14807
rect 11428 14764 11480 14773
rect 12808 14832 12860 14884
rect 14096 14875 14148 14884
rect 14096 14841 14105 14875
rect 14105 14841 14139 14875
rect 14139 14841 14148 14875
rect 14096 14832 14148 14841
rect 14004 14764 14056 14816
rect 14832 14832 14884 14884
rect 24124 14909 24133 14943
rect 24133 14909 24167 14943
rect 24167 14909 24176 14943
rect 24124 14900 24176 14909
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1952 14560 2004 14612
rect 3700 14603 3752 14612
rect 3700 14569 3709 14603
rect 3709 14569 3743 14603
rect 3743 14569 3752 14603
rect 3700 14560 3752 14569
rect 3792 14560 3844 14612
rect 5264 14603 5316 14612
rect 5264 14569 5273 14603
rect 5273 14569 5307 14603
rect 5307 14569 5316 14603
rect 5264 14560 5316 14569
rect 6368 14603 6420 14612
rect 6368 14569 6377 14603
rect 6377 14569 6411 14603
rect 6411 14569 6420 14603
rect 6368 14560 6420 14569
rect 6828 14560 6880 14612
rect 12532 14603 12584 14612
rect 1676 14535 1728 14544
rect 1676 14501 1685 14535
rect 1685 14501 1719 14535
rect 1719 14501 1728 14535
rect 1676 14492 1728 14501
rect 2228 14492 2280 14544
rect 2596 14535 2648 14544
rect 2596 14501 2599 14535
rect 2599 14501 2633 14535
rect 2633 14501 2648 14535
rect 2596 14492 2648 14501
rect 3976 14492 4028 14544
rect 6552 14492 6604 14544
rect 6000 14424 6052 14476
rect 7656 14492 7708 14544
rect 8760 14492 8812 14544
rect 10784 14492 10836 14544
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 12900 14560 12952 14612
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 14004 14603 14056 14612
rect 14004 14569 14013 14603
rect 14013 14569 14047 14603
rect 14047 14569 14056 14603
rect 14004 14560 14056 14569
rect 14096 14560 14148 14612
rect 11428 14492 11480 14544
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 4252 14356 4304 14408
rect 8392 14424 8444 14476
rect 12072 14424 12124 14476
rect 9864 14356 9916 14408
rect 5540 14220 5592 14272
rect 8760 14220 8812 14272
rect 9036 14220 9088 14272
rect 9496 14220 9548 14272
rect 11888 14220 11940 14272
rect 12808 14424 12860 14476
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15384 14288 15436 14340
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2320 14016 2372 14068
rect 2596 14016 2648 14068
rect 3976 14016 4028 14068
rect 6000 14016 6052 14068
rect 6276 14059 6328 14068
rect 6276 14025 6285 14059
rect 6285 14025 6319 14059
rect 6319 14025 6328 14059
rect 6276 14016 6328 14025
rect 6368 14016 6420 14068
rect 9036 14016 9088 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 14004 14016 14056 14068
rect 14556 14016 14608 14068
rect 14832 14016 14884 14068
rect 15384 14016 15436 14068
rect 6552 13991 6604 14000
rect 6552 13957 6561 13991
rect 6561 13957 6595 13991
rect 6595 13957 6604 13991
rect 6552 13948 6604 13957
rect 8852 13991 8904 14000
rect 8852 13957 8861 13991
rect 8861 13957 8895 13991
rect 8895 13957 8904 13991
rect 8852 13948 8904 13957
rect 10784 13948 10836 14000
rect 12256 13948 12308 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2688 13812 2740 13864
rect 3424 13812 3476 13864
rect 4068 13880 4120 13932
rect 6828 13923 6880 13932
rect 4252 13855 4304 13864
rect 4252 13821 4261 13855
rect 4261 13821 4295 13855
rect 4295 13821 4304 13855
rect 4252 13812 4304 13821
rect 1676 13744 1728 13796
rect 1860 13744 1912 13796
rect 4528 13812 4580 13864
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 8576 13880 8628 13932
rect 5540 13855 5592 13864
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 9864 13880 9916 13932
rect 14096 13880 14148 13932
rect 14740 13923 14792 13932
rect 14740 13889 14749 13923
rect 14749 13889 14783 13923
rect 14783 13889 14792 13923
rect 14740 13880 14792 13889
rect 14832 13880 14884 13932
rect 6552 13744 6604 13796
rect 7380 13744 7432 13796
rect 8760 13744 8812 13796
rect 3884 13676 3936 13728
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 11980 13812 12032 13864
rect 18236 13855 18288 13864
rect 18236 13821 18245 13855
rect 18245 13821 18279 13855
rect 18279 13821 18288 13855
rect 18236 13812 18288 13821
rect 11704 13744 11756 13796
rect 14832 13787 14884 13796
rect 14832 13753 14841 13787
rect 14841 13753 14875 13787
rect 14875 13753 14884 13787
rect 14832 13744 14884 13753
rect 16212 13787 16264 13796
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 16212 13744 16264 13753
rect 9864 13676 9916 13685
rect 11796 13676 11848 13728
rect 12072 13676 12124 13728
rect 12900 13676 12952 13728
rect 14372 13676 14424 13728
rect 18420 13719 18472 13728
rect 18420 13685 18429 13719
rect 18429 13685 18463 13719
rect 18463 13685 18472 13719
rect 18420 13676 18472 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1676 13515 1728 13524
rect 1676 13481 1685 13515
rect 1685 13481 1719 13515
rect 1719 13481 1728 13515
rect 1676 13472 1728 13481
rect 2228 13472 2280 13524
rect 4528 13472 4580 13524
rect 1492 13404 1544 13456
rect 1952 13404 2004 13456
rect 2688 13404 2740 13456
rect 4160 13379 4212 13388
rect 4160 13345 4169 13379
rect 4169 13345 4203 13379
rect 4203 13345 4212 13379
rect 4160 13336 4212 13345
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 4528 13336 4580 13345
rect 2136 13268 2188 13320
rect 7380 13472 7432 13524
rect 6092 13404 6144 13456
rect 6736 13404 6788 13456
rect 10784 13472 10836 13524
rect 11704 13472 11756 13524
rect 11980 13515 12032 13524
rect 11980 13481 11989 13515
rect 11989 13481 12023 13515
rect 12023 13481 12032 13515
rect 11980 13472 12032 13481
rect 12072 13472 12124 13524
rect 18236 13472 18288 13524
rect 12256 13447 12308 13456
rect 6276 13336 6328 13388
rect 6644 13336 6696 13388
rect 7380 13268 7432 13320
rect 9680 13336 9732 13388
rect 12256 13413 12265 13447
rect 12265 13413 12299 13447
rect 12299 13413 12308 13447
rect 12256 13404 12308 13413
rect 12624 13404 12676 13456
rect 12808 13447 12860 13456
rect 12808 13413 12817 13447
rect 12817 13413 12851 13447
rect 12851 13413 12860 13447
rect 12808 13404 12860 13413
rect 12992 13404 13044 13456
rect 2412 13200 2464 13252
rect 4988 13200 5040 13252
rect 8024 13200 8076 13252
rect 8576 13200 8628 13252
rect 9128 13200 9180 13252
rect 9772 13200 9824 13252
rect 10784 13268 10836 13320
rect 13176 13336 13228 13388
rect 3700 13132 3752 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 7012 13132 7064 13141
rect 7748 13132 7800 13184
rect 8300 13132 8352 13184
rect 8852 13132 8904 13184
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 11060 13132 11112 13184
rect 14280 13336 14332 13388
rect 14648 13336 14700 13388
rect 14832 13336 14884 13388
rect 15568 13336 15620 13388
rect 16028 13336 16080 13388
rect 17316 13336 17368 13388
rect 24676 13336 24728 13388
rect 14372 13268 14424 13320
rect 13544 13200 13596 13252
rect 14188 13200 14240 13252
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 15384 13132 15436 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1768 12928 1820 12980
rect 1952 12928 2004 12980
rect 4528 12928 4580 12980
rect 6368 12928 6420 12980
rect 8116 12928 8168 12980
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 8760 12928 8812 12980
rect 9956 12928 10008 12980
rect 13176 12928 13228 12980
rect 14188 12971 14240 12980
rect 14188 12937 14212 12971
rect 14212 12937 14240 12971
rect 14188 12928 14240 12937
rect 14464 12971 14516 12980
rect 14464 12937 14473 12971
rect 14473 12937 14507 12971
rect 14507 12937 14516 12971
rect 14464 12928 14516 12937
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 2320 12903 2372 12912
rect 2320 12869 2329 12903
rect 2329 12869 2363 12903
rect 2363 12869 2372 12903
rect 2320 12860 2372 12869
rect 4160 12860 4212 12912
rect 7380 12860 7432 12912
rect 7472 12860 7524 12912
rect 8300 12903 8352 12912
rect 8300 12869 8309 12903
rect 8309 12869 8343 12903
rect 8343 12869 8352 12903
rect 8300 12860 8352 12869
rect 9588 12860 9640 12912
rect 9772 12903 9824 12912
rect 9772 12869 9796 12903
rect 9796 12869 9824 12903
rect 9772 12860 9824 12869
rect 2872 12792 2924 12844
rect 8024 12792 8076 12844
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 8576 12792 8628 12844
rect 9036 12792 9088 12844
rect 12808 12860 12860 12912
rect 13912 12860 13964 12912
rect 14280 12903 14332 12912
rect 14280 12869 14289 12903
rect 14289 12869 14323 12903
rect 14323 12869 14332 12903
rect 14280 12860 14332 12869
rect 14832 12860 14884 12912
rect 10048 12792 10100 12844
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 14372 12835 14424 12844
rect 1768 12724 1820 12776
rect 2412 12767 2464 12776
rect 2412 12733 2421 12767
rect 2421 12733 2455 12767
rect 2455 12733 2464 12767
rect 2412 12724 2464 12733
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 7012 12767 7064 12776
rect 5448 12724 5500 12733
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 8300 12724 8352 12776
rect 13452 12724 13504 12776
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 14464 12792 14516 12844
rect 15384 12724 15436 12776
rect 15476 12724 15528 12776
rect 16028 12767 16080 12776
rect 16028 12733 16037 12767
rect 16037 12733 16071 12767
rect 16071 12733 16080 12767
rect 16028 12724 16080 12733
rect 2320 12656 2372 12708
rect 2688 12656 2740 12708
rect 7748 12656 7800 12708
rect 8668 12656 8720 12708
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 7564 12588 7616 12640
rect 8392 12588 8444 12640
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 9680 12656 9732 12708
rect 10876 12656 10928 12708
rect 16212 12656 16264 12708
rect 9772 12588 9824 12640
rect 10048 12588 10100 12640
rect 15660 12631 15712 12640
rect 15660 12597 15669 12631
rect 15669 12597 15703 12631
rect 15703 12597 15712 12631
rect 15660 12588 15712 12597
rect 17316 12631 17368 12640
rect 17316 12597 17325 12631
rect 17325 12597 17359 12631
rect 17359 12597 17368 12631
rect 17316 12588 17368 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1584 12384 1636 12436
rect 2044 12384 2096 12436
rect 2780 12384 2832 12436
rect 5448 12384 5500 12436
rect 6368 12384 6420 12436
rect 7840 12427 7892 12436
rect 7840 12393 7849 12427
rect 7849 12393 7883 12427
rect 7883 12393 7892 12427
rect 7840 12384 7892 12393
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 1952 12359 2004 12368
rect 1952 12325 1961 12359
rect 1961 12325 1995 12359
rect 1995 12325 2004 12359
rect 1952 12316 2004 12325
rect 2412 12359 2464 12368
rect 2412 12325 2421 12359
rect 2421 12325 2455 12359
rect 2455 12325 2464 12359
rect 2412 12316 2464 12325
rect 2872 12316 2924 12368
rect 5264 12316 5316 12368
rect 8852 12316 8904 12368
rect 8944 12316 8996 12368
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 4344 12248 4396 12300
rect 5172 12248 5224 12300
rect 5540 12248 5592 12300
rect 6092 12248 6144 12300
rect 6644 12248 6696 12300
rect 8208 12248 8260 12300
rect 9956 12248 10008 12300
rect 10784 12316 10836 12368
rect 15660 12384 15712 12436
rect 16028 12384 16080 12436
rect 13176 12359 13228 12368
rect 13176 12325 13185 12359
rect 13185 12325 13219 12359
rect 13219 12325 13228 12359
rect 13176 12316 13228 12325
rect 13544 12359 13596 12368
rect 13544 12325 13553 12359
rect 13553 12325 13587 12359
rect 13587 12325 13596 12359
rect 13544 12316 13596 12325
rect 14372 12316 14424 12368
rect 15384 12316 15436 12368
rect 15568 12316 15620 12368
rect 11704 12248 11756 12300
rect 11796 12248 11848 12300
rect 18236 12248 18288 12300
rect 2504 12180 2556 12232
rect 4620 12223 4672 12232
rect 4620 12189 4629 12223
rect 4629 12189 4663 12223
rect 4663 12189 4672 12223
rect 4620 12180 4672 12189
rect 6000 12223 6052 12232
rect 6000 12189 6009 12223
rect 6009 12189 6043 12223
rect 6043 12189 6052 12223
rect 7564 12223 7616 12232
rect 6000 12180 6052 12189
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 9772 12180 9824 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14004 12223 14056 12232
rect 14004 12189 14013 12223
rect 14013 12189 14047 12223
rect 14047 12189 14056 12223
rect 14004 12180 14056 12189
rect 14740 12180 14792 12232
rect 6552 12112 6604 12164
rect 9588 12112 9640 12164
rect 14280 12112 14332 12164
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 4804 12044 4856 12096
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 6184 12044 6236 12096
rect 6644 12087 6696 12096
rect 6644 12053 6653 12087
rect 6653 12053 6687 12087
rect 6687 12053 6696 12087
rect 6644 12044 6696 12053
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7472 12087 7524 12096
rect 7472 12053 7481 12087
rect 7481 12053 7515 12087
rect 7515 12053 7524 12087
rect 7472 12044 7524 12053
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 9404 12087 9456 12096
rect 9404 12053 9413 12087
rect 9413 12053 9447 12087
rect 9447 12053 9456 12087
rect 9404 12044 9456 12053
rect 9680 12044 9732 12096
rect 10140 12087 10192 12096
rect 10140 12053 10149 12087
rect 10149 12053 10183 12087
rect 10183 12053 10192 12087
rect 10140 12044 10192 12053
rect 15476 12112 15528 12164
rect 17316 12112 17368 12164
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2688 11840 2740 11892
rect 3332 11840 3384 11892
rect 4068 11840 4120 11892
rect 4252 11840 4304 11892
rect 2872 11772 2924 11824
rect 3792 11772 3844 11824
rect 1952 11704 2004 11756
rect 3424 11704 3476 11756
rect 6000 11840 6052 11892
rect 6276 11840 6328 11892
rect 7564 11840 7616 11892
rect 8484 11840 8536 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 9588 11883 9640 11892
rect 9588 11849 9597 11883
rect 9597 11849 9631 11883
rect 9631 11849 9640 11883
rect 9588 11840 9640 11849
rect 11796 11840 11848 11892
rect 12900 11883 12952 11892
rect 12900 11849 12909 11883
rect 12909 11849 12943 11883
rect 12943 11849 12952 11883
rect 12900 11840 12952 11849
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 15292 11840 15344 11892
rect 6184 11815 6236 11824
rect 6184 11781 6193 11815
rect 6193 11781 6227 11815
rect 6227 11781 6236 11815
rect 6184 11772 6236 11781
rect 7472 11772 7524 11824
rect 8392 11815 8444 11824
rect 8392 11781 8401 11815
rect 8401 11781 8435 11815
rect 8435 11781 8444 11815
rect 8392 11772 8444 11781
rect 8852 11772 8904 11824
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 7932 11704 7984 11756
rect 1584 11611 1636 11620
rect 1584 11577 1593 11611
rect 1593 11577 1627 11611
rect 1627 11577 1636 11611
rect 1584 11568 1636 11577
rect 3148 11568 3200 11620
rect 3332 11611 3384 11620
rect 3332 11577 3335 11611
rect 3335 11577 3369 11611
rect 3369 11577 3384 11611
rect 3332 11568 3384 11577
rect 4252 11568 4304 11620
rect 5172 11636 5224 11688
rect 6460 11636 6512 11688
rect 6644 11568 6696 11620
rect 7012 11636 7064 11688
rect 8024 11636 8076 11688
rect 9404 11636 9456 11688
rect 10048 11636 10100 11688
rect 14832 11772 14884 11824
rect 15476 11815 15528 11824
rect 15476 11781 15485 11815
rect 15485 11781 15519 11815
rect 15519 11781 15528 11815
rect 15476 11772 15528 11781
rect 11704 11704 11756 11756
rect 12900 11704 12952 11756
rect 10692 11636 10744 11688
rect 10876 11636 10928 11688
rect 11336 11636 11388 11688
rect 13176 11636 13228 11688
rect 8392 11568 8444 11620
rect 9588 11568 9640 11620
rect 9772 11568 9824 11620
rect 11520 11611 11572 11620
rect 11520 11577 11529 11611
rect 11529 11577 11563 11611
rect 11563 11577 11572 11611
rect 11520 11568 11572 11577
rect 2964 11500 3016 11552
rect 4804 11543 4856 11552
rect 4804 11509 4813 11543
rect 4813 11509 4847 11543
rect 4847 11509 4856 11543
rect 4804 11500 4856 11509
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8208 11500 8260 11552
rect 9680 11500 9732 11552
rect 12992 11568 13044 11620
rect 14740 11704 14792 11756
rect 15568 11704 15620 11756
rect 15200 11568 15252 11620
rect 27620 11636 27672 11688
rect 14188 11500 14240 11552
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 18236 11543 18288 11552
rect 18236 11509 18245 11543
rect 18245 11509 18279 11543
rect 18279 11509 18288 11543
rect 18236 11500 18288 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2412 11296 2464 11348
rect 3608 11296 3660 11348
rect 2504 11271 2556 11280
rect 2504 11237 2513 11271
rect 2513 11237 2547 11271
rect 2547 11237 2556 11271
rect 2504 11228 2556 11237
rect 2964 11228 3016 11280
rect 3148 11271 3200 11280
rect 3148 11237 3157 11271
rect 3157 11237 3191 11271
rect 3191 11237 3200 11271
rect 3148 11228 3200 11237
rect 3976 11228 4028 11280
rect 4252 11228 4304 11280
rect 5540 11228 5592 11280
rect 2320 11160 2372 11212
rect 4620 11160 4672 11212
rect 7472 11296 7524 11348
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 14188 11296 14240 11348
rect 15200 11296 15252 11348
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 9864 11228 9916 11280
rect 10140 11228 10192 11280
rect 11336 11271 11388 11280
rect 6092 11160 6144 11212
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 7012 11160 7064 11212
rect 7564 11160 7616 11212
rect 8668 11160 8720 11212
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 12348 11228 12400 11280
rect 12900 11228 12952 11280
rect 14372 11228 14424 11280
rect 11244 11160 11296 11212
rect 11520 11160 11572 11212
rect 12256 11160 12308 11212
rect 15752 11203 15804 11212
rect 4344 11092 4396 11144
rect 4436 11092 4488 11144
rect 8116 11092 8168 11144
rect 11704 11092 11756 11144
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 15844 11092 15896 11144
rect 6184 11024 6236 11076
rect 8392 11024 8444 11076
rect 1952 10999 2004 11008
rect 1952 10965 1961 10999
rect 1961 10965 1995 10999
rect 1995 10965 2004 10999
rect 1952 10956 2004 10965
rect 3700 10956 3752 11008
rect 3792 10956 3844 11008
rect 5172 10956 5224 11008
rect 7840 10956 7892 11008
rect 8484 10956 8536 11008
rect 9772 10956 9824 11008
rect 10048 10956 10100 11008
rect 13084 10999 13136 11008
rect 13084 10965 13093 10999
rect 13093 10965 13127 10999
rect 13127 10965 13136 10999
rect 13084 10956 13136 10965
rect 13728 10956 13780 11008
rect 14740 10956 14792 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4068 10752 4120 10804
rect 4252 10752 4304 10804
rect 4528 10795 4580 10804
rect 4528 10761 4537 10795
rect 4537 10761 4571 10795
rect 4571 10761 4580 10795
rect 4528 10752 4580 10761
rect 6368 10752 6420 10804
rect 7012 10752 7064 10804
rect 9404 10752 9456 10804
rect 10140 10752 10192 10804
rect 10692 10795 10744 10804
rect 10692 10761 10701 10795
rect 10701 10761 10735 10795
rect 10735 10761 10744 10795
rect 10692 10752 10744 10761
rect 12348 10752 12400 10804
rect 13084 10752 13136 10804
rect 13452 10752 13504 10804
rect 3608 10727 3660 10736
rect 3608 10693 3617 10727
rect 3617 10693 3651 10727
rect 3651 10693 3660 10727
rect 3608 10684 3660 10693
rect 3700 10684 3752 10736
rect 3424 10616 3476 10668
rect 6092 10616 6144 10668
rect 7196 10684 7248 10736
rect 8484 10727 8536 10736
rect 8484 10693 8493 10727
rect 8493 10693 8527 10727
rect 8527 10693 8536 10727
rect 8484 10684 8536 10693
rect 9680 10727 9732 10736
rect 4528 10548 4580 10600
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 7472 10616 7524 10668
rect 8116 10616 8168 10668
rect 8576 10659 8628 10668
rect 8576 10625 8582 10659
rect 8582 10625 8616 10659
rect 8616 10625 8628 10659
rect 9680 10693 9689 10727
rect 9689 10693 9723 10727
rect 9723 10693 9732 10727
rect 9680 10684 9732 10693
rect 13176 10727 13228 10736
rect 13176 10693 13185 10727
rect 13185 10693 13219 10727
rect 13219 10693 13228 10727
rect 13176 10684 13228 10693
rect 14096 10752 14148 10804
rect 15844 10795 15896 10804
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 19340 10752 19392 10804
rect 16948 10684 17000 10736
rect 8576 10616 8628 10625
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 2044 10412 2096 10464
rect 3056 10412 3108 10464
rect 6552 10480 6604 10532
rect 4528 10412 4580 10464
rect 7656 10412 7708 10464
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 9956 10616 10008 10668
rect 13360 10616 13412 10668
rect 9864 10548 9916 10600
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11244 10591 11296 10600
rect 11244 10557 11253 10591
rect 11253 10557 11287 10591
rect 11287 10557 11296 10591
rect 11244 10548 11296 10557
rect 14004 10591 14056 10600
rect 14004 10557 14013 10591
rect 14013 10557 14047 10591
rect 14047 10557 14056 10591
rect 14004 10548 14056 10557
rect 15292 10591 15344 10600
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 15752 10548 15804 10600
rect 23756 10591 23808 10600
rect 23756 10557 23774 10591
rect 23774 10557 23808 10591
rect 8944 10523 8996 10532
rect 8944 10489 8953 10523
rect 8953 10489 8987 10523
rect 8987 10489 8996 10523
rect 8944 10480 8996 10489
rect 11520 10523 11572 10532
rect 11520 10489 11529 10523
rect 11529 10489 11563 10523
rect 11563 10489 11572 10523
rect 11520 10480 11572 10489
rect 13360 10523 13412 10532
rect 13360 10489 13369 10523
rect 13369 10489 13403 10523
rect 13403 10489 13412 10523
rect 13360 10480 13412 10489
rect 13452 10523 13504 10532
rect 13452 10489 13461 10523
rect 13461 10489 13495 10523
rect 13495 10489 13504 10523
rect 23756 10548 23808 10557
rect 13452 10480 13504 10489
rect 10968 10412 11020 10464
rect 14740 10412 14792 10464
rect 18144 10412 18196 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2228 10208 2280 10260
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 6460 10208 6512 10260
rect 1676 10140 1728 10192
rect 2964 10183 3016 10192
rect 2964 10149 2973 10183
rect 2973 10149 3007 10183
rect 3007 10149 3016 10183
rect 2964 10140 3016 10149
rect 7012 10183 7064 10192
rect 7012 10149 7021 10183
rect 7021 10149 7055 10183
rect 7055 10149 7064 10183
rect 8116 10208 8168 10260
rect 8576 10208 8628 10260
rect 8944 10208 8996 10260
rect 9496 10208 9548 10260
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 12348 10208 12400 10260
rect 7012 10140 7064 10149
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 4528 10072 4580 10124
rect 5172 10115 5224 10124
rect 1768 10004 1820 10056
rect 2320 10004 2372 10056
rect 3700 10047 3752 10056
rect 3700 10013 3709 10047
rect 3709 10013 3743 10047
rect 3743 10013 3752 10047
rect 3700 10004 3752 10013
rect 4804 10004 4856 10056
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 10968 10140 11020 10192
rect 8392 10072 8444 10124
rect 10140 10072 10192 10124
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 12808 10072 12860 10124
rect 14464 10140 14516 10192
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 7288 10004 7340 10056
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 2596 9936 2648 9988
rect 4620 9936 4672 9988
rect 8484 9936 8536 9988
rect 9680 9936 9732 9988
rect 18236 10004 18288 10056
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 8392 9868 8444 9920
rect 9864 9911 9916 9920
rect 9864 9877 9888 9911
rect 9888 9877 9916 9911
rect 9864 9868 9916 9877
rect 11152 9868 11204 9920
rect 15292 9868 15344 9920
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1676 9707 1728 9716
rect 1676 9673 1685 9707
rect 1685 9673 1719 9707
rect 1719 9673 1728 9707
rect 1676 9664 1728 9673
rect 3240 9664 3292 9716
rect 2688 9528 2740 9580
rect 6184 9664 6236 9716
rect 6552 9707 6604 9716
rect 6552 9673 6561 9707
rect 6561 9673 6595 9707
rect 6595 9673 6604 9707
rect 6552 9664 6604 9673
rect 7564 9664 7616 9716
rect 8392 9664 8444 9716
rect 10876 9664 10928 9716
rect 13268 9664 13320 9716
rect 5172 9596 5224 9648
rect 7748 9596 7800 9648
rect 11336 9596 11388 9648
rect 12900 9639 12952 9648
rect 12900 9605 12909 9639
rect 12909 9605 12943 9639
rect 12943 9605 12952 9639
rect 12900 9596 12952 9605
rect 6092 9528 6144 9580
rect 6552 9460 6604 9512
rect 1860 9392 1912 9444
rect 4896 9435 4948 9444
rect 4896 9401 4905 9435
rect 4905 9401 4939 9435
rect 4939 9401 4948 9435
rect 4896 9392 4948 9401
rect 6736 9392 6788 9444
rect 8024 9460 8076 9512
rect 9036 9528 9088 9580
rect 10784 9528 10836 9580
rect 15384 9664 15436 9716
rect 15936 9664 15988 9716
rect 14648 9528 14700 9580
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 9772 9435 9824 9444
rect 9772 9401 9781 9435
rect 9781 9401 9815 9435
rect 9815 9401 9824 9435
rect 9772 9392 9824 9401
rect 2044 9324 2096 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 7656 9324 7708 9376
rect 7932 9324 7984 9376
rect 8392 9324 8444 9376
rect 9680 9324 9732 9376
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10876 9392 10928 9444
rect 11888 9392 11940 9444
rect 12900 9392 12952 9444
rect 16948 9392 17000 9444
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 4528 9120 4580 9172
rect 4804 9120 4856 9172
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 9036 9163 9088 9172
rect 9036 9129 9045 9163
rect 9045 9129 9079 9163
rect 9079 9129 9088 9163
rect 9036 9120 9088 9129
rect 11520 9120 11572 9172
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 15292 9120 15344 9172
rect 2044 9095 2096 9104
rect 2044 9061 2053 9095
rect 2053 9061 2087 9095
rect 2087 9061 2096 9095
rect 2044 9052 2096 9061
rect 2596 9095 2648 9104
rect 2596 9061 2605 9095
rect 2605 9061 2639 9095
rect 2639 9061 2648 9095
rect 2596 9052 2648 9061
rect 7196 9095 7248 9104
rect 7196 9061 7205 9095
rect 7205 9061 7239 9095
rect 7239 9061 7248 9095
rect 7196 9052 7248 9061
rect 11336 9095 11388 9104
rect 11336 9061 11345 9095
rect 11345 9061 11379 9095
rect 11379 9061 11388 9095
rect 11336 9052 11388 9061
rect 12900 9052 12952 9104
rect 15936 9120 15988 9172
rect 6276 8984 6328 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 7288 8984 7340 9036
rect 7932 8984 7984 9036
rect 8944 8984 8996 9036
rect 9496 8984 9548 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 16948 9027 17000 9036
rect 16948 8993 16957 9027
rect 16957 8993 16991 9027
rect 16991 8993 17000 9027
rect 16948 8984 17000 8993
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 4620 8916 4672 8968
rect 6920 8916 6972 8968
rect 9956 8916 10008 8968
rect 11612 8916 11664 8968
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 14740 8916 14792 8968
rect 15660 8916 15712 8968
rect 16120 8916 16172 8968
rect 16212 8916 16264 8968
rect 8668 8848 8720 8900
rect 10048 8848 10100 8900
rect 1768 8780 1820 8832
rect 3976 8780 4028 8832
rect 5540 8780 5592 8832
rect 7840 8780 7892 8832
rect 8024 8780 8076 8832
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 10784 8780 10836 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2320 8508 2372 8560
rect 4436 8508 4488 8560
rect 1952 8440 2004 8492
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 3976 8440 4028 8449
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 1860 8304 1912 8356
rect 2964 8304 3016 8356
rect 4068 8304 4120 8356
rect 5264 8576 5316 8628
rect 7748 8576 7800 8628
rect 6828 8508 6880 8560
rect 8208 8508 8260 8560
rect 9680 8576 9732 8628
rect 10048 8576 10100 8628
rect 12900 8576 12952 8628
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 9864 8508 9916 8560
rect 10508 8508 10560 8560
rect 5448 8440 5500 8492
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 13728 8440 13780 8492
rect 14372 8440 14424 8492
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 7840 8372 7892 8424
rect 5540 8304 5592 8356
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 5264 8236 5316 8288
rect 5908 8279 5960 8288
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 6276 8279 6328 8288
rect 6276 8245 6285 8279
rect 6285 8245 6319 8279
rect 6319 8245 6328 8279
rect 6276 8236 6328 8245
rect 6736 8304 6788 8356
rect 7288 8236 7340 8288
rect 8208 8279 8260 8288
rect 8208 8245 8217 8279
rect 8217 8245 8251 8279
rect 8251 8245 8260 8279
rect 10048 8304 10100 8356
rect 12900 8304 12952 8356
rect 8208 8236 8260 8245
rect 10692 8236 10744 8288
rect 11336 8236 11388 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 25136 8372 25188 8424
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 15844 8347 15896 8356
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 15844 8313 15853 8347
rect 15853 8313 15887 8347
rect 15887 8313 15896 8347
rect 15844 8304 15896 8313
rect 14096 8236 14148 8245
rect 15568 8236 15620 8288
rect 18604 8236 18656 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 2044 8032 2096 8084
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 4988 8032 5040 8084
rect 7288 8075 7340 8084
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 13084 8075 13136 8084
rect 13084 8041 13093 8075
rect 13093 8041 13127 8075
rect 13127 8041 13136 8075
rect 13084 8032 13136 8041
rect 15292 8032 15344 8084
rect 15844 8032 15896 8084
rect 1768 8007 1820 8016
rect 1768 7973 1777 8007
rect 1777 7973 1811 8007
rect 1811 7973 1820 8007
rect 1768 7964 1820 7973
rect 4804 7964 4856 8016
rect 5448 8007 5500 8016
rect 5448 7973 5457 8007
rect 5457 7973 5491 8007
rect 5491 7973 5500 8007
rect 5448 7964 5500 7973
rect 5908 7964 5960 8016
rect 6368 7964 6420 8016
rect 10048 7964 10100 8016
rect 12256 8007 12308 8016
rect 8576 7896 8628 7948
rect 9772 7896 9824 7948
rect 10968 7896 11020 7948
rect 12256 7973 12265 8007
rect 12265 7973 12299 8007
rect 12299 7973 12308 8007
rect 12256 7964 12308 7973
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 14372 8007 14424 8016
rect 13820 7964 13872 7973
rect 14372 7973 14381 8007
rect 14381 7973 14415 8007
rect 14415 7973 14424 8007
rect 14372 7964 14424 7973
rect 15384 7964 15436 8016
rect 16212 7964 16264 8016
rect 25504 7896 25556 7948
rect 1952 7871 2004 7880
rect 1584 7760 1636 7812
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 5080 7828 5132 7880
rect 6460 7828 6512 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 11888 7828 11940 7880
rect 12624 7828 12676 7880
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 15660 7871 15712 7880
rect 1860 7760 1912 7812
rect 2596 7760 2648 7812
rect 3700 7760 3752 7812
rect 5448 7760 5500 7812
rect 15660 7837 15669 7871
rect 15669 7837 15703 7871
rect 15703 7837 15712 7871
rect 15660 7828 15712 7837
rect 16212 7692 16264 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 6092 7531 6144 7540
rect 6092 7497 6101 7531
rect 6101 7497 6135 7531
rect 6135 7497 6144 7531
rect 6092 7488 6144 7497
rect 6368 7531 6420 7540
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 9128 7488 9180 7540
rect 10048 7488 10100 7540
rect 10876 7531 10928 7540
rect 6276 7420 6328 7472
rect 8576 7420 8628 7472
rect 1860 7352 1912 7404
rect 1952 7352 2004 7404
rect 7196 7352 7248 7404
rect 3148 7284 3200 7336
rect 4528 7284 4580 7336
rect 6092 7284 6144 7336
rect 7656 7284 7708 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 10876 7497 10885 7531
rect 10885 7497 10919 7531
rect 10919 7497 10928 7531
rect 10876 7488 10928 7497
rect 12256 7488 12308 7540
rect 15384 7531 15436 7540
rect 15384 7497 15393 7531
rect 15393 7497 15427 7531
rect 15427 7497 15436 7531
rect 15384 7488 15436 7497
rect 16212 7488 16264 7540
rect 10876 7352 10928 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 13820 7352 13872 7404
rect 24124 7352 24176 7404
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 16120 7284 16172 7336
rect 27620 7284 27672 7336
rect 3240 7259 3292 7268
rect 3240 7225 3249 7259
rect 3249 7225 3283 7259
rect 3283 7225 3292 7259
rect 3240 7216 3292 7225
rect 8668 7216 8720 7268
rect 12532 7259 12584 7268
rect 12532 7225 12541 7259
rect 12541 7225 12575 7259
rect 12575 7225 12584 7259
rect 12532 7216 12584 7225
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 4988 7148 5040 7200
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 12164 7191 12216 7200
rect 12164 7157 12173 7191
rect 12173 7157 12207 7191
rect 12207 7157 12216 7191
rect 12164 7148 12216 7157
rect 15844 7148 15896 7200
rect 25504 7191 25556 7200
rect 25504 7157 25513 7191
rect 25513 7157 25547 7191
rect 25547 7157 25556 7191
rect 25504 7148 25556 7157
rect 26516 7148 26568 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1768 6944 1820 6996
rect 3240 6944 3292 6996
rect 5080 6944 5132 6996
rect 6828 6944 6880 6996
rect 8116 6944 8168 6996
rect 9680 6944 9732 6996
rect 2964 6876 3016 6928
rect 4896 6876 4948 6928
rect 5172 6876 5224 6928
rect 9588 6876 9640 6928
rect 10692 6987 10744 6996
rect 10692 6953 10701 6987
rect 10701 6953 10735 6987
rect 10735 6953 10744 6987
rect 10692 6944 10744 6953
rect 10968 6987 11020 6996
rect 10968 6953 10977 6987
rect 10977 6953 11011 6987
rect 11011 6953 11020 6987
rect 10968 6944 11020 6953
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 12624 6944 12676 6996
rect 14096 6987 14148 6996
rect 14096 6953 14105 6987
rect 14105 6953 14139 6987
rect 14139 6953 14148 6987
rect 14096 6944 14148 6953
rect 12164 6919 12216 6928
rect 12164 6885 12173 6919
rect 12173 6885 12207 6919
rect 12207 6885 12216 6919
rect 12164 6876 12216 6885
rect 2320 6808 2372 6860
rect 6368 6808 6420 6860
rect 6644 6808 6696 6860
rect 6736 6808 6788 6860
rect 9772 6808 9824 6860
rect 12256 6808 12308 6860
rect 12808 6808 12860 6860
rect 15844 6851 15896 6860
rect 15844 6817 15853 6851
rect 15853 6817 15887 6851
rect 15887 6817 15896 6851
rect 15844 6808 15896 6817
rect 17040 6808 17092 6860
rect 7196 6740 7248 6792
rect 8484 6740 8536 6792
rect 13268 6740 13320 6792
rect 13728 6740 13780 6792
rect 6460 6672 6512 6724
rect 1860 6604 1912 6656
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 5356 6604 5408 6656
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 7748 6604 7800 6656
rect 8024 6604 8076 6656
rect 9220 6604 9272 6656
rect 13452 6604 13504 6656
rect 16672 6604 16724 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 6368 6400 6420 6452
rect 7196 6400 7248 6452
rect 7748 6400 7800 6452
rect 8116 6443 8168 6452
rect 8116 6409 8125 6443
rect 8125 6409 8159 6443
rect 8159 6409 8168 6443
rect 8116 6400 8168 6409
rect 11152 6400 11204 6452
rect 12256 6400 12308 6452
rect 12808 6400 12860 6452
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 9220 6375 9272 6384
rect 9220 6341 9229 6375
rect 9229 6341 9263 6375
rect 9263 6341 9272 6375
rect 9220 6332 9272 6341
rect 22928 6332 22980 6384
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 2228 6264 2280 6316
rect 3148 6264 3200 6316
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 6736 6264 6788 6316
rect 8668 6264 8720 6316
rect 12532 6264 12584 6316
rect 5540 6196 5592 6248
rect 20812 6239 20864 6248
rect 20812 6205 20821 6239
rect 20821 6205 20855 6239
rect 20855 6205 20864 6239
rect 20812 6196 20864 6205
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 1860 6171 1912 6180
rect 1860 6137 1869 6171
rect 1869 6137 1903 6171
rect 1903 6137 1912 6171
rect 1860 6128 1912 6137
rect 7656 6128 7708 6180
rect 8392 6128 8444 6180
rect 2964 6060 3016 6112
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 17040 6103 17092 6112
rect 17040 6069 17049 6103
rect 17049 6069 17083 6103
rect 17083 6069 17092 6103
rect 17040 6060 17092 6069
rect 18604 6060 18656 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1768 5856 1820 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 2228 5788 2280 5840
rect 2412 5788 2464 5840
rect 8484 5788 8536 5840
rect 4068 5720 4120 5772
rect 7196 5720 7248 5772
rect 7840 5720 7892 5772
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8300 5584 8352 5636
rect 7564 5516 7616 5568
rect 7932 5559 7984 5568
rect 7932 5525 7941 5559
rect 7941 5525 7975 5559
rect 7975 5525 7984 5559
rect 7932 5516 7984 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 6644 5312 6696 5364
rect 10140 5312 10192 5364
rect 4068 5287 4120 5296
rect 4068 5253 4077 5287
rect 4077 5253 4111 5287
rect 4111 5253 4120 5287
rect 4068 5244 4120 5253
rect 8024 5244 8076 5296
rect 9772 5244 9824 5296
rect 3056 5176 3108 5228
rect 1676 5108 1728 5160
rect 3792 5108 3844 5160
rect 1216 5040 1268 5092
rect 7288 5040 7340 5092
rect 8484 5083 8536 5092
rect 8484 5049 8493 5083
rect 8493 5049 8527 5083
rect 8527 5049 8536 5083
rect 8484 5040 8536 5049
rect 5172 4972 5224 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 9404 5015 9456 5024
rect 9404 4981 9413 5015
rect 9413 4981 9447 5015
rect 9447 4981 9456 5015
rect 9404 4972 9456 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1768 4768 1820 4820
rect 2596 4811 2648 4820
rect 2596 4777 2605 4811
rect 2605 4777 2639 4811
rect 2639 4777 2648 4811
rect 2596 4768 2648 4777
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 8484 4768 8536 4820
rect 10784 4700 10836 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 7288 4675 7340 4684
rect 7288 4641 7297 4675
rect 7297 4641 7331 4675
rect 7331 4641 7340 4675
rect 7288 4632 7340 4641
rect 7472 4632 7524 4684
rect 9404 4632 9456 4684
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 112 4224 164 4276
rect 2412 4267 2464 4276
rect 2412 4233 2421 4267
rect 2421 4233 2455 4267
rect 2455 4233 2464 4267
rect 2412 4224 2464 4233
rect 7380 4224 7432 4276
rect 1676 4156 1728 4208
rect 7472 4156 7524 4208
rect 10692 4088 10744 4140
rect 12348 4088 12400 4140
rect 1308 4020 1360 4072
rect 10784 3952 10836 4004
rect 11428 3884 11480 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1492 3680 1544 3732
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 11428 3612 11480 3664
rect 13360 3612 13412 3664
rect 13452 3587 13504 3596
rect 13452 3553 13461 3587
rect 13461 3553 13495 3587
rect 13495 3553 13504 3587
rect 13452 3544 13504 3553
rect 11520 3476 11572 3528
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3424 3136 3476 3188
rect 10876 3136 10928 3188
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 13360 3000 13412 3052
rect 112 2932 164 2984
rect 14464 2932 14516 2984
rect 10784 2839 10836 2848
rect 10784 2805 10793 2839
rect 10793 2805 10827 2839
rect 10827 2805 10836 2839
rect 10784 2796 10836 2805
rect 11520 2796 11572 2848
rect 12900 2864 12952 2916
rect 14004 2796 14056 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1768 2592 1820 2644
rect 4712 2592 4764 2644
rect 11520 2592 11572 2644
rect 12532 2592 12584 2644
rect 756 2388 808 2440
rect 9128 2456 9180 2508
rect 6644 2252 6696 2304
rect 14004 2456 14056 2508
rect 12532 2252 12584 2304
rect 14556 2252 14608 2304
rect 16028 2252 16080 2304
rect 20628 2252 20680 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 23756 76 23808 128
rect 24860 76 24912 128
<< metal2 >>
rect 938 27520 994 28000
rect 2870 27520 2926 28000
rect 4894 27520 4950 28000
rect 6918 27520 6974 28000
rect 8850 27520 8906 28000
rect 10874 27520 10930 28000
rect 12898 27554 12954 28000
rect 12728 27526 12954 27554
rect 110 24576 166 24585
rect 110 24511 166 24520
rect 124 23186 152 24511
rect 112 23180 164 23186
rect 112 23122 164 23128
rect 952 19378 980 27520
rect 2502 26752 2558 26761
rect 2502 26687 2558 26696
rect 1306 25392 1362 25401
rect 1306 25327 1362 25336
rect 1320 23730 1348 25327
rect 1308 23724 1360 23730
rect 1308 23666 1360 23672
rect 1124 23520 1176 23526
rect 1124 23462 1176 23468
rect 940 19372 992 19378
rect 940 19314 992 19320
rect 1136 15706 1164 23462
rect 1214 22672 1270 22681
rect 1214 22607 1270 22616
rect 1228 22166 1256 22607
rect 1216 22160 1268 22166
rect 1216 22102 1268 22108
rect 1228 21690 1256 22102
rect 1216 21684 1268 21690
rect 1216 21626 1268 21632
rect 1582 21312 1638 21321
rect 1582 21247 1638 21256
rect 1596 20602 1624 21247
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1582 20088 1638 20097
rect 1582 20023 1638 20032
rect 1596 18970 1624 20023
rect 1688 19514 1716 20334
rect 1952 20052 2004 20058
rect 1872 20012 1952 20040
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1872 19334 1900 20012
rect 1952 19994 2004 20000
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 1780 19306 1900 19334
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1780 18834 1808 19306
rect 1964 19174 1992 19858
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1582 18728 1638 18737
rect 1582 18663 1638 18672
rect 1596 18426 1624 18663
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17134 1532 17478
rect 1492 17128 1544 17134
rect 1492 17070 1544 17076
rect 1124 15700 1176 15706
rect 1124 15642 1176 15648
rect 1504 13462 1532 17070
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 15910 1624 16594
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1596 15745 1624 15846
rect 1582 15736 1638 15745
rect 1582 15671 1638 15680
rect 1688 15026 1716 16390
rect 1766 16008 1822 16017
rect 1766 15943 1822 15952
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1688 13938 1716 14486
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1688 13530 1716 13738
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 1780 12986 1808 15943
rect 1872 13802 1900 16934
rect 1964 16561 1992 19110
rect 2056 18426 2084 19654
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 18426 2360 18770
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2320 18420 2372 18426
rect 2320 18362 2372 18368
rect 2056 18222 2084 18362
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16046 1992 16390
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 14890 1992 15982
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1964 14618 1992 14826
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1952 13456 2004 13462
rect 1952 13398 2004 13404
rect 1964 12986 1992 13398
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1780 12782 1808 12922
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1596 11626 1624 12378
rect 1964 12374 1992 12922
rect 2056 12442 2084 17478
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2148 15638 2176 15846
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 2148 15162 2176 15574
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2240 14550 2268 15914
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2240 13530 2268 14350
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2228 13524 2280 13530
rect 2228 13466 2280 13472
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1952 12368 2004 12374
rect 1952 12310 2004 12316
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1584 11620 1636 11626
rect 1584 11562 1636 11568
rect 1964 11014 1992 11698
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 1688 10198 1716 10406
rect 1676 10192 1728 10198
rect 1676 10134 1728 10140
rect 1688 9722 1716 10134
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1490 9344 1546 9353
rect 1490 9279 1546 9288
rect 1306 7984 1362 7993
rect 1306 7919 1362 7928
rect 1216 5092 1268 5098
rect 1216 5034 1268 5040
rect 110 4584 166 4593
rect 110 4519 166 4528
rect 124 4282 152 4519
rect 112 4276 164 4282
rect 112 4218 164 4224
rect 110 3224 166 3233
rect 110 3159 166 3168
rect 124 2990 152 3159
rect 112 2984 164 2990
rect 112 2926 164 2932
rect 756 2440 808 2446
rect 756 2382 808 2388
rect 768 2281 796 2382
rect 754 2272 810 2281
rect 754 2207 810 2216
rect 938 82 994 480
rect 1228 82 1256 5034
rect 1320 4078 1348 7919
rect 1400 4684 1452 4690
rect 1504 4672 1532 9279
rect 1780 8838 1808 9998
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1872 8362 1900 9386
rect 2056 9382 2084 10406
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9110 2084 9318
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1964 8498 1992 8910
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1584 7812 1636 7818
rect 1584 7754 1636 7760
rect 1452 4644 1532 4672
rect 1400 4626 1452 4632
rect 1308 4072 1360 4078
rect 1308 4014 1360 4020
rect 1504 3738 1532 4644
rect 1596 4196 1624 7754
rect 1780 7002 1808 7958
rect 1964 7886 1992 8434
rect 2056 8090 2084 9046
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7410 1900 7754
rect 1964 7410 1992 7822
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1674 6760 1730 6769
rect 1674 6695 1730 6704
rect 1688 5166 1716 6695
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6186 1900 6598
rect 2148 6322 2176 13262
rect 2332 12918 2360 14010
rect 2424 13920 2452 19110
rect 2516 18222 2544 26687
rect 2884 19514 2912 27520
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 3240 22976 3292 22982
rect 3240 22918 3292 22924
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2884 19310 2912 19450
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2976 18737 3004 19110
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2962 18728 3018 18737
rect 2962 18663 3018 18672
rect 3068 18426 3096 18770
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2884 16998 2912 17682
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2596 15428 2648 15434
rect 2596 15370 2648 15376
rect 2608 15026 2636 15370
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2608 14074 2636 14486
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2424 13892 2636 13920
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2320 12912 2372 12918
rect 2320 12854 2372 12860
rect 2332 12714 2360 12854
rect 2424 12782 2452 13194
rect 2412 12776 2464 12782
rect 2412 12718 2464 12724
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2424 11354 2452 12310
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2516 11286 2544 12174
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2240 8430 2268 10202
rect 2332 10062 2360 11154
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2608 9994 2636 13892
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2700 13462 2728 13806
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2700 11898 2728 12650
rect 2792 12442 2820 16390
rect 2884 13814 2912 16934
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2976 16250 3004 16594
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2976 15162 3004 16186
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2884 13786 3004 13814
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12753 2912 12786
rect 2870 12744 2926 12753
rect 2870 12679 2926 12688
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2884 11830 2912 12310
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2976 11558 3004 13786
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11286 3004 11494
rect 3160 11286 3188 11562
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2976 10198 3004 11222
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 9110 2636 9930
rect 2700 9586 2728 10066
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2332 6866 2360 8502
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 1780 5914 1808 6122
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 2148 5710 2176 6258
rect 2240 5846 2268 6258
rect 2228 5840 2280 5846
rect 2332 5828 2360 6802
rect 2412 5840 2464 5846
rect 2332 5800 2412 5828
rect 2228 5782 2280 5788
rect 2412 5782 2464 5788
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1780 4826 1808 5646
rect 2240 5370 2268 5782
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2608 4826 2636 7754
rect 2976 6934 3004 8298
rect 2964 6928 3016 6934
rect 2964 6870 3016 6876
rect 2976 6118 3004 6870
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 1676 4208 1728 4214
rect 1596 4168 1676 4196
rect 1676 4150 1728 4156
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1780 2650 1808 4762
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2424 4282 2452 4626
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 938 54 1256 82
rect 2870 82 2926 480
rect 2976 82 3004 6054
rect 3068 5370 3096 10406
rect 3252 9722 3280 22918
rect 4080 22778 4108 23122
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4908 22098 4936 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6932 23866 6960 27520
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 4528 22092 4580 22098
rect 4528 22034 4580 22040
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4540 21690 4568 22034
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 5276 21554 5304 21830
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3436 19174 3464 19858
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3436 13870 3464 19110
rect 3606 17368 3662 17377
rect 3606 17303 3662 17312
rect 3620 16658 3648 17303
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3712 16794 3740 17070
rect 3896 17066 3924 19654
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3344 11626 3372 11834
rect 3436 11762 3464 12038
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3436 9926 3464 10610
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3436 9625 3464 9862
rect 3422 9616 3478 9625
rect 3422 9551 3478 9560
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 7546 3188 8230
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3160 7342 3188 7482
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 7002 3280 7210
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3160 6322 3188 6598
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 5137 3096 5170
rect 3054 5128 3110 5137
rect 3054 5063 3110 5072
rect 3528 4154 3556 16458
rect 3620 16250 3648 16594
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3712 14618 3740 14962
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3804 14618 3832 14826
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3896 13814 3924 17002
rect 3988 15706 4016 20878
rect 4712 20528 4764 20534
rect 4712 20470 4764 20476
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4344 19372 4396 19378
rect 4068 19346 4120 19352
rect 4344 19314 4396 19320
rect 4068 19288 4120 19294
rect 4160 19304 4212 19310
rect 4080 19174 4108 19288
rect 4160 19246 4212 19252
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4172 18426 4200 19246
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4356 18358 4384 19314
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4448 19174 4476 19246
rect 4632 19174 4660 19858
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4344 18352 4396 18358
rect 4344 18294 4396 18300
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4264 18086 4292 18158
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4264 17746 4292 18022
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4172 15026 4200 17478
rect 4264 16998 4292 17682
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16046 4292 16934
rect 4356 16658 4384 17002
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4252 16040 4304 16046
rect 4252 15982 4304 15988
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3988 14074 4016 14486
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4080 13938 4108 14350
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3896 13786 4016 13814
rect 3884 13728 3936 13734
rect 3804 13705 3884 13716
rect 3790 13696 3884 13705
rect 3846 13688 3884 13696
rect 3884 13670 3936 13676
rect 3790 13631 3846 13640
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12889 3740 13126
rect 3698 12880 3754 12889
rect 3698 12815 3754 12824
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3620 10742 3648 11290
rect 3804 11014 3832 11766
rect 3988 11286 4016 13786
rect 4172 13394 4200 14962
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4264 13870 4292 14350
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4172 12918 4200 13330
rect 4160 12912 4212 12918
rect 4080 12860 4160 12866
rect 4080 12854 4212 12860
rect 4080 12838 4200 12854
rect 4080 12306 4108 12838
rect 4172 12789 4200 12838
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4080 11898 4108 12242
rect 4264 11898 4292 13806
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4264 11286 4292 11562
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4252 11280 4304 11286
rect 4252 11222 4304 11228
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3712 10742 3740 10950
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3700 10736 3752 10742
rect 3700 10678 3752 10684
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3712 7818 3740 9998
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3804 5166 3832 10950
rect 4264 10810 4292 11222
rect 4356 11150 4384 12242
rect 4448 11234 4476 19110
rect 4632 18086 4660 19110
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 15638 4660 16526
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4632 15162 4660 15574
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4540 13530 4568 13806
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4540 13394 4568 13466
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4540 12986 4568 13330
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4448 11206 4568 11234
rect 4632 11218 4660 12174
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3988 8498 4016 8774
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4080 8362 4108 10746
rect 4448 8566 4476 11086
rect 4540 10810 4568 11206
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4540 10606 4568 10746
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4540 10130 4568 10406
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4632 9994 4660 11154
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4540 7342 4568 9114
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8090 4660 8910
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4080 5409 4108 5714
rect 4066 5400 4122 5409
rect 4066 5335 4122 5344
rect 4080 5302 4108 5335
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3436 4126 3556 4154
rect 3436 3194 3464 4126
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4724 2650 4752 20470
rect 5000 20466 5028 21286
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5184 20534 5212 20742
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5368 20058 5396 20266
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5460 19938 5488 23462
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7484 22166 7512 22374
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6932 21554 6960 21898
rect 7484 21690 7512 22102
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 5552 20942 5580 21490
rect 6932 21146 6960 21490
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 7024 21078 7052 21354
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 5540 20936 5592 20942
rect 5540 20878 5592 20884
rect 5552 20602 5580 20878
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6288 20602 6316 21014
rect 7576 21010 7604 21898
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 7760 20602 7788 22510
rect 8312 22438 8340 23122
rect 8864 22778 8892 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9864 23180 9916 23186
rect 9864 23122 9916 23128
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8220 21690 8248 21966
rect 8312 21962 8340 22374
rect 9232 22001 9260 22918
rect 9324 22778 9352 22918
rect 9876 22778 9904 23122
rect 10152 22982 10180 24142
rect 10888 23866 10916 27520
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 11060 23656 11112 23662
rect 11060 23598 11112 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10876 23248 10928 23254
rect 10876 23190 10928 23196
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9324 22574 9352 22714
rect 9312 22568 9364 22574
rect 9312 22510 9364 22516
rect 9218 21992 9274 22001
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8484 21956 8536 21962
rect 9218 21927 9274 21936
rect 8484 21898 8536 21904
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8496 21554 8524 21898
rect 9876 21554 9904 22714
rect 10428 22642 10456 22918
rect 10416 22636 10468 22642
rect 10416 22578 10468 22584
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22166 10180 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10796 22234 10824 23054
rect 10888 22438 10916 23190
rect 11072 23118 11100 23598
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12440 23248 12492 23254
rect 12440 23190 12492 23196
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22642 11100 23054
rect 12452 22778 12480 23190
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10876 22432 10928 22438
rect 10876 22374 10928 22380
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 10784 22228 10836 22234
rect 10784 22170 10836 22176
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10888 22098 10916 22374
rect 12360 22098 12388 22374
rect 12452 22166 12480 22714
rect 12544 22642 12572 23462
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12544 22216 12572 22578
rect 12624 22228 12676 22234
rect 12544 22188 12624 22216
rect 12624 22170 12676 22176
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 10876 22092 10928 22098
rect 10876 22034 10928 22040
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 10888 21690 10916 22034
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 8576 21412 8628 21418
rect 8576 21354 8628 21360
rect 8588 21146 8616 21354
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6288 19990 6316 20198
rect 6276 19984 6328 19990
rect 5460 19910 5580 19938
rect 6276 19926 6328 19932
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19446 5212 19654
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 5184 19310 5212 19382
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4816 18426 4844 19110
rect 5368 18970 5396 19178
rect 5460 18970 5488 19790
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4908 18426 4936 18770
rect 5552 18766 5580 19910
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6288 19514 6316 19926
rect 6748 19718 6776 20334
rect 7656 19984 7708 19990
rect 7656 19926 7708 19932
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6288 19174 6316 19450
rect 6748 19378 6776 19654
rect 7668 19514 7696 19926
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4896 18420 4948 18426
rect 4948 18380 5028 18408
rect 4896 18362 4948 18368
rect 4816 16028 4844 18362
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4908 17882 4936 18158
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 5000 17814 5028 18380
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 5092 16998 5120 18566
rect 5552 17882 5580 18702
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18426 6040 18838
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6196 18290 6224 18702
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 6196 17814 6224 18226
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 6184 17808 6236 17814
rect 6184 17750 6236 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4896 16040 4948 16046
rect 4816 16000 4896 16028
rect 4896 15982 4948 15988
rect 4908 15638 4936 15982
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 5092 13814 5120 16934
rect 5184 16794 5212 17614
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17134 5304 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6012 17338 6040 17750
rect 6288 17338 6316 19110
rect 6932 18970 6960 19110
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7300 18630 7328 19246
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6656 18086 6684 18158
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6656 17338 6684 18022
rect 7116 17338 7144 18090
rect 7484 17882 7512 18702
rect 7576 18358 7604 18838
rect 7760 18766 7788 20334
rect 8312 20058 8340 20946
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8036 18816 8064 19314
rect 8220 19174 8248 19790
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8116 18828 8168 18834
rect 8036 18788 8116 18816
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 7760 18290 7788 18702
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 6012 16794 6040 17274
rect 6092 17060 6144 17066
rect 6092 17002 6144 17008
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5184 16522 5212 16730
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5172 16516 5224 16522
rect 5172 16458 5224 16464
rect 5368 16250 5396 16662
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5460 15706 5488 16594
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6104 16017 6132 17002
rect 6288 16726 6316 17274
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6840 16794 6868 17070
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 6090 16008 6146 16017
rect 6090 15943 6146 15952
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5184 15094 5212 15438
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5184 14385 5212 15030
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5276 14618 5304 14962
rect 5368 14890 5396 15438
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 6012 14482 6040 14894
rect 6276 14884 6328 14890
rect 6276 14826 6328 14832
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5170 14376 5226 14385
rect 5170 14311 5226 14320
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13870 5580 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 14074 6040 14418
rect 6288 14074 6316 14826
rect 6380 14618 6408 15506
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6380 14074 6408 14554
rect 6564 14550 6592 16662
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15026 6868 15846
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 5540 13864 5592 13870
rect 5092 13786 5212 13814
rect 5540 13806 5592 13812
rect 6288 13814 6316 14010
rect 6564 14006 6592 14486
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6288 13786 6408 13814
rect 6564 13802 6592 13942
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 5000 12646 5028 13194
rect 5184 12782 5212 13786
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5172 12776 5224 12782
rect 5448 12776 5500 12782
rect 5224 12736 5304 12764
rect 5172 12718 5224 12724
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5276 12374 5304 12736
rect 5448 12718 5500 12724
rect 5460 12442 5488 12718
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 6104 12306 6132 13398
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6288 13190 6316 13330
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5184 12102 5212 12242
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4816 11558 4844 12038
rect 5184 11694 5212 12038
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 5552 11286 5580 12242
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11898 6040 12174
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6196 11830 6224 12038
rect 6288 11898 6316 13126
rect 6380 12986 6408 13786
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6748 13462 6776 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6840 13938 6868 14554
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6656 12646 6684 13330
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 12782 7052 13126
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 5540 11280 5592 11286
rect 5368 11240 5540 11268
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 10606 5212 10950
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10130 5212 10542
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4816 9178 4844 9998
rect 5184 9654 5212 10066
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4816 7206 4844 7958
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 6322 4844 7142
rect 4908 6934 4936 9386
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5000 8090 5028 8366
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5000 7206 5028 8026
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5092 7002 5120 7822
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5184 6934 5212 9590
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5276 8634 5304 9114
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5276 8294 5304 8570
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 5172 6928 5224 6934
rect 5172 6870 5224 6876
rect 5368 6662 5396 11240
rect 5540 11222 5592 11228
rect 6380 11218 6408 12378
rect 6656 12306 6684 12582
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6550 12200 6606 12209
rect 6550 12135 6552 12144
rect 6604 12135 6606 12144
rect 6552 12106 6604 12112
rect 6564 11762 6592 12106
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6104 10674 6132 11154
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6196 10130 6224 11018
rect 6380 10810 6408 11154
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6366 10704 6422 10713
rect 6366 10639 6422 10648
rect 6380 10266 6408 10639
rect 6472 10266 6500 11630
rect 6656 11626 6684 12038
rect 7024 11694 7052 12038
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 7024 11218 7052 11630
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7024 10810 7052 11154
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6196 9722 6224 10066
rect 6564 9722 6592 10474
rect 7024 10198 7052 10746
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5460 8022 5488 8434
rect 5552 8362 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5460 7818 5488 7958
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 5552 6254 5580 8298
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 8022 5948 8230
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6104 7546 6132 9522
rect 6564 9518 6592 9658
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8294 6316 8978
rect 6748 8362 6776 9386
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8566 6868 8978
rect 6932 8974 6960 9318
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6104 7342 6132 7482
rect 6288 7478 6316 8230
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6380 7546 6408 7958
rect 6748 7886 6776 8298
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6380 6866 6408 7482
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6380 6458 6408 6802
rect 6472 6730 6500 7822
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 7002 6868 7142
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 6656 6118 6684 6802
rect 6748 6662 6776 6802
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6322 6776 6598
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6656 5370 6684 6054
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 2870 54 3004 82
rect 4894 82 4950 480
rect 5184 82 5212 4966
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 7116 4154 7144 16390
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7208 9110 7236 10678
rect 7300 10062 7328 16934
rect 7484 16794 7512 17818
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7392 15570 7420 15914
rect 7380 15564 7432 15570
rect 7380 15506 7432 15512
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7392 14822 7420 15506
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 14958 7696 15302
rect 7760 15162 7788 15506
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7760 14958 7788 15098
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7668 14550 7696 14894
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13530 7420 13738
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7392 12918 7420 13262
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7484 12102 7512 12854
rect 7760 12714 7788 13126
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 12238 7604 12582
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11830 7512 12038
rect 7576 11898 7604 12174
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7484 11354 7512 11766
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7484 10062 7512 10610
rect 7576 10130 7604 11154
rect 7760 10996 7788 12650
rect 7852 12442 7880 18566
rect 8036 17746 8064 18788
rect 8116 18770 8168 18776
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 16998 8064 17682
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8220 15094 8248 19110
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8496 17746 8524 18838
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 16726 8340 17070
rect 8496 16998 8524 17682
rect 8680 17542 8708 18566
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8220 14822 8248 14894
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8404 14482 8432 14894
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8036 12850 8064 13194
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7944 11558 7972 11698
rect 8036 11694 8064 12786
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7840 11008 7892 11014
rect 7760 10968 7840 10996
rect 7840 10950 7892 10956
rect 7852 10470 7880 10950
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7208 7410 7236 9046
rect 7300 9042 7328 9998
rect 7576 9722 7604 10066
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7668 9674 7696 10406
rect 7944 10062 7972 11494
rect 8128 11150 8156 12922
rect 8312 12918 8340 13126
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8404 12850 8432 13670
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 12102 8248 12242
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11558 8248 12038
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10674 8156 11086
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10266 8156 10610
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7668 9654 7788 9674
rect 7668 9648 7800 9654
rect 7668 9646 7748 9648
rect 7748 9590 7800 9596
rect 7760 9500 7788 9590
rect 7576 9472 7788 9500
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 8090 7328 8230
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7208 6798 7236 7346
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7208 6458 7236 6734
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 4826 7236 5714
rect 7576 5574 7604 9472
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 7342 7696 9318
rect 7852 8838 7880 9862
rect 7944 9382 7972 9998
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9518 8064 9862
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7760 6662 7788 8570
rect 7944 8498 7972 8978
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7852 7886 7880 8366
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6458 7788 6598
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7300 4690 7328 5034
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7300 4264 7328 4626
rect 7380 4276 7432 4282
rect 7300 4236 7380 4264
rect 7380 4218 7432 4224
rect 7484 4214 7512 4626
rect 7668 4622 7696 6122
rect 7852 5778 7880 7822
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7944 5692 7972 7278
rect 8036 6662 8064 8774
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8220 8294 8248 8502
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8128 6458 8156 6938
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8024 5704 8076 5710
rect 7944 5664 8024 5692
rect 8024 5646 8076 5652
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5030 7972 5510
rect 8036 5302 8064 5646
rect 8220 5624 8248 8230
rect 8312 5914 8340 12718
rect 8404 12646 8432 12786
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8496 11898 8524 16934
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8588 13258 8616 13874
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8680 12986 8708 17478
rect 8772 17066 8800 18226
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8772 16726 8800 17002
rect 8760 16720 8812 16726
rect 8760 16662 8812 16668
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8772 15570 8800 15982
rect 9140 15638 9168 21490
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 20482 10732 21354
rect 10888 20534 10916 21626
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 20874 11008 21490
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11992 21010 12020 21354
rect 12360 21350 12388 22034
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 11256 20534 11284 20878
rect 11348 20602 11376 20878
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11992 20534 12020 20946
rect 10876 20528 10928 20534
rect 10704 20466 10824 20482
rect 10876 20470 10928 20476
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 10704 20460 10836 20466
rect 10704 20454 10784 20460
rect 10784 20402 10836 20408
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9312 19304 9364 19310
rect 9416 19281 9444 20198
rect 9876 19990 9904 20266
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9692 19378 9720 19790
rect 9876 19514 9904 19926
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9312 19246 9364 19252
rect 9402 19272 9458 19281
rect 9324 18766 9352 19246
rect 9402 19207 9458 19216
rect 9692 18970 9720 19314
rect 10704 19174 10732 20334
rect 11992 20058 12020 20470
rect 12360 20058 12388 21286
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11440 19514 11468 19926
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 10888 18902 10916 19246
rect 11440 18902 11468 19450
rect 11716 19174 11744 19790
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9876 18426 9904 18770
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 10520 18154 10548 18634
rect 11440 18426 11468 18838
rect 11428 18420 11480 18426
rect 11428 18362 11480 18368
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 10048 18148 10100 18154
rect 10048 18090 10100 18096
rect 10508 18148 10560 18154
rect 10508 18090 10560 18096
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 9232 17202 9260 18090
rect 10060 17814 10088 18090
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 17814 10180 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10336 17338 10364 17682
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9600 16114 9628 16662
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16250 9720 16526
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9876 16182 9904 17070
rect 10980 17066 11008 17274
rect 11164 17202 11192 18090
rect 11716 17678 11744 19110
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11808 18426 11836 18702
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17746 11928 18022
rect 12728 17882 12756 27526
rect 12898 27520 12954 27526
rect 14922 27520 14978 28000
rect 16854 27520 16910 28000
rect 18878 27520 18934 28000
rect 20902 27554 20958 28000
rect 20732 27526 20958 27554
rect 14936 26738 14964 27520
rect 14844 26710 14964 26738
rect 14844 23866 14872 26710
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 16868 23866 16896 27520
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 14372 23520 14424 23526
rect 14372 23462 14424 23468
rect 13452 23112 13504 23118
rect 13452 23054 13504 23060
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12820 22642 12848 22986
rect 13464 22778 13492 23054
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 13464 22545 13492 22714
rect 13450 22536 13506 22545
rect 13450 22471 13506 22480
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20466 12940 20742
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 12912 20369 12940 20402
rect 12898 20360 12954 20369
rect 12898 20295 12954 20304
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 13004 19990 13032 20266
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12820 19242 12848 19654
rect 13188 19378 13216 20402
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13740 19514 13768 19858
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13740 19242 13768 19450
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 12820 18329 12848 19178
rect 12912 18970 12940 19178
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 12990 18728 13046 18737
rect 12990 18663 13046 18672
rect 12806 18320 12862 18329
rect 12806 18255 12862 18264
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 13004 17814 13032 18663
rect 13188 18426 13216 18770
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13188 17814 13216 18362
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11900 17338 11928 17682
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 12544 17134 12572 17478
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10888 16726 10916 17002
rect 10980 16794 11008 17002
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 12176 16726 12204 16934
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 11980 16584 12032 16590
rect 11518 16552 11574 16561
rect 11980 16526 12032 16532
rect 11518 16487 11574 16496
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15638 9628 16050
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9128 15632 9180 15638
rect 9128 15574 9180 15580
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 8760 15564 8812 15570
rect 8760 15506 8812 15512
rect 8772 15162 8800 15506
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8772 14958 8800 15098
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 9140 14890 9168 15574
rect 9876 15366 9904 15982
rect 10152 15706 10180 15982
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8772 14278 8800 14486
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13802 8800 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8772 12986 8800 13738
rect 8864 13190 8892 13942
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8392 11824 8444 11830
rect 8588 11778 8616 12786
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8680 12102 8708 12650
rect 8956 12374 8984 14758
rect 9218 14512 9274 14521
rect 9218 14447 9274 14456
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 14074 9076 14214
rect 9232 14074 9260 14447
rect 9508 14278 9536 14826
rect 9876 14414 9904 15302
rect 10336 15162 10364 15506
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 11256 15026 11284 15438
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11440 14822 11468 15574
rect 11532 15502 11560 16487
rect 11992 16250 12020 16526
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12176 15978 12204 16662
rect 12544 16590 12572 17070
rect 13004 16658 13032 17750
rect 13188 17270 13216 17750
rect 13464 17338 13492 18022
rect 13832 17338 13860 18702
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 14016 17542 14044 18090
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 13188 16794 13216 17206
rect 14016 17202 14044 17478
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13556 15978 13584 16050
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 15094 11560 15438
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 11440 14550 11468 14758
rect 12544 14618 12572 14826
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9876 13938 9904 14350
rect 10796 14006 10824 14486
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9048 12850 9076 13126
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9140 12646 9168 13194
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8444 11772 8616 11778
rect 8392 11766 8616 11772
rect 8404 11750 8616 11766
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8404 11082 8432 11562
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8404 10130 8432 11018
rect 8496 11014 8524 11750
rect 8680 11218 8708 12038
rect 8864 11830 8892 12310
rect 9140 12209 9168 12582
rect 9126 12200 9182 12209
rect 9600 12170 9628 12854
rect 9692 12714 9720 13330
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 12918 9812 13194
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 12238 9812 12582
rect 9772 12232 9824 12238
rect 9678 12200 9734 12209
rect 9126 12135 9182 12144
rect 9588 12164 9640 12170
rect 9140 11898 9168 12135
rect 9772 12174 9824 12180
rect 9678 12135 9734 12144
rect 9588 12106 9640 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10742 8524 10950
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8496 9994 8524 10678
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10266 8616 10610
rect 8944 10532 8996 10538
rect 8944 10474 8996 10480
rect 8956 10266 8984 10474
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8404 9722 8432 9862
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8404 9382 8432 9658
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 6186 8432 9318
rect 8588 8106 8616 10202
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 9178 9076 9522
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8496 8078 8616 8106
rect 8496 6798 8524 8078
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7478 8616 7890
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8496 5846 8524 6734
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8300 5636 8352 5642
rect 8220 5596 8300 5624
rect 8300 5578 8352 5584
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 8312 4486 8340 5578
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8496 4826 8524 5034
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8588 4729 8616 7414
rect 8680 7274 8708 8842
rect 8956 8090 8984 8978
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9140 7546 9168 11834
rect 9416 11694 9444 12038
rect 9600 11898 9628 12106
rect 9692 12102 9720 12135
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 10810 9444 11630
rect 9784 11626 9812 12174
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9508 9518 9536 10202
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 9042 9536 9454
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8680 6322 8708 7210
rect 9600 6934 9628 11562
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 10742 9720 11494
rect 9876 11286 9904 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10796 13530 10824 13942
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 13530 11744 13738
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 10784 13524 10836 13530
rect 10704 13484 10784 13512
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9968 12306 9996 12922
rect 10704 12850 10732 13484
rect 10784 13466 10836 13472
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10060 12646 10088 12786
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10796 12374 10824 13262
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10888 12442 10916 12650
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9968 11354 9996 12242
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9772 11008 9824 11014
rect 9824 10968 9904 10996
rect 9772 10950 9824 10956
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9876 10606 9904 10968
rect 9968 10674 9996 11290
rect 10060 11014 10088 11630
rect 10152 11286 10180 12038
rect 10888 11694 10916 12378
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9382 9720 9930
rect 9876 9926 9904 10542
rect 10060 10062 10088 10950
rect 10152 10810 10180 11222
rect 10704 11218 10732 11630
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10704 10810 10732 11154
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9042 9720 9318
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8634 9720 8978
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9692 7002 9720 8570
rect 9784 7954 9812 9386
rect 9876 8566 9904 9862
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9968 8498 9996 8910
rect 10060 8906 10088 9998
rect 10152 9382 10180 10066
rect 10888 9722 10916 11630
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10980 10470 11008 10542
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 10198 11008 10406
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9968 8090 9996 8434
rect 10060 8362 10088 8570
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10060 8022 10088 8298
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 10060 7546 10088 7958
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 6390 9260 6598
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8680 5914 8708 6258
rect 9784 6118 9812 6802
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 9784 5302 9812 6054
rect 10152 5370 10180 9318
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10796 8838 10824 9522
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10520 8566 10548 8774
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 7342 10732 8230
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 7002 10732 7278
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 9772 5296 9824 5302
rect 9770 5264 9772 5273
rect 9824 5264 9826 5273
rect 9770 5199 9826 5208
rect 9784 5173 9812 5199
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 8574 4720 8630 4729
rect 9416 4690 9444 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10796 4758 10824 8774
rect 10888 7546 10916 9386
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 8574 4655 8630 4664
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 6932 4126 7144 4154
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 4894 54 5212 82
rect 6656 82 6684 2246
rect 6932 2009 6960 4126
rect 6918 2000 6974 2009
rect 6918 1935 6974 1944
rect 8312 1193 8340 4422
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 8298 1184 8354 1193
rect 8298 1119 8354 1128
rect 6918 82 6974 480
rect 6656 54 6974 82
rect 938 0 994 54
rect 2870 0 2926 54
rect 4894 0 4950 54
rect 6918 0 6974 54
rect 8850 82 8906 480
rect 9140 82 9168 2450
rect 9416 105 9444 4626
rect 10888 4604 10916 7346
rect 10980 7002 11008 7890
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10796 4576 10916 4604
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3738 10732 4082
rect 10796 4010 10824 4576
rect 11072 4154 11100 13126
rect 11808 12306 11836 13670
rect 11900 12442 11928 14214
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11992 13530 12020 13806
rect 12084 13734 12112 14418
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13530 12112 13670
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12268 13462 12296 13942
rect 12728 13814 12756 14962
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 14482 12848 14826
rect 12912 14618 12940 15914
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15366 13400 15846
rect 13556 15706 13584 15914
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12728 13786 12848 13814
rect 12820 13462 12848 13786
rect 12912 13734 12940 14554
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12808 13456 12860 13462
rect 12808 13398 12860 13404
rect 12636 12442 12664 13398
rect 12820 12918 12848 13398
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11716 11762 11744 12242
rect 11808 11898 11836 12242
rect 12912 11898 12940 13670
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12912 11762 12940 11834
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11348 11286 11376 11630
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11532 11218 11560 11562
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11256 10606 11284 11154
rect 11716 11150 11744 11698
rect 12912 11286 12940 11698
rect 13004 11626 13032 13398
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13188 12986 13216 13330
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13188 12374 13216 12922
rect 13372 12753 13400 15302
rect 13556 14618 13584 15642
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13740 15065 13768 15438
rect 13832 15162 13860 15574
rect 14108 15502 14136 15914
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13726 15056 13782 15065
rect 13726 14991 13782 15000
rect 14108 14890 14136 15438
rect 14292 15434 14320 15846
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 14618 14044 14758
rect 14108 14618 14136 14826
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14016 14074 14044 14554
rect 14292 14521 14320 15370
rect 14278 14512 14334 14521
rect 14278 14447 14334 14456
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13464 12782 13492 13126
rect 13452 12776 13504 12782
rect 13358 12744 13414 12753
rect 13452 12718 13504 12724
rect 13358 12679 13414 12688
rect 13556 12374 13584 13194
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12918 13952 13126
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13176 12368 13228 12374
rect 13176 12310 13228 12316
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13556 12209 13584 12310
rect 13728 12232 13780 12238
rect 13542 12200 13598 12209
rect 13728 12174 13780 12180
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13542 12135 13598 12144
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11520 10532 11572 10538
rect 11520 10474 11572 10480
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 6458 11192 9862
rect 11348 9654 11376 10066
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11532 9178 11560 10474
rect 12268 10266 12296 11154
rect 12360 10810 12388 11222
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 11888 9444 11940 9450
rect 11888 9386 11940 9392
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11336 9104 11388 9110
rect 11336 9046 11388 9052
rect 11348 8294 11376 9046
rect 11900 8974 11928 9386
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11624 8294 11652 8910
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 7993 11652 8230
rect 11610 7984 11666 7993
rect 11610 7919 11666 7928
rect 11900 7886 11928 8910
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12268 7546 12296 7958
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12176 6934 12204 7142
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12268 6866 12296 7482
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12268 6458 12296 6802
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 10888 4126 11100 4154
rect 12360 4146 12388 10202
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12820 9178 12848 10066
rect 12912 9654 12940 11222
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10810 13124 10950
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 13188 10742 13216 11630
rect 13740 11354 13768 12174
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13372 10538 13400 10610
rect 13464 10538 13492 10746
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13280 9722 13308 10066
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12912 9450 12940 9590
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12452 8498 12480 9114
rect 12912 9110 12940 9386
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12912 8634 12940 9046
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12912 8362 12940 8570
rect 12900 8356 12952 8362
rect 12900 8298 12952 8304
rect 13096 8090 13124 8910
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12544 7002 12572 7210
rect 12636 7002 12664 7822
rect 12820 7410 12848 7822
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12544 6322 12572 6938
rect 12820 6866 12848 7346
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 6458 12848 6802
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 13280 5137 13308 6734
rect 13266 5128 13322 5137
rect 13266 5063 13322 5072
rect 12348 4140 12400 4146
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10888 3194 10916 4126
rect 12348 4082 12400 4088
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3670 11468 3878
rect 13372 3670 13400 10474
rect 13740 8498 13768 10950
rect 14016 10606 14044 12174
rect 14108 10810 14136 13874
rect 14384 13814 14412 23462
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 18892 22098 18920 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 17052 21690 17080 22034
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 18616 20369 18644 20742
rect 18602 20360 18658 20369
rect 18602 20295 18658 20304
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 18616 19281 18644 20198
rect 18602 19272 18658 19281
rect 18602 19207 18658 19216
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15488 17814 15516 18090
rect 15672 18086 15700 18770
rect 18326 18728 18382 18737
rect 18248 18698 18326 18714
rect 18236 18692 18326 18698
rect 18288 18686 18326 18692
rect 18326 18663 18382 18672
rect 18236 18634 18288 18640
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15476 17808 15528 17814
rect 15476 17750 15528 17756
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14476 17066 14504 17274
rect 14464 17060 14516 17066
rect 14464 17002 14516 17008
rect 14660 16998 14688 17478
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15488 17338 15516 17750
rect 15672 17678 15700 18022
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 14648 16992 14700 16998
rect 15580 16980 15608 17546
rect 15660 16992 15712 16998
rect 15580 16952 15660 16980
rect 14648 16934 14700 16940
rect 15660 16934 15712 16940
rect 14462 16008 14518 16017
rect 14462 15943 14518 15952
rect 14292 13786 14412 13814
rect 14292 13394 14320 13786
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14384 13326 14412 13670
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12986 14228 13194
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14292 12170 14320 12854
rect 14384 12850 14412 13262
rect 14476 12986 14504 15943
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14384 11558 14412 12310
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14200 11354 14228 11494
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14384 11286 14412 11494
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14476 10198 14504 12786
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 14292 8362 14320 8774
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 6798 13768 7822
rect 13832 7410 13860 7958
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 14108 7342 14136 8230
rect 14292 7857 14320 8298
rect 14384 8022 14412 8434
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14278 7848 14334 7857
rect 14278 7783 14334 7792
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14108 7002 14136 7278
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 5137 13492 6598
rect 13450 5128 13506 5137
rect 13450 5063 13506 5072
rect 14568 4154 14596 14010
rect 14660 13841 14688 16934
rect 15672 16726 15700 16934
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16046 15332 16526
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15304 15434 15332 15982
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15396 15162 15424 15506
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14752 13938 14780 14350
rect 14844 14074 14872 14826
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14844 13938 14872 14010
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14832 13932 14884 13938
rect 15304 13920 15332 14894
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 14346 15424 14418
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15396 14074 15424 14282
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 14832 13874 14884 13880
rect 15120 13892 15332 13920
rect 14646 13832 14702 13841
rect 15120 13814 15148 13892
rect 14844 13802 15148 13814
rect 14646 13767 14702 13776
rect 14832 13796 15148 13802
rect 14884 13786 15148 13796
rect 15290 13832 15346 13841
rect 15290 13767 15346 13776
rect 14832 13738 14884 13744
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14660 9586 14688 13330
rect 14844 12918 14872 13330
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11898 14780 12174
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11830 14872 12854
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11898 15332 13767
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 12782 15424 13126
rect 15488 12782 15516 15914
rect 15580 15910 15608 16594
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 13394 15608 15846
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16040 12782 16068 13330
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15396 12374 15424 12718
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12442 15700 12582
rect 16040 12442 16068 12718
rect 16224 12714 16252 13738
rect 18248 13530 18276 13806
rect 18432 13734 18460 15914
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15065 18644 15846
rect 18602 15056 18658 15065
rect 18602 14991 18658 15000
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 16212 12708 16264 12714
rect 16212 12650 16264 12656
rect 17328 12646 17356 13330
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15488 11830 15516 12106
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15580 11762 15608 12310
rect 17328 12170 17356 12582
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 14752 11014 14780 11698
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15212 11354 15240 11562
rect 18248 11558 18276 12242
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14752 8974 14780 10406
rect 15304 9926 15332 10542
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15396 9722 15424 11290
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 15764 10606 15792 11154
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10810 15884 11086
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16960 10742 16988 11154
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8090 15332 9114
rect 15580 8634 15608 9862
rect 15948 9722 15976 10066
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 8974 15700 9522
rect 15948 9178 15976 9658
rect 18156 9625 18184 10406
rect 18248 10062 18276 11494
rect 19352 10810 19380 23598
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20732 15978 20760 27526
rect 20902 27520 20958 27526
rect 22834 27520 22890 28000
rect 24858 27520 24914 28000
rect 26882 27520 26938 28000
rect 22848 23866 22876 27520
rect 24674 26344 24730 26353
rect 24674 26279 24730 26288
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 21192 22545 21220 23530
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 21178 22536 21234 22545
rect 21178 22471 21234 22480
rect 22848 22438 22876 23122
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22848 22001 22876 22374
rect 22834 21992 22890 22001
rect 22834 21927 22890 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 24596 18737 24624 18770
rect 24582 18728 24638 18737
rect 24582 18663 24638 18672
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24584 18352 24636 18358
rect 24490 18320 24546 18329
rect 24546 18300 24584 18306
rect 24546 18294 24636 18300
rect 24546 18278 24624 18294
rect 24490 18255 24546 18264
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16046 24716 26279
rect 24872 23322 24900 27520
rect 25134 24168 25190 24177
rect 25134 24103 25190 24112
rect 25148 23866 25176 24103
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25148 23662 25176 23802
rect 25136 23656 25188 23662
rect 25136 23598 25188 23604
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24766 21992 24822 22001
rect 24766 21927 24822 21936
rect 24780 20602 24808 21927
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25240 20602 25268 20946
rect 26896 20602 26924 27520
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 26884 20596 26936 20602
rect 26884 20538 26936 20544
rect 24766 19816 24822 19825
rect 24766 19751 24822 19760
rect 24780 18970 24808 19751
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 25412 18828 25464 18834
rect 25412 18770 25464 18776
rect 25424 18426 25452 18770
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27632 18193 27660 18226
rect 27618 18184 27674 18193
rect 27618 18119 27674 18128
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 24766 15600 24822 15609
rect 24676 15564 24728 15570
rect 24766 15535 24822 15544
rect 24676 15506 24728 15512
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15506
rect 24780 15434 24808 15535
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24124 14952 24176 14958
rect 24124 14894 24176 14900
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 24136 14385 24164 14894
rect 24122 14376 24178 14385
rect 24122 14311 24178 14320
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24674 13696 24730 13705
rect 19622 13628 19918 13648
rect 24674 13631 24730 13640
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 24688 13394 24716 13631
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12986 24716 13330
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 27618 11792 27674 11801
rect 27618 11727 27674 11736
rect 27632 11694 27660 11727
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 23756 10600 23808 10606
rect 23756 10542 23808 10548
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18142 9616 18198 9625
rect 18142 9551 18198 9560
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16960 9042 16988 9386
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15580 8294 15608 8570
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15396 7546 15424 7958
rect 15672 7886 15700 8910
rect 16132 8498 16160 8910
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15856 8090 15884 8298
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 16132 7342 16160 8434
rect 16224 8022 16252 8910
rect 16960 8634 16988 8978
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 16212 8016 16264 8022
rect 18616 7993 18644 8230
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 16212 7958 16264 7964
rect 18602 7984 18658 7993
rect 18602 7919 18658 7928
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7546 16252 7686
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 6866 15884 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15856 6458 15884 6802
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14476 4126 14596 4154
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 11440 3194 11468 3606
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11532 2854 11560 3470
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12544 3058 12572 3334
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 8850 54 9168 82
rect 9402 96 9458 105
rect 8850 0 8906 54
rect 10796 82 10824 2790
rect 11532 2650 11560 2790
rect 12544 2650 12572 2994
rect 12912 2922 12940 3470
rect 13372 3058 13400 3606
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13464 3194 13492 3538
rect 14476 3194 14504 4126
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 14476 2990 14504 3130
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 14004 2848 14056 2854
rect 14004 2790 14056 2796
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 14016 2514 14044 2790
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 10874 82 10930 480
rect 10796 54 10930 82
rect 12544 82 12572 2246
rect 12898 82 12954 480
rect 12544 54 12954 82
rect 14568 82 14596 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 16040 2009 16068 2246
rect 16026 2000 16082 2009
rect 16026 1935 16082 1944
rect 14922 82 14978 480
rect 14568 54 14978 82
rect 16684 82 16712 6598
rect 17052 6118 17080 6802
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 16854 82 16910 480
rect 16684 54 16910 82
rect 18616 82 18644 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20824 5137 20852 6190
rect 20810 5128 20866 5137
rect 20810 5063 20866 5072
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 18878 82 18934 480
rect 18616 54 18934 82
rect 20640 82 20668 2246
rect 20902 82 20958 480
rect 20640 54 20958 82
rect 9402 31 9458 40
rect 10874 0 10930 54
rect 12898 0 12954 54
rect 14922 0 14978 54
rect 16854 0 16910 54
rect 18878 0 18934 54
rect 20902 0 20958 54
rect 22834 82 22890 480
rect 22940 82 22968 6326
rect 23768 134 23796 10542
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 25134 9072 25190 9081
rect 25134 9007 25190 9016
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 25148 8634 25176 9007
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25148 8430 25176 8570
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 24122 7848 24178 7857
rect 24122 7783 24178 7792
rect 24136 7410 24164 7783
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 25516 7206 25544 7890
rect 27618 7440 27674 7449
rect 27618 7375 27674 7384
rect 27632 7342 27660 7375
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 22834 54 22968 82
rect 23756 128 23808 134
rect 23756 70 23808 76
rect 24858 128 24914 480
rect 24858 76 24860 128
rect 24912 76 24914 128
rect 22834 0 22890 54
rect 24858 0 24914 76
rect 26528 82 26556 7142
rect 26606 5264 26662 5273
rect 26606 5199 26662 5208
rect 26620 3641 26648 5199
rect 26606 3632 26662 3641
rect 26606 3567 26662 3576
rect 27618 1048 27674 1057
rect 27618 983 27674 992
rect 26882 82 26938 480
rect 27632 105 27660 983
rect 26528 54 26938 82
rect 26882 0 26938 54
rect 27618 96 27674 105
rect 27618 31 27674 40
<< via2 >>
rect 110 24520 166 24576
rect 2502 26696 2558 26752
rect 1306 25336 1362 25392
rect 1214 22616 1270 22672
rect 1582 21256 1638 21312
rect 1582 20032 1638 20088
rect 1582 18672 1638 18728
rect 1582 15680 1638 15736
rect 1766 15952 1822 16008
rect 1950 16496 2006 16552
rect 1490 9288 1546 9344
rect 1306 7928 1362 7984
rect 110 4528 166 4584
rect 110 3168 166 3224
rect 754 2216 810 2272
rect 1674 6704 1730 6760
rect 2962 18672 3018 18728
rect 2870 12688 2926 12744
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 3606 17312 3662 17368
rect 3422 9560 3478 9616
rect 3054 5072 3110 5128
rect 3790 13640 3846 13696
rect 3698 12824 3754 12880
rect 4066 5344 4122 5400
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9218 21936 9274 21992
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 6090 15952 6146 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5170 14320 5226 14376
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6550 12164 6606 12200
rect 6550 12144 6552 12164
rect 6552 12144 6604 12164
rect 6604 12144 6606 12164
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6366 10648 6422 10704
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9402 19216 9458 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 13450 22480 13506 22536
rect 12898 20304 12954 20360
rect 12990 18672 13046 18728
rect 12806 18264 12862 18320
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 11518 16496 11574 16552
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9218 14456 9274 14512
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9126 12144 9182 12200
rect 9678 12144 9734 12200
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 9770 5244 9772 5264
rect 9772 5244 9824 5264
rect 9824 5244 9826 5264
rect 9770 5208 9826 5244
rect 8574 4664 8630 4720
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6918 1944 6974 2000
rect 8298 1128 8354 1184
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 13726 15000 13782 15056
rect 14278 14456 14334 14512
rect 13358 12688 13414 12744
rect 13542 12144 13598 12200
rect 11610 7928 11666 7984
rect 13266 5072 13322 5128
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 18602 20304 18658 20360
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 18602 19216 18658 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 18326 18672 18382 18728
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14462 15952 14518 16008
rect 14278 7792 14334 7848
rect 13450 5072 13506 5128
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14646 13776 14702 13832
rect 15290 13776 15346 13832
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 18602 15000 18658 15056
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 24674 26288 24730 26344
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 21178 22480 21234 22536
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 22834 21936 22890 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24582 18672 24638 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24490 18264 24546 18320
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25134 24112 25190 24168
rect 24766 21936 24822 21992
rect 24766 19760 24822 19816
rect 27618 18128 27674 18184
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 24766 15544 24822 15600
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 24122 14320 24178 14376
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24674 13640 24730 13696
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 27618 11736 27674 11792
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18142 9560 18198 9616
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 18602 7928 18658 7984
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 9402 40 9458 96
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 16026 1944 16082 2000
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20810 5072 20866 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 25134 9016 25190 9072
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24122 7792 24178 7848
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 27618 7384 27674 7440
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 26606 5208 26662 5264
rect 26606 3576 26662 3632
rect 27618 992 27674 1048
rect 27618 40 27674 96
<< metal3 >>
rect 0 27208 480 27328
rect 62 26754 122 27208
rect 27520 26800 28000 26920
rect 2497 26754 2563 26757
rect 62 26752 2563 26754
rect 62 26696 2502 26752
rect 2558 26696 2563 26752
rect 62 26694 2563 26696
rect 2497 26691 2563 26694
rect 24669 26346 24735 26349
rect 27662 26346 27722 26800
rect 24669 26344 27722 26346
rect 24669 26288 24674 26344
rect 24730 26288 27722 26344
rect 24669 26286 27722 26288
rect 24669 26283 24735 26286
rect 0 25848 480 25968
rect 62 25394 122 25848
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1301 25394 1367 25397
rect 62 25392 1367 25394
rect 62 25336 1306 25392
rect 1362 25336 1367 25392
rect 62 25334 1367 25336
rect 1301 25331 1367 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 27520 24624 28000 24744
rect 0 24576 480 24608
rect 0 24520 110 24576
rect 166 24520 480 24576
rect 0 24488 480 24520
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 25129 24170 25195 24173
rect 27662 24170 27722 24624
rect 25129 24168 27722 24170
rect 25129 24112 25134 24168
rect 25190 24112 27722 24168
rect 25129 24110 27722 24112
rect 25129 24107 25195 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 62 22674 122 23128
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1209 22674 1275 22677
rect 62 22672 1275 22674
rect 62 22616 1214 22672
rect 1270 22616 1275 22672
rect 62 22614 1275 22616
rect 1209 22611 1275 22614
rect 13445 22538 13511 22541
rect 21173 22538 21239 22541
rect 13445 22536 21239 22538
rect 13445 22480 13450 22536
rect 13506 22480 21178 22536
rect 21234 22480 21239 22536
rect 13445 22478 21239 22480
rect 13445 22475 13511 22478
rect 21173 22475 21239 22478
rect 27520 22448 28000 22568
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 9213 21994 9279 21997
rect 22829 21994 22895 21997
rect 9213 21992 22895 21994
rect 9213 21936 9218 21992
rect 9274 21936 22834 21992
rect 22890 21936 22895 21992
rect 9213 21934 22895 21936
rect 9213 21931 9279 21934
rect 22829 21931 22895 21934
rect 24761 21994 24827 21997
rect 27662 21994 27722 22448
rect 24761 21992 27722 21994
rect 24761 21936 24766 21992
rect 24822 21936 27722 21992
rect 24761 21934 27722 21936
rect 24761 21931 24827 21934
rect 0 21768 480 21888
rect 5610 21792 5930 21793
rect 62 21314 122 21768
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1577 21314 1643 21317
rect 62 21312 1643 21314
rect 62 21256 1582 21312
rect 1638 21256 1643 21312
rect 62 21254 1643 21256
rect 1577 21251 1643 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 5610 20704 5930 20705
rect 0 20544 480 20664
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 62 20090 122 20544
rect 12893 20362 12959 20365
rect 18597 20362 18663 20365
rect 12893 20360 18663 20362
rect 12893 20304 12898 20360
rect 12954 20304 18602 20360
rect 18658 20304 18663 20360
rect 12893 20302 18663 20304
rect 12893 20299 12959 20302
rect 18597 20299 18663 20302
rect 27520 20272 28000 20392
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1577 20090 1643 20093
rect 62 20088 1643 20090
rect 62 20032 1582 20088
rect 1638 20032 1643 20088
rect 62 20030 1643 20032
rect 1577 20027 1643 20030
rect 24761 19818 24827 19821
rect 27662 19818 27722 20272
rect 24761 19816 27722 19818
rect 24761 19760 24766 19816
rect 24822 19760 27722 19816
rect 24761 19758 27722 19760
rect 24761 19755 24827 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19184 480 19304
rect 9397 19274 9463 19277
rect 18597 19274 18663 19277
rect 9397 19272 18663 19274
rect 9397 19216 9402 19272
rect 9458 19216 18602 19272
rect 18658 19216 18663 19272
rect 9397 19214 18663 19216
rect 9397 19211 9463 19214
rect 18597 19211 18663 19214
rect 62 18730 122 19184
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 1577 18730 1643 18733
rect 62 18728 1643 18730
rect 62 18672 1582 18728
rect 1638 18672 1643 18728
rect 62 18670 1643 18672
rect 1577 18667 1643 18670
rect 2957 18730 3023 18733
rect 12985 18730 13051 18733
rect 2957 18728 13051 18730
rect 2957 18672 2962 18728
rect 3018 18672 12990 18728
rect 13046 18672 13051 18728
rect 2957 18670 13051 18672
rect 2957 18667 3023 18670
rect 12985 18667 13051 18670
rect 18321 18730 18387 18733
rect 24577 18730 24643 18733
rect 18321 18728 24643 18730
rect 18321 18672 18326 18728
rect 18382 18672 24582 18728
rect 24638 18672 24643 18728
rect 18321 18670 24643 18672
rect 18321 18667 18387 18670
rect 24577 18667 24643 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 12801 18322 12867 18325
rect 24485 18322 24551 18325
rect 12801 18320 24551 18322
rect 12801 18264 12806 18320
rect 12862 18264 24490 18320
rect 24546 18264 24551 18320
rect 12801 18262 24551 18264
rect 12801 18259 12867 18262
rect 24485 18259 24551 18262
rect 27520 18184 28000 18216
rect 27520 18128 27618 18184
rect 27674 18128 28000 18184
rect 27520 18096 28000 18128
rect 10277 17984 10597 17985
rect 0 17824 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 62 17370 122 17824
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 3601 17370 3667 17373
rect 62 17368 3667 17370
rect 62 17312 3606 17368
rect 3662 17312 3667 17368
rect 62 17310 3667 17312
rect 3601 17307 3667 17310
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16464 480 16584
rect 1945 16554 2011 16557
rect 11513 16554 11579 16557
rect 1945 16552 11579 16554
rect 1945 16496 1950 16552
rect 2006 16496 11518 16552
rect 11574 16496 11579 16552
rect 1945 16494 11579 16496
rect 1945 16491 2011 16494
rect 11513 16491 11579 16494
rect 62 16010 122 16464
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 1761 16010 1827 16013
rect 62 16008 1827 16010
rect 62 15952 1766 16008
rect 1822 15952 1827 16008
rect 62 15950 1827 15952
rect 1761 15947 1827 15950
rect 6085 16010 6151 16013
rect 14457 16010 14523 16013
rect 6085 16008 14523 16010
rect 6085 15952 6090 16008
rect 6146 15952 14462 16008
rect 14518 15952 14523 16008
rect 6085 15950 14523 15952
rect 6085 15947 6151 15950
rect 14457 15947 14523 15950
rect 27520 15920 28000 16040
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1577 15738 1643 15741
rect 62 15736 1643 15738
rect 62 15680 1582 15736
rect 1638 15680 1643 15736
rect 62 15678 1643 15680
rect 62 15224 122 15678
rect 1577 15675 1643 15678
rect 24761 15602 24827 15605
rect 27662 15602 27722 15920
rect 24761 15600 27722 15602
rect 24761 15544 24766 15600
rect 24822 15544 27722 15600
rect 24761 15542 27722 15544
rect 24761 15539 24827 15542
rect 5610 15264 5930 15265
rect 0 15104 480 15224
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 13721 15058 13787 15061
rect 18597 15058 18663 15061
rect 13721 15056 18663 15058
rect 13721 15000 13726 15056
rect 13782 15000 18602 15056
rect 18658 15000 18663 15056
rect 13721 14998 18663 15000
rect 13721 14995 13787 14998
rect 18597 14995 18663 14998
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 9213 14514 9279 14517
rect 14273 14514 14339 14517
rect 9213 14512 14339 14514
rect 9213 14456 9218 14512
rect 9274 14456 14278 14512
rect 14334 14456 14339 14512
rect 9213 14454 14339 14456
rect 9213 14451 9279 14454
rect 14273 14451 14339 14454
rect 5165 14378 5231 14381
rect 24117 14378 24183 14381
rect 5165 14376 24183 14378
rect 5165 14320 5170 14376
rect 5226 14320 24122 14376
rect 24178 14320 24183 14376
rect 5165 14318 24183 14320
rect 5165 14315 5231 14318
rect 24117 14315 24183 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13972 480 14000
rect 0 13908 60 13972
rect 124 13908 480 13972
rect 0 13880 480 13908
rect 27520 13880 28000 14000
rect 14641 13834 14707 13837
rect 15285 13834 15351 13837
rect 14641 13832 15351 13834
rect 14641 13776 14646 13832
rect 14702 13776 15290 13832
rect 15346 13776 15351 13832
rect 14641 13774 15351 13776
rect 14641 13771 14707 13774
rect 15285 13771 15351 13774
rect 54 13636 60 13700
rect 124 13698 130 13700
rect 3785 13698 3851 13701
rect 124 13696 3851 13698
rect 124 13640 3790 13696
rect 3846 13640 3851 13696
rect 124 13638 3851 13640
rect 124 13636 130 13638
rect 3785 13635 3851 13638
rect 24669 13698 24735 13701
rect 27662 13698 27722 13880
rect 24669 13696 27722 13698
rect 24669 13640 24674 13696
rect 24730 13640 27722 13696
rect 24669 13638 27722 13640
rect 24669 13635 24735 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 3693 12882 3759 12885
rect 62 12880 3759 12882
rect 62 12824 3698 12880
rect 3754 12824 3759 12880
rect 62 12822 3759 12824
rect 62 12640 122 12822
rect 3693 12819 3759 12822
rect 2865 12746 2931 12749
rect 13353 12746 13419 12749
rect 2865 12744 13419 12746
rect 2865 12688 2870 12744
rect 2926 12688 13358 12744
rect 13414 12688 13419 12744
rect 2865 12686 13419 12688
rect 2865 12683 2931 12686
rect 13353 12683 13419 12686
rect 0 12520 480 12640
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 6545 12202 6611 12205
rect 9121 12202 9187 12205
rect 9673 12202 9739 12205
rect 13537 12202 13603 12205
rect 6545 12200 13603 12202
rect 6545 12144 6550 12200
rect 6606 12144 9126 12200
rect 9182 12144 9678 12200
rect 9734 12144 13542 12200
rect 13598 12144 13603 12200
rect 6545 12142 13603 12144
rect 6545 12139 6611 12142
rect 9121 12139 9187 12142
rect 9673 12139 9739 12142
rect 13537 12139 13603 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27520 11792 28000 11824
rect 27520 11736 27618 11792
rect 27674 11736 28000 11792
rect 27520 11704 28000 11736
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 0 11160 480 11280
rect 62 10706 122 11160
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 6361 10706 6427 10709
rect 62 10704 6427 10706
rect 62 10648 6366 10704
rect 6422 10648 6427 10704
rect 62 10646 6427 10648
rect 6361 10643 6427 10646
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 0 9800 480 9920
rect 5610 9824 5930 9825
rect 62 9346 122 9800
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 3417 9618 3483 9621
rect 18137 9618 18203 9621
rect 3417 9616 18203 9618
rect 3417 9560 3422 9616
rect 3478 9560 18142 9616
rect 18198 9560 18203 9616
rect 3417 9558 18203 9560
rect 3417 9555 3483 9558
rect 18137 9555 18203 9558
rect 27520 9528 28000 9648
rect 1485 9346 1551 9349
rect 62 9344 1551 9346
rect 62 9288 1490 9344
rect 1546 9288 1551 9344
rect 62 9286 1551 9288
rect 1485 9283 1551 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 25129 9074 25195 9077
rect 27662 9074 27722 9528
rect 25129 9072 27722 9074
rect 25129 9016 25134 9072
rect 25190 9016 27722 9072
rect 25129 9014 27722 9016
rect 25129 9011 25195 9014
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 0 8440 480 8560
rect 62 7986 122 8440
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 1301 7986 1367 7989
rect 62 7984 1367 7986
rect 62 7928 1306 7984
rect 1362 7928 1367 7984
rect 62 7926 1367 7928
rect 1301 7923 1367 7926
rect 11605 7986 11671 7989
rect 18597 7986 18663 7989
rect 11605 7984 18663 7986
rect 11605 7928 11610 7984
rect 11666 7928 18602 7984
rect 18658 7928 18663 7984
rect 11605 7926 18663 7928
rect 11605 7923 11671 7926
rect 18597 7923 18663 7926
rect 14273 7850 14339 7853
rect 24117 7850 24183 7853
rect 14273 7848 24183 7850
rect 14273 7792 14278 7848
rect 14334 7792 24122 7848
rect 24178 7792 24183 7848
rect 14273 7790 24183 7792
rect 14273 7787 14339 7790
rect 24117 7787 24183 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7440 28000 7472
rect 27520 7384 27618 7440
rect 27674 7384 28000 7440
rect 27520 7352 28000 7384
rect 0 7216 480 7336
rect 62 6762 122 7216
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 1669 6762 1735 6765
rect 62 6760 1735 6762
rect 62 6704 1674 6760
rect 1730 6704 1735 6760
rect 62 6702 1735 6704
rect 1669 6699 1735 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 10277 6016 10597 6017
rect 0 5856 480 5976
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 62 5402 122 5856
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 4061 5402 4127 5405
rect 62 5400 4127 5402
rect 62 5344 4066 5400
rect 4122 5344 4127 5400
rect 62 5342 4127 5344
rect 4061 5339 4127 5342
rect 9765 5266 9831 5269
rect 26601 5266 26667 5269
rect 9765 5264 26667 5266
rect 9765 5208 9770 5264
rect 9826 5208 26606 5264
rect 26662 5208 26667 5264
rect 9765 5206 26667 5208
rect 9765 5203 9831 5206
rect 26601 5203 26667 5206
rect 27520 5176 28000 5296
rect 3049 5130 3115 5133
rect 13261 5130 13327 5133
rect 3049 5128 13327 5130
rect 3049 5072 3054 5128
rect 3110 5072 13266 5128
rect 13322 5072 13327 5128
rect 3049 5070 13327 5072
rect 3049 5067 3115 5070
rect 13261 5067 13327 5070
rect 13445 5130 13511 5133
rect 20805 5130 20871 5133
rect 13445 5128 20871 5130
rect 13445 5072 13450 5128
rect 13506 5072 20810 5128
rect 20866 5072 20871 5128
rect 13445 5070 20871 5072
rect 13445 5067 13511 5070
rect 20805 5067 20871 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 8569 4722 8635 4725
rect 27662 4722 27722 5176
rect 8569 4720 27722 4722
rect 8569 4664 8574 4720
rect 8630 4664 27722 4720
rect 8569 4662 27722 4664
rect 8569 4659 8635 4662
rect 0 4584 480 4616
rect 0 4528 110 4584
rect 166 4528 480 4584
rect 0 4496 480 4528
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 26601 3634 26667 3637
rect 26601 3632 27722 3634
rect 26601 3576 26606 3632
rect 26662 3576 27722 3632
rect 26601 3574 27722 3576
rect 26601 3571 26667 3574
rect 5610 3296 5930 3297
rect 0 3224 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 0 3168 110 3224
rect 166 3168 480 3224
rect 0 3136 480 3168
rect 27662 3120 27722 3574
rect 27520 3000 28000 3120
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 749 2274 815 2277
rect 62 2272 815 2274
rect 62 2216 754 2272
rect 810 2216 815 2272
rect 62 2214 815 2216
rect 62 1896 122 2214
rect 749 2211 815 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6913 2002 6979 2005
rect 16021 2002 16087 2005
rect 6913 2000 16087 2002
rect 6913 1944 6918 2000
rect 6974 1944 16026 2000
rect 16082 1944 16087 2000
rect 6913 1942 16087 1944
rect 6913 1939 6979 1942
rect 16021 1939 16087 1942
rect 0 1776 480 1896
rect 8293 1186 8359 1189
rect 62 1184 8359 1186
rect 62 1128 8298 1184
rect 8354 1128 8359 1184
rect 62 1126 8359 1128
rect 62 672 122 1126
rect 8293 1123 8359 1126
rect 27520 1048 28000 1080
rect 27520 992 27618 1048
rect 27674 992 28000 1048
rect 27520 960 28000 992
rect 0 552 480 672
rect 9397 98 9463 101
rect 27613 98 27679 101
rect 9397 96 27679 98
rect 9397 40 9402 96
rect 9458 40 27618 96
rect 27674 40 27679 96
rect 9397 38 27679 40
rect 9397 35 9463 38
rect 27613 35 27679 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 60 13908 124 13972
rect 60 13636 124 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 59 13972 125 13973
rect 59 13908 60 13972
rect 124 13908 125 13972
rect 59 13907 125 13908
rect 62 13701 122 13907
rect 59 13700 125 13701
rect 59 13636 60 13700
rect 124 13636 125 13700
rect 59 13635 125 13636
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_fill_2  FILLER_1_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_22 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_44 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_53
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_46
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_57 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_61
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_97
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_101
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _230_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_193
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_197
timestamp 1586364061
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_201
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_8  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_28
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_60
timestamp 1586364061
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_69
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_17
timestamp 1586364061
transform 1 0 2668 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_64
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_58
timestamp 1586364061
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_76
timestamp 1586364061
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_87
timestamp 1586364061
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_91
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_103
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_35
timestamp 1586364061
transform 1 0 4324 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_49
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_59
timestamp 1586364061
transform 1 0 6532 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_67
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_68
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 866 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 8648 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_72
timestamp 1586364061
transform 1 0 7728 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 406 592
use scs8hd_conb_1  _211_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_126
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_131
timestamp 1586364061
transform 1 0 13156 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_159
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_162
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_182
timestamp 1586364061
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_218
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_242
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_8
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_38
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_51
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_55
timestamp 1586364061
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _103_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 590 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_96
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_150
timestamp 1586364061
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_175
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_199
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_32
timestamp 1586364061
transform 1 0 4048 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _151_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_55
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_82
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 774 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_93
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_97
timestamp 1586364061
transform 1 0 10028 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_102
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_164
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_168
timestamp 1586364061
transform 1 0 16560 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_9_274
timestamp 1586364061
transform 1 0 26312 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_14
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_26
timestamp 1586364061
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_48
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_69
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_82
timestamp 1586364061
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_90
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_198
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_8
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_23
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 406 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_34
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_181
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_258
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_262
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_17
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_40
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 774 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 682 592
use scs8hd_decap_3  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_72
timestamp 1586364061
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_118
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_122
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_192
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_14
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_35
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_59
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_83
timestamp 1586364061
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 9292 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_87
timestamp 1586364061
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_91
timestamp 1586364061
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_123
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_151
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_161
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_165
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_181
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_199
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_211
timestamp 1586364061
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_47
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 406 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_128
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_141
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_145
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_173
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_177
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_252
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_264
timestamp 1586364061
transform 1 0 25392 0 1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_60
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 10580 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_101
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12144 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_112
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_131
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 130 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_142
timestamp 1586364061
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_192
timestamp 1586364061
transform 1 0 18768 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_31
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_35
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_48
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_52
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_56
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_65
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 406 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 130 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_85
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_127
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_188
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_200
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_212
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_258
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_262
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_41
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_45
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_58
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_87
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_91
timestamp 1586364061
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_107
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_111
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_4  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_18_174
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 774 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_185
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_6
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_10
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_25
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_17
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_29
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_33
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_37
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_54
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_57
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_67
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 314 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 866 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_78
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_84
timestamp 1586364061
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 866 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_115
timestamp 1586364061
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_166
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_170
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_174
timestamp 1586364061
transform 1 0 17112 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_178
timestamp 1586364061
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_182
timestamp 1586364061
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_198
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_210
timestamp 1586364061
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_40
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_44
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_52
timestamp 1586364061
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_73
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_139
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_143
timestamp 1586364061
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_181
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_190
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_194
timestamp 1586364061
transform 1 0 18952 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_206
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_242
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_29
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_43
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_47
timestamp 1586364061
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use scs8hd_nor3_4  _170_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_58
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_62
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_79
timestamp 1586364061
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_110
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_118
timestamp 1586364061
transform 1 0 11960 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_198
timestamp 1586364061
transform 1 0 19320 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_210
timestamp 1586364061
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_19
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_23
timestamp 1586364061
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 7360 0 1 14688
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_81
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_85
timestamp 1586364061
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_102
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 406 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_23_182
timestamp 1586364061
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_248
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_252
timestamp 1586364061
transform 1 0 24288 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_18
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_30
timestamp 1586364061
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_53
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_63
timestamp 1586364061
transform 1 0 6900 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 130 592
use scs8hd_nor3_4  _169_
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 1234 592
use scs8hd_fill_1  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_96
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_100
timestamp 1586364061
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_118
timestamp 1586364061
transform 1 0 11960 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_199
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_211
timestamp 1586364061
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_17
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_21
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 590 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5244 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_42
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_65
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_69
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_73
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_95
timestamp 1586364061
transform 1 0 9844 0 1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_262
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_25_274
timestamp 1586364061
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_14
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_18
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_29
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_67
timestamp 1586364061
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_71
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_85
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12512 0 1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_116
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_139
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_160
timestamp 1586364061
transform 1 0 15824 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_172
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_199
timestamp 1586364061
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_39
timestamp 1586364061
transform 1 0 4692 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_42
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_60
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_67
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_4  FILLER_28_71
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_97
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 774 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_120
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_137
timestamp 1586364061
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_175
timestamp 1586364061
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_187
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_199
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_211
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_18
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_26
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 590 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_72
timestamp 1586364061
transform 1 0 7728 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_165
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_177
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_262
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 4232 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_43
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_47
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_83
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_86
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_139
timestamp 1586364061
transform 1 0 13892 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_151
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_169
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_181
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_205
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_14
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_19
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 590 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_36
timestamp 1586364061
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_40
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_79
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_139
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_151
timestamp 1586364061
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_9
timestamp 1586364061
transform 1 0 1932 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_20
timestamp 1586364061
transform 1 0 2944 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_28
timestamp 1586364061
transform 1 0 3680 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_39
timestamp 1586364061
transform 1 0 4692 0 -1 20128
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_43
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_58
timestamp 1586364061
transform 1 0 6440 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_79
timestamp 1586364061
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_91
timestamp 1586364061
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_32_123
timestamp 1586364061
transform 1 0 12420 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_140
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_36
timestamp 1586364061
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_40
timestamp 1586364061
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_35
timestamp 1586364061
transform 1 0 4324 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_43
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_46
timestamp 1586364061
transform 1 0 5336 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 590 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_73
timestamp 1586364061
transform 1 0 7820 0 1 20128
box -38 -48 590 592
use scs8hd_decap_6  FILLER_34_73
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_84
timestamp 1586364061
transform 1 0 8832 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_6  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_99
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_34_109
timestamp 1586364061
transform 1 0 11132 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_116
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_130
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_148
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_142
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_150
timestamp 1586364061
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_172
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_180
timestamp 1586364061
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_259
timestamp 1586364061
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_258
timestamp 1586364061
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_263
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_275
timestamp 1586364061
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_270
timestamp 1586364061
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_274
timestamp 1586364061
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_38
timestamp 1586364061
transform 1 0 4600 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_99
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_112
timestamp 1586364061
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use scs8hd_decap_4  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_35_174
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_182
timestamp 1586364061
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_18
timestamp 1586364061
transform 1 0 2760 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_30
timestamp 1586364061
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_36_39
timestamp 1586364061
transform 1 0 4692 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_43
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_46
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_54
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 314 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 6348 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_60
timestamp 1586364061
transform 1 0 6624 0 -1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_77
timestamp 1586364061
transform 1 0 8188 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_81
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_89
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_112
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_175
timestamp 1586364061
transform 1 0 17204 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_187
timestamp 1586364061
transform 1 0 18308 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_34
timestamp 1586364061
transform 1 0 4232 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_46
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 6992 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_58
timestamp 1586364061
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_73
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_77
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_80
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_90
timestamp 1586364061
transform 1 0 9384 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_113
timestamp 1586364061
transform 1 0 11500 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_136
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_238
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_35
timestamp 1586364061
transform 1 0 4324 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_47
timestamp 1586364061
transform 1 0 5428 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_59
timestamp 1586364061
transform 1 0 6532 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8280 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_77
timestamp 1586364061
transform 1 0 8188 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_81
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_38_89
timestamp 1586364061
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_4  FILLER_38_96
timestamp 1586364061
transform 1 0 9936 0 -1 23392
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10304 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12236 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_113
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_38_130
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_142
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_150
timestamp 1586364061
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_235
timestamp 1586364061
transform 1 0 22724 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 22816 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_240
timestamp 1586364061
transform 1 0 23184 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_252
timestamp 1586364061
transform 1 0 24288 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_264
timestamp 1586364061
transform 1 0 25392 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_272
timestamp 1586364061
transform 1 0 26128 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_52
timestamp 1586364061
transform 1 0 5888 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_56
timestamp 1586364061
transform 1 0 6256 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_60
timestamp 1586364061
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_94
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 314 592
use scs8hd_decap_6  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 590 592
use scs8hd_conb_1  _222_
timestamp 1586364061
transform 1 0 10212 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_105
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_112
timestamp 1586364061
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_116
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 590 592
use scs8hd_decap_4  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_114
timestamp 1586364061
transform 1 0 11592 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_134
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_126
timestamp 1586364061
transform 1 0 12696 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_138
timestamp 1586364061
transform 1 0 13800 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_146
timestamp 1586364061
transform 1 0 14536 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_150
timestamp 1586364061
transform 1 0 14904 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_157
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_161
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_173
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_181
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_234
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_242
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_262
timestamp 1586364061
transform 1 0 25208 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 938 27520 994 28000 6 address[0]
port 0 nsew default input
rlabel metal3 s 27520 960 28000 1080 6 address[1]
port 1 nsew default input
rlabel metal2 s 4894 0 4950 480 6 address[2]
port 2 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 552 480 672 6 address[4]
port 4 nsew default input
rlabel metal3 s 27520 5176 28000 5296 6 address[5]
port 5 nsew default input
rlabel metal2 s 6918 0 6974 480 6 bottom_left_grid_pin_13_
port 6 nsew default input
rlabel metal2 s 10874 0 10930 480 6 bottom_right_grid_pin_11_
port 7 nsew default input
rlabel metal3 s 0 4496 480 4616 6 bottom_right_grid_pin_13_
port 8 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 bottom_right_grid_pin_15_
port 9 nsew default input
rlabel metal3 s 0 1776 480 1896 6 bottom_right_grid_pin_1_
port 10 nsew default input
rlabel metal3 s 27520 7352 28000 7472 6 bottom_right_grid_pin_3_
port 11 nsew default input
rlabel metal2 s 8850 0 8906 480 6 bottom_right_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 2870 27520 2926 28000 6 bottom_right_grid_pin_7_
port 13 nsew default input
rlabel metal3 s 0 3136 480 3256 6 bottom_right_grid_pin_9_
port 14 nsew default input
rlabel metal2 s 4894 27520 4950 28000 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal2 s 12898 0 12954 480 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 9800 480 9920 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal2 s 10874 27520 10930 28000 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal3 s 0 11160 480 11280 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal2 s 12898 27520 12954 28000 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal2 s 14922 27520 14978 28000 6 chany_bottom_in[0]
port 33 nsew default input
rlabel metal2 s 18878 0 18934 480 6 chany_bottom_in[1]
port 34 nsew default input
rlabel metal3 s 0 15104 480 15224 6 chany_bottom_in[2]
port 35 nsew default input
rlabel metal3 s 0 16464 480 16584 6 chany_bottom_in[3]
port 36 nsew default input
rlabel metal3 s 0 17824 480 17944 6 chany_bottom_in[4]
port 37 nsew default input
rlabel metal2 s 16854 27520 16910 28000 6 chany_bottom_in[5]
port 38 nsew default input
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_in[6]
port 39 nsew default input
rlabel metal2 s 18878 27520 18934 28000 6 chany_bottom_in[7]
port 40 nsew default input
rlabel metal3 s 27520 18096 28000 18216 6 chany_bottom_in[8]
port 41 nsew default input
rlabel metal3 s 0 19184 480 19304 6 chany_bottom_out[0]
port 42 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_bottom_out[1]
port 43 nsew default tristate
rlabel metal2 s 22834 27520 22890 28000 6 chany_bottom_out[2]
port 44 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chany_bottom_out[3]
port 45 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chany_bottom_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chany_bottom_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chany_bottom_out[6]
port 48 nsew default tristate
rlabel metal2 s 22834 0 22890 480 6 chany_bottom_out[7]
port 49 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_bottom_out[8]
port 50 nsew default tristate
rlabel metal2 s 2870 0 2926 480 6 data_in
port 51 nsew default input
rlabel metal2 s 938 0 994 480 6 enable
port 52 nsew default input
rlabel metal3 s 0 23128 480 23248 6 left_bottom_grid_pin_12_
port 53 nsew default input
rlabel metal2 s 24858 0 24914 480 6 left_top_grid_pin_11_
port 54 nsew default input
rlabel metal2 s 26882 0 26938 480 6 left_top_grid_pin_13_
port 55 nsew default input
rlabel metal3 s 0 27208 480 27328 6 left_top_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 26882 27520 26938 28000 6 left_top_grid_pin_1_
port 57 nsew default input
rlabel metal3 s 27520 24624 28000 24744 6 left_top_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 24488 480 24608 6 left_top_grid_pin_5_
port 59 nsew default input
rlabel metal3 s 0 25848 480 25968 6 left_top_grid_pin_7_
port 60 nsew default input
rlabel metal3 s 27520 26800 28000 26920 6 left_top_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
