* NGSPICE file created from sb_2__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_dfxbp_1 abstract view
.subckt scs8hd_dfxbp_1 CLK D Q QN vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_mux2_1 abstract view
.subckt scs8hd_mux2_1 A0 A1 S X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

.subckt sb_2__1_ bottom_left_grid_pin_34_ bottom_left_grid_pin_35_ bottom_left_grid_pin_36_
+ bottom_left_grid_pin_37_ bottom_left_grid_pin_38_ bottom_left_grid_pin_39_ bottom_left_grid_pin_40_
+ bottom_left_grid_pin_41_ bottom_right_grid_pin_1_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_top_grid_pin_42_ left_top_grid_pin_43_ left_top_grid_pin_44_
+ left_top_grid_pin_45_ left_top_grid_pin_46_ left_top_grid_pin_47_ left_top_grid_pin_48_
+ left_top_grid_pin_49_ prog_clk top_left_grid_pin_34_ top_left_grid_pin_35_ top_left_grid_pin_36_
+ top_left_grid_pin_37_ top_left_grid_pin_38_ top_left_grid_pin_39_ top_left_grid_pin_40_
+ top_left_grid_pin_41_ top_right_grid_pin_1_ vpwr vgnd
XFILLER_39_222 vpwr vgnd scs8hd_fill_2
XFILLER_22_199 vgnd vpwr scs8hd_decap_12
XFILLER_22_122 vpwr vgnd scs8hd_fill_2
XFILLER_7_7 vgnd vpwr scs8hd_decap_3
Xmem_left_track_19.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_19.mux_l1_in_0_/S mux_left_track_19.mux_l2_in_0_/S
+ mem_left_track_19.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_41 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_25.scs8hd_buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X _081_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_9_126 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_2__S mux_top_track_16.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_1_ bottom_left_grid_pin_36_ bottom_left_grid_pin_34_
+ mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_67 vpwr vgnd scs8hd_fill_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XFILLER_12_43 vpwr vgnd scs8hd_fill_2
XFILLER_37_95 vgnd vpwr scs8hd_fill_1
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_15_217 vgnd vpwr scs8hd_decap_12
X_062_ _062_/A chanx_left_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_68 vpwr vgnd scs8hd_fill_2
XFILLER_9_33 vpwr vgnd scs8hd_fill_2
XFILLER_9_99 vgnd vpwr scs8hd_decap_4
Xmux_left_track_13.scs8hd_buf_4_0_ mux_left_track_13.mux_l3_in_0_/X _067_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l3_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_86 vgnd vpwr scs8hd_fill_1
XFILLER_7_224 vgnd vpwr scs8hd_decap_6
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_045_ _045_/HI _045_/LO vgnd vpwr scs8hd_conb_1
Xmem_bottom_track_3.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l4_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_172 vpwr vgnd scs8hd_fill_2
XFILLER_37_161 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_3_/S
+ mux_bottom_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l2_in_0__S mux_left_track_17.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_205 vpwr vgnd scs8hd_fill_2
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_10 vpwr vgnd scs8hd_fill_2
XFILLER_20_32 vpwr vgnd scs8hd_fill_2
XFILLER_29_30 vpwr vgnd scs8hd_fill_2
X_028_ _028_/HI _028_/LO vgnd vpwr scs8hd_conb_1
XFILLER_34_131 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_33.scs8hd_buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X _077_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_25_164 vpwr vgnd scs8hd_fill_2
XFILLER_15_32 vpwr vgnd scs8hd_fill_2
XFILLER_40_145 vgnd vpwr scs8hd_decap_8
XFILLER_40_123 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_42 vpwr vgnd scs8hd_fill_2
XFILLER_31_97 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_31_134 vpwr vgnd scs8hd_fill_2
XFILLER_31_123 vpwr vgnd scs8hd_fill_2
XFILLER_31_101 vgnd vpwr scs8hd_fill_1
XFILLER_16_120 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_7.mux_l1_in_0__S mux_left_track_7.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_145 vgnd vpwr scs8hd_decap_4
Xmem_left_track_19.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_17.mux_l2_in_0_/S mux_left_track_19.mux_l1_in_0_/S
+ mem_left_track_19.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_26_75 vpwr vgnd scs8hd_fill_2
XFILLER_13_101 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
XFILLER_13_134 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_149 vgnd vpwr scs8hd_decap_3
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_1_/S
+ mux_bottom_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__D mux_top_track_8.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_21.scs8hd_buf_4_0_ mux_left_track_21.mux_l2_in_0_/X _063_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XFILLER_23_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_15_229 vgnd vpwr scs8hd_decap_12
X_061_ _061_/A chanx_left_out[12] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A0 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_2_188 vpwr vgnd scs8hd_fill_2
XFILLER_2_166 vgnd vpwr scs8hd_fill_1
XFILLER_9_12 vpwr vgnd scs8hd_fill_2
XFILLER_9_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_1.mux_l1_in_0_/S mux_left_track_1.mux_l2_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_18_65 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_7_203 vpwr vgnd scs8hd_fill_2
XFILLER_11_221 vgnd vpwr scs8hd_decap_12
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
X_044_ _044_/HI _044_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_3__S mux_left_track_7.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__S mux_left_track_5.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l3_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_1__A0 mux_bottom_track_1.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__D mux_top_track_24.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
X_027_ _027_/HI _027_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_68 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_3_ _032_/HI left_top_grid_pin_49_ mux_left_track_7.mux_l1_in_2_/S
+ mux_left_track_7.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l4_in_0__S mux_top_track_8.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_40_135 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_21.scs8hd_dfxbp_1_0__D mux_left_track_19.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D mux_bottom_track_5.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_15.mux_l3_in_0_ mux_left_track_15.mux_l2_in_1_/X mux_left_track_15.mux_l2_in_0_/X
+ mux_left_track_15.mux_l3_in_0_/S mux_left_track_15.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l4_in_0__A0 mux_bottom_track_1.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_3_ _034_/HI chanx_left_in[14] mux_top_track_0.mux_l2_in_1_/S
+ mux_top_track_0.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_22_102 vpwr vgnd scs8hd_fill_2
XFILLER_13_157 vgnd vpwr scs8hd_decap_4
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_21.mux_l1_in_0__S mux_left_track_21.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_75 vpwr vgnd scs8hd_fill_2
XFILLER_37_53 vpwr vgnd scs8hd_fill_2
XFILLER_37_42 vpwr vgnd scs8hd_fill_2
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_1_ _051_/HI left_top_grid_pin_45_ mux_left_track_15.mux_l2_in_1_/S
+ mux_left_track_15.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.mux_l1_in_3__S mux_top_track_24.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_131 vpwr vgnd scs8hd_fill_2
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_5_197 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ mux_left_track_7.mux_l3_in_0_/S mux_left_track_7.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_060_ left_top_grid_pin_43_ chanx_left_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_4
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XFILLER_2_134 vpwr vgnd scs8hd_fill_2
XFILLER_2_112 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_2__A1 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ mux_top_track_0.mux_l4_in_0_/S mux_top_track_0.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_59 vgnd vpwr scs8hd_decap_3
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l3_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_15.scs8hd_buf_4_0__A mux_left_track_15.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__061__A _061_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_22 vpwr vgnd scs8hd_fill_2
XFILLER_18_44 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_decap_3
XFILLER_34_10 vpwr vgnd scs8hd_fill_2
Xmem_left_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_33.mux_l3_in_0_/S mux_left_track_1.mux_l1_in_0_/S
+ mem_left_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
X_112_ _112_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_34_87 vgnd vpwr scs8hd_decap_4
XFILLER_34_65 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.mux_l2_in_1_ mux_left_track_7.mux_l1_in_3_/X mux_left_track_7.mux_l1_in_2_/X
+ mux_left_track_7.mux_l2_in_1_/S mux_left_track_7.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
X_043_ _043_/HI _043_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__D mux_bottom_track_9.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_237 vgnd vpwr scs8hd_decap_6
XFILLER_11_233 vgnd vpwr scs8hd_decap_8
XFILLER_38_108 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_3.mux_l1_in_1_/S mux_bottom_track_3.mux_l2_in_0_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l3_in_1__A1 mux_bottom_track_1.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__056__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_20_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_45 vpwr vgnd scs8hd_fill_2
XFILLER_20_89 vgnd vpwr scs8hd_decap_3
XFILLER_29_87 vpwr vgnd scs8hd_fill_2
XFILLER_28_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_6 vpwr vgnd scs8hd_fill_2
XFILLER_34_144 vgnd vpwr scs8hd_decap_8
XFILLER_19_152 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.mux_l1_in_2_ left_top_grid_pin_47_ left_top_grid_pin_45_ mux_left_track_7.mux_l1_in_2_/S
+ mux_left_track_7.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_40_158 vgnd vpwr scs8hd_decap_8
XFILLER_15_12 vgnd vpwr scs8hd_decap_4
XFILLER_31_66 vgnd vpwr scs8hd_decap_3
XFILLER_31_11 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l2_in_0__S mux_left_track_13.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l4_in_0__A1 mux_bottom_track_1.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_188 vgnd vpwr scs8hd_decap_12
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_2_ chanx_left_in[7] chanx_left_in[0] mux_top_track_0.mux_l2_in_1_/S
+ mux_top_track_0.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_203 vpwr vgnd scs8hd_fill_2
XFILLER_22_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_19.mux_l1_in_1__S mux_left_track_19.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_11 vpwr vgnd scs8hd_fill_2
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_21_180 vgnd vpwr scs8hd_decap_3
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_26 vpwr vgnd scs8hd_fill_2
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XFILLER_8_140 vpwr vgnd scs8hd_fill_2
XFILLER_8_162 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_5.scs8hd_buf_4_0_ mux_bottom_track_5.mux_l4_in_0_/X _091_/A vgnd
+ vpwr scs8hd_buf_1
XANTENNA_mux_left_track_3.mux_l1_in_0__S mux_left_track_3.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_128 vgnd vpwr scs8hd_fill_1
XANTENNA__064__A _064_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_35 vpwr vgnd scs8hd_fill_2
XFILLER_12_68 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_0_ chany_bottom_in[19] mux_left_track_15.mux_l1_in_0_/X
+ mux_left_track_15.mux_l2_in_1_/S mux_left_track_15.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_154 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA__059__A chany_top_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_9.mux_l1_in_0_/S mux_left_track_9.mux_l2_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A0 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_20_212 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vpwr vgnd scs8hd_fill_2
XFILLER_18_89 vgnd vpwr scs8hd_decap_3
X_111_ _111_/A chany_top_out[2] vgnd vpwr scs8hd_buf_2
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S mux_left_track_7.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
X_042_ _042_/HI _042_/LO vgnd vpwr scs8hd_conb_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__D mux_top_track_16.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_bottom_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_1.mux_l4_in_0_/S mux_bottom_track_3.mux_l1_in_1_/S
+ mem_bottom_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_153 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_219 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _072_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vpwr vgnd scs8hd_fill_2
XFILLER_28_142 vpwr vgnd scs8hd_fill_2
XFILLER_6_26 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_32.mux_l1_in_1__S mux_top_track_32.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l3_in_1__A0 mux_top_track_0.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_34_123 vpwr vgnd scs8hd_fill_2
XFILLER_34_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_3__S mux_left_track_3.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l3_in_0__S mux_left_track_1.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_7.mux_l1_in_1_ left_top_grid_pin_43_ chany_bottom_in[6] mux_left_track_7.mux_l1_in_2_/S
+ mux_left_track_7.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_25_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 mux_bottom_track_5.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_156 vpwr vgnd scs8hd_fill_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_15_68 vpwr vgnd scs8hd_fill_2
XFILLER_31_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D mux_left_track_25.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_233 vpwr vgnd scs8hd_fill_2
XFILLER_0_222 vgnd vpwr scs8hd_decap_6
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_31_104 vgnd vpwr scs8hd_fill_1
XFILLER_16_145 vpwr vgnd scs8hd_fill_2
XFILLER_16_167 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_7.mux_l2_in_1__S mux_left_track_7.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_1_ chany_bottom_in[12] mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_1_/S
+ mux_top_track_0.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_226 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_30_181 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0__A0 chany_bottom_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_26_89 vgnd vpwr scs8hd_fill_1
XFILLER_26_45 vpwr vgnd scs8hd_fill_2
XFILLER_26_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__A0 _044_/HI vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_11 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.scs8hd_buf_4_0_ mux_left_track_9.mux_l3_in_0_/X _069_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_4.mux_l4_in_0__S mux_top_track_4.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__A0 mux_top_track_0.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_185 vpwr vgnd scs8hd_fill_2
XFILLER_12_192 vpwr vgnd scs8hd_fill_2
XFILLER_10_107 vpwr vgnd scs8hd_fill_2
XANTENNA__080__A chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_37_11 vgnd vpwr scs8hd_decap_4
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_99 vgnd vpwr scs8hd_decap_12
XFILLER_37_88 vgnd vpwr scs8hd_decap_4
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[2] top_right_grid_pin_1_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_2.scs8hd_buf_4_0_ mux_top_track_2.mux_l4_in_0_/X _112_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A0 mux_left_track_1.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XFILLER_23_79 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_23_35 vgnd vpwr scs8hd_decap_3
XANTENNA__075__A chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_2_158 vpwr vgnd scs8hd_fill_2
XFILLER_9_37 vgnd vpwr scs8hd_decap_4
XFILLER_14_210 vgnd vpwr scs8hd_decap_4
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
Xmem_left_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_7.mux_l3_in_0_/S mux_left_track_9.mux_l1_in_0_/S
+ mem_left_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_0.mux_l2_in_2__A1 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_ chany_bottom_in[12] chany_top_in[12] mux_left_track_15.mux_l1_in_0_/S
+ mux_left_track_15.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
X_110_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_34_78 vpwr vgnd scs8hd_fill_2
XFILLER_34_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
X_041_ _041_/HI _041_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l2_in_1__S mux_top_track_24.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_165 vgnd vpwr scs8hd_decap_4
XFILLER_1_71 vgnd vpwr scs8hd_decap_4
XFILLER_37_176 vpwr vgnd scs8hd_fill_2
XFILLER_4_209 vpwr vgnd scs8hd_fill_2
XFILLER_28_154 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l2_in_3_ _047_/HI chanx_left_in[18] mux_bottom_track_9.mux_l2_in_3_/S
+ mux_bottom_track_9.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l3_in_1__A1 mux_top_track_0.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_110 vpwr vgnd scs8hd_fill_2
Xmux_left_track_7.mux_l1_in_0_ chany_bottom_in[3] chany_top_in[6] mux_left_track_7.mux_l1_in_2_/S
+ mux_left_track_7.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_168 vgnd vpwr scs8hd_decap_12
XANTENNA__083__A chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_15_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_212 vpwr vgnd scs8hd_fill_2
XFILLER_0_245 vgnd vpwr scs8hd_decap_3
XFILLER_31_138 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S mux_top_track_0.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_249 vpwr vgnd scs8hd_fill_2
XFILLER_39_238 vgnd vpwr scs8hd_decap_6
XFILLER_30_193 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0__A1 mux_left_track_11.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_79 vpwr vgnd scs8hd_fill_2
XANTENNA__078__A chany_top_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__A1 mux_top_track_0.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_42_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_15.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ mux_bottom_track_9.mux_l4_in_0_/S mux_bottom_track_9.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_1_ top_left_grid_pin_40_ top_left_grid_pin_38_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0__A1 mux_left_track_1.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_3
XFILLER_4_82 vpwr vgnd scs8hd_fill_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_9_16 vpwr vgnd scs8hd_fill_2
XFILLER_13_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.scs8hd_buf_4_0__A mux_left_track_7.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S mux_bottom_track_9.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_36 vpwr vgnd scs8hd_fill_2
XFILLER_18_69 vpwr vgnd scs8hd_fill_2
XANTENNA__086__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_207 vpwr vgnd scs8hd_fill_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
Xmux_left_track_19.scs8hd_buf_4_0_ mux_left_track_19.mux_l2_in_0_/X _064_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_1_3 vgnd vpwr scs8hd_decap_4
X_040_ _040_/HI _040_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_6_240 vgnd vpwr scs8hd_fill_1
XFILLER_37_188 vgnd vpwr scs8hd_decap_12
XFILLER_37_111 vgnd vpwr scs8hd_decap_8
XFILLER_1_50 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_29_13 vpwr vgnd scs8hd_fill_2
XFILLER_28_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_5__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XFILLER_3_210 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[4] mux_bottom_track_9.mux_l2_in_3_/S
+ mux_bottom_track_9.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_133 vpwr vgnd scs8hd_fill_2
XFILLER_19_144 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_34_158 vgnd vpwr scs8hd_decap_12
XFILLER_40_117 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_3__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_23.scs8hd_buf_4_0__A mux_left_track_23.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_257 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_3
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_217 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 mux_top_track_4.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_106 vgnd vpwr scs8hd_decap_8
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_26_58 vpwr vgnd scs8hd_fill_2
XFILLER_21_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_36_209 vgnd vpwr scs8hd_decap_4
XFILLER_8_154 vgnd vpwr scs8hd_fill_1
XFILLER_12_161 vpwr vgnd scs8hd_fill_2
XFILLER_32_90 vpwr vgnd scs8hd_fill_2
XFILLER_8_165 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A mux_bottom_track_17.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_3__A0 _036_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l2_in_1__S mux_left_track_3.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l1_in_0__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_37_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA__089__A _089_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.mux_l1_in_0_ top_left_grid_pin_36_ top_left_grid_pin_34_ mux_top_track_0.mux_l1_in_0_/S
+ mux_top_track_0.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_3__S mux_top_track_2.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l4_in_0__S mux_top_track_0.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_61 vgnd vpwr scs8hd_fill_1
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_138 vpwr vgnd scs8hd_fill_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_5__A0 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l2_in_1_ _043_/HI mux_bottom_track_25.mux_l1_in_2_/X mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_81 vpwr vgnd scs8hd_fill_2
XFILLER_1_193 vgnd vpwr scs8hd_decap_3
XFILLER_1_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S mux_bottom_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_20_204 vgnd vpwr scs8hd_decap_8
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_26 vpwr vgnd scs8hd_fill_2
XFILLER_40_90 vpwr vgnd scs8hd_fill_2
X_099_ chany_bottom_in[13] chany_top_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_37_156 vgnd vpwr scs8hd_fill_1
XFILLER_37_134 vgnd vpwr scs8hd_decap_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l1_in_2__A0 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l2_in_1__A0 _050_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_49 vpwr vgnd scs8hd_fill_2
XFILLER_28_134 vgnd vpwr scs8hd_decap_6
XFILLER_28_101 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__097__A _097_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_178 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_25.mux_l1_in_2_ chanx_left_in[13] chanx_left_in[6] mux_bottom_track_25.mux_l1_in_2_/S
+ mux_bottom_track_25.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
XFILLER_3_233 vpwr vgnd scs8hd_fill_2
XFILLER_3_222 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_1_ bottom_left_grid_pin_41_ bottom_left_grid_pin_37_
+ mux_bottom_track_9.mux_l2_in_3_/S mux_bottom_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 bottom_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vgnd vpwr scs8hd_fill_1
XFILLER_0_269 vgnd vpwr scs8hd_decap_8
XFILLER_16_137 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_207 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_3.mux_l2_in_1__A0 mux_left_track_3.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l3_in_0__A0 mux_left_track_13.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_11_6 vpwr vgnd scs8hd_fill_2
XFILLER_22_118 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__D mux_bottom_track_33.mux_l2_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_23.mux_l1_in_0__A0 chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_7_83 vpwr vgnd scs8hd_fill_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_129 vgnd vpwr scs8hd_decap_3
XFILLER_21_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_16_70 vpwr vgnd scs8hd_fill_2
XFILLER_8_144 vpwr vgnd scs8hd_fill_2
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_3__A1 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l1_in_0__A1 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_37_36 vgnd vpwr scs8hd_decap_4
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A0 mux_left_track_3.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A mux_bottom_track_5.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_4_40 vgnd vpwr scs8hd_decap_4
XFILLER_4_180 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__D mux_left_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_5__A1 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_29_7 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_2__S mux_bottom_track_25.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_48 vpwr vgnd scs8hd_fill_2
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
X_098_ chany_bottom_in[14] chany_top_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_1_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_2__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l2_in_1__A1 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_29_26 vpwr vgnd scs8hd_fill_2
XFILLER_28_146 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_25.mux_l1_in_1_ bottom_left_grid_pin_39_ bottom_left_grid_pin_35_
+ mux_bottom_track_25.mux_l1_in_2_/S mux_bottom_track_25.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_ bottom_right_grid_pin_1_ mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_3_/S mux_bottom_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_127 vpwr vgnd scs8hd_fill_2
XFILLER_34_116 vgnd vpwr scs8hd_decap_4
XFILLER_19_81 vgnd vpwr scs8hd_decap_4
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_31_49 vpwr vgnd scs8hd_fill_2
XFILLER_31_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_237 vgnd vpwr scs8hd_decap_8
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 mux_left_track_3.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l3_in_0__A1 mux_left_track_13.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_3_ _035_/HI chanx_left_in[17] mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_23.mux_l1_in_0__A1 chany_top_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_38_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__D mux_left_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 mux_top_track_24.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_196 vgnd vpwr scs8hd_decap_12
XFILLER_21_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_3__S mux_bottom_track_5.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l4_in_0__S mux_bottom_track_3.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XFILLER_8_189 vpwr vgnd scs8hd_fill_2
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_12_196 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_3__A0 _042_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_1__S mux_bottom_track_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__A1 mux_left_track_3.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.scs8hd_buf_4_0__A mux_top_track_0.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D mux_bottom_track_9.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_11.scs8hd_dfxbp_1_2__D mux_left_track_11.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_74 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_9 vpwr vgnd scs8hd_fill_2
XFILLER_2_107 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 top_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__S mux_left_track_5.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_3_ _030_/HI left_top_grid_pin_49_ mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_5__A0 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l1_in_1__A0 chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_17.mux_l1_in_1_/S mux_left_track_17.mux_l2_in_0_/S
+ mem_left_track_17.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_4.mux_l1_in_4__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_1__S mux_top_track_2.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
XFILLER_6_210 vgnd vpwr scs8hd_fill_1
XFILLER_41_7 vpwr vgnd scs8hd_fill_2
X_097_ _097_/A chany_top_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_9.mux_l2_in_0__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_6 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l3_in_0_ mux_left_track_11.mux_l2_in_1_/X mux_left_track_11.mux_l2_in_0_/X
+ mux_left_track_11.mux_l3_in_0_/S mux_left_track_11.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_16.mux_l2_in_1_ mux_top_track_16.mux_l1_in_3_/X mux_top_track_16.mux_l1_in_2_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_2__S mux_top_track_8.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D mux_left_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_2_/S
+ mux_bottom_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D mux_top_track_24.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_19_71 vgnd vpwr scs8hd_decap_4
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_35_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 mux_top_track_32.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1__A0 _052_/HI vgnd vpwr scs8hd_diode_2
XFILLER_0_216 vgnd vpwr scs8hd_fill_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__D mux_left_track_13.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_11.mux_l2_in_1_ _049_/HI left_top_grid_pin_43_ mux_left_track_11.mux_l2_in_1_/S
+ mux_left_track_11.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_16.mux_l1_in_2_ chanx_left_in[10] chanx_left_in[3] mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ mux_left_track_3.mux_l3_in_0_/S mux_left_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_0_/S
+ mux_bottom_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_16_83 vpwr vgnd scs8hd_fill_2
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l3_in_0__S mux_top_track_32.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_3__A1 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A0 mux_left_track_17.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A0 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_1.mux_l3_in_1_/S mux_bottom_track_1.mux_l4_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A0 _047_/HI vgnd vpwr scs8hd_diode_2
XFILLER_5_116 vgnd vpwr scs8hd_decap_4
XFILLER_5_127 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_82 vpwr vgnd scs8hd_fill_2
XFILLER_27_71 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D mux_top_track_0.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_4_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l1_in_3__A0 _031_/HI vgnd vpwr scs8hd_diode_2
XFILLER_4_86 vgnd vpwr scs8hd_decap_3
XFILLER_4_64 vgnd vpwr scs8hd_fill_1
Xmem_top_track_4.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_4.mux_l3_in_1_/S mux_top_track_4.mux_l4_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_top_track_8.scs8hd_buf_4_0_ mux_top_track_8.mux_l4_in_0_/X _109_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_left_track_7.mux_l2_in_0__A0 mux_left_track_7.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_51 vgnd vpwr scs8hd_decap_4
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_95 vgnd vpwr scs8hd_decap_4
XFILLER_38_81 vgnd vpwr scs8hd_decap_8
XANTENNA__100__A chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l1_in_2_ left_top_grid_pin_47_ left_top_grid_pin_45_ mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_1__A1 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_5__A1 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_15.mux_l3_in_0_/S mux_left_track_17.mux_l1_in_1_/S
+ mem_left_track_17.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A mux_bottom_track_25.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_50 vgnd vpwr scs8hd_fill_1
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
X_096_ chany_bottom_in[16] chany_top_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__D mux_left_track_13.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A0 _029_/HI vgnd vpwr scs8hd_diode_2
XFILLER_1_54 vgnd vpwr scs8hd_fill_1
XFILLER_1_98 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_5.mux_l1_in_6_ chanx_left_in[17] chanx_left_in[10] mux_bottom_track_5.mux_l1_in_6_/S
+ mux_bottom_track_5.mux_l1_in_6_/X vgnd vpwr scs8hd_mux2_1
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_3_214 vpwr vgnd scs8hd_fill_2
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_23.mux_l2_in_0__S mux_left_track_23.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_50 vgnd vpwr scs8hd_decap_3
XFILLER_19_137 vpwr vgnd scs8hd_fill_2
XFILLER_19_148 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_079_ chany_top_in[13] chany_bottom_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_19 vpwr vgnd scs8hd_fill_2
XFILLER_18_181 vgnd vpwr scs8hd_decap_3
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_228 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_0__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A0 mux_left_track_25.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_11.mux_l2_in_0_ chany_bottom_in[11] mux_left_track_11.mux_l1_in_0_/X
+ mux_left_track_11.mux_l2_in_1_/S mux_left_track_11.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[17] chany_bottom_in[8] mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__D mux_top_track_0.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_121 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_140 vpwr vgnd scs8hd_fill_2
XFILLER_7_31 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_38_232 vgnd vpwr scs8hd_decap_12
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__D mux_left_track_7.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XFILLER_8_136 vpwr vgnd scs8hd_fill_2
XFILLER_12_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_165 vpwr vgnd scs8hd_fill_2
XFILLER_16_40 vgnd vpwr scs8hd_decap_4
XFILLER_8_158 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA__103__A chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0__A1 mux_left_track_17.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.scs8hd_buf_4_0__A mux_top_track_8.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l3_in_1_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_50 vgnd vpwr scs8hd_decap_4
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_3__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_1_/S
+ mem_top_track_4.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_7.mux_l2_in_0__A1 mux_left_track_7.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l3_in_1__S mux_bottom_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_85 vgnd vpwr scs8hd_decap_4
XFILLER_1_175 vpwr vgnd scs8hd_fill_2
XFILLER_9_242 vpwr vgnd scs8hd_fill_2
Xmux_left_track_3.mux_l1_in_1_ left_top_grid_pin_43_ chany_bottom_in[4] mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_095_ chany_bottom_in[17] chany_top_out[18] vgnd vpwr scs8hd_buf_2
XFILLER_40_61 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l3_in_0__S mux_left_track_15.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_84 vpwr vgnd scs8hd_fill_2
XFILLER_6_245 vgnd vpwr scs8hd_decap_12
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__D mux_top_track_2.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__S mux_bottom_track_17.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D mux_left_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_237 vgnd vpwr scs8hd_decap_6
XFILLER_3_226 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_5_ chanx_left_in[3] bottom_left_grid_pin_41_ mux_bottom_track_5.mux_l1_in_6_/S
+ mux_bottom_track_5.mux_l1_in_5_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_53 vgnd vpwr scs8hd_fill_1
XFILLER_35_94 vgnd vpwr scs8hd_decap_4
XFILLER_35_50 vgnd vpwr scs8hd_decap_3
XANTENNA__106__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
X_078_ chany_top_in[14] chany_bottom_out[15] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_5.mux_l2_in_0__S mux_left_track_5.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_19 vpwr vgnd scs8hd_fill_2
XFILLER_0_218 vpwr vgnd scs8hd_fill_2
XFILLER_24_163 vgnd vpwr scs8hd_decap_12
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_25.mux_l2_in_0__A1 mux_left_track_25.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_96 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_2__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_ top_left_grid_pin_39_ top_left_grid_pin_35_ mux_top_track_16.mux_l1_in_0_/S
+ mux_top_track_16.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_152 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_left_track_7.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_7.mux_l2_in_1_/S mux_left_track_7.mux_l3_in_0_/S
+ mem_left_track_7.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_13.scs8hd_buf_4_0__A mux_left_track_13.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_87 vpwr vgnd scs8hd_fill_2
XFILLER_38_244 vgnd vpwr scs8hd_decap_12
XFILLER_38_200 vgnd vpwr scs8hd_decap_12
XFILLER_26_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_9.mux_l3_in_1_/S mux_bottom_track_9.mux_l4_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_32_73 vpwr vgnd scs8hd_fill_2
XFILLER_32_51 vpwr vgnd scs8hd_fill_2
XFILLER_8_148 vgnd vpwr scs8hd_decap_3
XFILLER_12_111 vgnd vpwr scs8hd_decap_3
XFILLER_12_144 vpwr vgnd scs8hd_fill_2
XFILLER_12_188 vpwr vgnd scs8hd_fill_2
XFILLER_32_84 vgnd vpwr scs8hd_decap_4
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_1.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l2_in_0_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_11.mux_l1_in_0_ chany_bottom_in[9] chany_top_in[9] mux_left_track_11.mux_l1_in_0_/S
+ mux_left_track_11.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_3__A0 _040_/HI vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
Xmux_left_track_23.mux_l2_in_0_ mux_left_track_23.mux_l1_in_1_/X mux_left_track_23.mux_l1_in_0_/X
+ mux_left_track_23.mux_l2_in_0_/S mux_left_track_23.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_17_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__D mux_top_track_4.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_99 vpwr vgnd scs8hd_fill_2
XFILLER_4_11 vgnd vpwr scs8hd_fill_1
XFILLER_4_162 vgnd vpwr scs8hd_fill_1
Xmem_top_track_4.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_1_/S
+ mem_top_track_4.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_13_20 vgnd vpwr scs8hd_fill_1
XFILLER_1_198 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_5.mux_l2_in_3_ _046_/HI mux_bottom_track_5.mux_l1_in_6_/X mux_bottom_track_5.mux_l2_in_3_/S
+ mux_bottom_track_5.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_210 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l1_in_0_ chany_bottom_in[0] chany_top_in[4] mux_left_track_3.mux_l1_in_1_/S
+ mux_left_track_3.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_7.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_209 vgnd vpwr scs8hd_decap_12
Xmux_left_track_23.mux_l1_in_1_ _028_/HI left_top_grid_pin_49_ mux_left_track_23.mux_l1_in_1_/S
+ mux_left_track_23.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_9 vpwr vgnd scs8hd_fill_2
XFILLER_24_74 vpwr vgnd scs8hd_fill_2
X_094_ chany_bottom_in[18] chany_top_out[19] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_6_213 vgnd vpwr scs8hd_fill_1
XFILLER_6_224 vgnd vpwr scs8hd_decap_12
XFILLER_6_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__D mux_left_track_19.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_34 vgnd vpwr scs8hd_decap_4
XFILLER_28_128 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.scs8hd_buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X _093_/A vgnd
+ vpwr scs8hd_buf_1
Xmux_bottom_track_5.mux_l1_in_4_ bottom_left_grid_pin_40_ bottom_left_grid_pin_39_
+ mux_bottom_track_5.mux_l1_in_6_/S mux_bottom_track_5.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_106 vpwr vgnd scs8hd_fill_2
XFILLER_35_73 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vpwr vgnd scs8hd_fill_2
X_077_ _077_/A chany_bottom_out[16] vgnd vpwr scs8hd_buf_2
XFILLER_33_142 vpwr vgnd scs8hd_fill_2
XFILLER_0_208 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ mux_bottom_track_5.mux_l4_in_0_/S mux_bottom_track_5.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_175 vgnd vpwr scs8hd_decap_12
XFILLER_24_131 vgnd vpwr scs8hd_decap_6
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_75 vpwr vgnd scs8hd_fill_2
XFILLER_21_53 vpwr vgnd scs8hd_fill_2
XFILLER_21_31 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_175 vpwr vgnd scs8hd_fill_2
Xmem_left_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_25.mux_l1_in_0_/S ccff_tail
+ mem_left_track_25.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_145 vgnd vpwr scs8hd_decap_8
Xmem_left_track_7.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_7.mux_l1_in_2_/S mux_left_track_7.mux_l2_in_1_/S
+ mem_left_track_7.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_38_256 vgnd vpwr scs8hd_decap_12
XFILLER_38_212 vpwr vgnd scs8hd_fill_2
XFILLER_42_19 vpwr vgnd scs8hd_fill_2
XFILLER_21_145 vpwr vgnd scs8hd_fill_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l2_in_1__S mux_bottom_track_33.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__A0 _033_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D mux_bottom_track_3.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_9.mux_l2_in_3_/S mux_bottom_track_9.mux_l3_in_1_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_25.mux_l1_in_1__S mux_left_track_25.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l1_in_0__S mux_left_track_13.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_bottom_track_1.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_32.mux_l3_in_0_/S mux_bottom_track_1.mux_l1_in_1_/S
+ mem_bottom_track_1.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XFILLER_5_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_3__A1 chanx_left_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_3__S mux_top_track_16.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_78 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l3_in_0__A0 mux_left_track_9.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_4.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_2.mux_l4_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ mem_top_track_4.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_1_144 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_2_ mux_bottom_track_5.mux_l1_in_5_/X mux_bottom_track_5.mux_l1_in_4_/X
+ mux_bottom_track_5.mux_l2_in_3_/S mux_bottom_track_5.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_222 vgnd vpwr scs8hd_decap_12
Xmux_left_track_23.mux_l1_in_0_ chany_bottom_in[17] chany_top_in[17] mux_left_track_23.mux_l1_in_1_/S
+ mux_left_track_23.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_39_192 vpwr vgnd scs8hd_fill_2
XFILLER_40_41 vgnd vpwr scs8hd_decap_3
X_093_ _093_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_236 vgnd vpwr scs8hd_decap_4
XFILLER_6_269 vgnd vpwr scs8hd_decap_6
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l3_in_1__S mux_bottom_track_1.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.scs8hd_buf_4_0_ mux_left_track_5.mux_l3_in_0_/X _071_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D mux_top_track_4.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_173 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.mux_l1_in_3_ bottom_left_grid_pin_38_ bottom_left_grid_pin_37_
+ mux_bottom_track_5.mux_l1_in_6_/S mux_bottom_track_5.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__D mux_bottom_track_5.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_77 vpwr vgnd scs8hd_fill_2
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_27_151 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XFILLER_32_7 vpwr vgnd scs8hd_fill_2
X_076_ chany_top_in[16] chany_bottom_out[17] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_11.mux_l3_in_0__S mux_left_track_11.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_140 vpwr vgnd scs8hd_fill_2
XFILLER_33_154 vgnd vpwr scs8hd_decap_12
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_187 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_30_113 vpwr vgnd scs8hd_fill_2
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_132 vpwr vgnd scs8hd_fill_2
Xmem_left_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_23.mux_l2_in_0_/S mux_left_track_25.mux_l1_in_0_/S
+ mem_left_track_25.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_157 vgnd vpwr scs8hd_decap_12
Xmem_left_track_7.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_5.mux_l3_in_0_/S mux_left_track_7.mux_l1_in_2_/S
+ mem_left_track_7.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A mux_bottom_track_33.mux_l3_in_0_/X
+ vgnd vpwr scs8hd_diode_2
X_059_ chany_top_in[19] chanx_left_out[14] vgnd vpwr scs8hd_buf_2
XFILLER_38_268 vgnd vpwr scs8hd_decap_6
XFILLER_21_168 vpwr vgnd scs8hd_fill_2
XFILLER_21_113 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_0__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_9.mux_l1_in_0_/S mux_bottom_track_9.mux_l2_in_3_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_102 vgnd vpwr scs8hd_decap_3
XFILLER_12_135 vgnd vpwr scs8hd_decap_3
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_fill_1
XFILLER_16_87 vgnd vpwr scs8hd_decap_3
XFILLER_32_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_2__S mux_top_track_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__S mux_left_track_7.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_86 vpwr vgnd scs8hd_fill_2
XFILLER_27_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_4_120 vpwr vgnd scs8hd_fill_2
XFILLER_4_57 vgnd vpwr scs8hd_decap_4
XFILLER_4_46 vpwr vgnd scs8hd_fill_2
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_3__D mux_top_track_8.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l3_in_0__A1 mux_left_track_9.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D mux_bottom_track_17.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_44 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_123 vpwr vgnd scs8hd_fill_2
XFILLER_38_96 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_3_/S mux_bottom_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_234 vgnd vpwr scs8hd_decap_8
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_241 vgnd vpwr scs8hd_decap_3
XFILLER_24_98 vpwr vgnd scs8hd_fill_2
XFILLER_24_43 vgnd vpwr scs8hd_fill_1
XFILLER_24_10 vpwr vgnd scs8hd_fill_2
XFILLER_10_200 vgnd vpwr scs8hd_fill_1
XFILLER_10_211 vgnd vpwr scs8hd_decap_3
X_092_ _092_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_37_119 vgnd vpwr scs8hd_fill_1
XFILLER_36_185 vgnd vpwr scs8hd_decap_12
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_36_ bottom_left_grid_pin_35_
+ mux_bottom_track_5.mux_l1_in_6_/S mux_bottom_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_12 vgnd vpwr scs8hd_decap_4
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_45 vpwr vgnd scs8hd_fill_2
XFILLER_35_31 vgnd vpwr scs8hd_decap_4
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_163 vgnd vpwr scs8hd_decap_12
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_075_ chany_top_in[17] chany_bottom_out[18] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_24.mux_l1_in_1__S mux_top_track_24.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_7 vgnd vpwr scs8hd_decap_4
XFILLER_33_166 vgnd vpwr scs8hd_decap_12
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__D mux_top_track_32.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_169 vgnd vpwr scs8hd_decap_12
XFILLER_30_125 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.scs8hd_buf_4_0__A mux_left_track_5.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_058_ chany_top_in[15] chanx_left_out[15] vgnd vpwr scs8hd_buf_2
XFILLER_7_35 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_9.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_5.mux_l4_in_0_/S mux_bottom_track_9.mux_l1_in_0_/S
+ mem_bottom_track_9.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__D mux_left_track_21.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_107 vgnd vpwr scs8hd_decap_3
XFILLER_16_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_180 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.scs8hd_buf_4_0_ mux_left_track_15.mux_l3_in_0_/X _066_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_7_140 vgnd vpwr scs8hd_fill_1
XFILLER_11_180 vgnd vpwr scs8hd_fill_1
XFILLER_7_162 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ mux_bottom_track_33.mux_l3_in_0_/S mux_bottom_track_33.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA__054__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_27_54 vgnd vpwr scs8hd_fill_1
XFILLER_27_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_40_231 vgnd vpwr scs8hd_decap_12
XFILLER_4_36 vpwr vgnd scs8hd_fill_2
XFILLER_4_165 vpwr vgnd scs8hd_fill_2
XFILLER_4_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_21.mux_l1_in_1__S mux_left_track_21.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_21.scs8hd_buf_4_0__A mux_left_track_21.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_12 vpwr vgnd scs8hd_fill_2
XFILLER_1_102 vpwr vgnd scs8hd_fill_2
XFILLER_38_20 vpwr vgnd scs8hd_fill_2
XFILLER_1_179 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_3_/S mux_bottom_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_bottom_track_33.mux_l2_in_1_ _045_/HI mux_bottom_track_33.mux_l1_in_2_/X mux_bottom_track_33.mux_l2_in_1_/S
+ mux_bottom_track_33.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 chany_bottom_in[12] vgnd vpwr scs8hd_diode_2
XFILLER_40_10 vpwr vgnd scs8hd_fill_2
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
X_091_ _091_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_40_65 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__S mux_top_track_16.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_197 vgnd vpwr scs8hd_decap_12
XFILLER_36_142 vpwr vgnd scs8hd_fill_2
XANTENNA__062__A _062_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l1_in_1_ bottom_left_grid_pin_34_ bottom_right_grid_pin_1_
+ mux_bottom_track_5.mux_l1_in_6_/S mux_bottom_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__D mux_left_track_21.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_33.mux_l1_in_2_ chanx_left_in[14] chanx_left_in[7] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_33 vpwr vgnd scs8hd_fill_2
XFILLER_19_55 vgnd vpwr scs8hd_decap_4
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_175 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_11.mux_l1_in_0__A0 chany_bottom_in[9] vgnd vpwr scs8hd_diode_2
X_074_ chany_top_in[18] chany_bottom_out[19] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_164 vpwr vgnd scs8hd_fill_2
XFILLER_18_186 vgnd vpwr scs8hd_decap_12
XFILLER_33_178 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XANTENNA__057__A chany_top_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_24_145 vpwr vgnd scs8hd_fill_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_23.scs8hd_buf_4_0_ mux_left_track_23.mux_l2_in_0_/X _062_/A vgnd vpwr
+ scs8hd_buf_1
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_2__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_057_ chany_top_in[11] chanx_left_out[16] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_38_226 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_32_55 vgnd vpwr scs8hd_decap_4
XFILLER_32_22 vgnd vpwr scs8hd_decap_3
XFILLER_32_11 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_8_119 vgnd vpwr scs8hd_decap_4
XFILLER_12_148 vpwr vgnd scs8hd_fill_2
XFILLER_32_77 vpwr vgnd scs8hd_fill_2
XFILLER_20_192 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_1__S mux_left_track_13.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_109_ _109_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XANTENNA__070__A _070_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 top_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_40_243 vgnd vpwr scs8hd_decap_12
XFILLER_4_133 vpwr vgnd scs8hd_fill_2
XFILLER_4_199 vpwr vgnd scs8hd_fill_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_1__S mux_left_track_3.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_1__A0 mux_bottom_track_3.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__065__A _065_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_76 vgnd vpwr scs8hd_decap_3
XFILLER_38_54 vgnd vpwr scs8hd_decap_3
XFILLER_38_32 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_1_/S mux_bottom_track_33.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 mux_top_track_0.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_23 vpwr vgnd scs8hd_fill_2
XFILLER_24_78 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
X_090_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_206 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_3.mux_l4_in_0__A0 mux_bottom_track_3.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_38 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_39_3 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_6_/S
+ mux_bottom_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A mux_bottom_track_3.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_33.mux_l1_in_1_ chanx_left_in[0] bottom_left_grid_pin_40_ mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_77 vpwr vgnd scs8hd_fill_2
XFILLER_35_55 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l1_in_0__A1 chany_top_in[9] vgnd vpwr scs8hd_diode_2
X_073_ _073_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_146 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_2__D mux_top_track_16.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_fill_1
XFILLER_18_198 vgnd vpwr scs8hd_decap_12
XFILLER_24_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_79 vpwr vgnd scs8hd_fill_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
XFILLER_21_35 vpwr vgnd scs8hd_fill_2
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l1_in_2__S mux_top_track_32.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
X_056_ chany_top_in[7] chanx_left_out[17] vgnd vpwr scs8hd_buf_2
XFILLER_30_7 vpwr vgnd scs8hd_fill_2
XFILLER_23_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l1_in_3_ _037_/HI chanx_left_in[16] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_0__A1 chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_46 vgnd vpwr scs8hd_fill_1
Xmem_left_track_15.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_15.mux_l2_in_1_/S mux_left_track_15.mux_l3_in_0_/S
+ mem_left_track_15.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_3.mux_l2_in_2__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
X_108_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_11_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
X_039_ _039_/HI _039_/LO vgnd vpwr scs8hd_conb_1
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_12 vpwr vgnd scs8hd_fill_2
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_40_255 vgnd vpwr scs8hd_decap_12
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l3_in_1__A1 mux_bottom_track_3.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_211 vgnd vpwr scs8hd_decap_3
XANTENNA__081__A _081_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_148 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_5_81 vpwr vgnd scs8hd_fill_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_3
XFILLER_24_46 vpwr vgnd scs8hd_fill_2
XFILLER_24_35 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_10_203 vgnd vpwr scs8hd_decap_8
XFILLER_40_78 vgnd vpwr scs8hd_decap_12
XFILLER_40_23 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l2_in_3_ _036_/HI chanx_left_in[13] mux_top_track_2.mux_l2_in_1_/S
+ mux_top_track_2.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l4_in_0__A1 mux_bottom_track_3.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_111 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.mux_l2_in_1_ mux_top_track_24.mux_l1_in_3_/X mux_top_track_24.mux_l1_in_2_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_19_46 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_33.mux_l1_in_0_ bottom_left_grid_pin_36_ chany_top_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_221 vgnd vpwr scs8hd_decap_8
X_072_ _072_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_114 vpwr vgnd scs8hd_fill_2
XFILLER_18_144 vgnd vpwr scs8hd_decap_3
XFILLER_24_114 vgnd vpwr scs8hd_decap_8
XFILLER_2_93 vpwr vgnd scs8hd_fill_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ mux_left_track_9.mux_l3_in_0_/S mux_left_track_9.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XFILLER_30_117 vpwr vgnd scs8hd_fill_2
XFILLER_30_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_136 vpwr vgnd scs8hd_fill_2
X_055_ chany_top_in[3] chanx_left_out[18] vgnd vpwr scs8hd_buf_2
Xmux_top_track_24.mux_l1_in_2_ chanx_left_in[9] chanx_left_in[2] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XFILLER_21_128 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ mux_top_track_2.mux_l4_in_0_/S mux_top_track_2.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_16_36 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_3
Xmem_left_track_15.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_15.mux_l1_in_0_/S mux_left_track_15.mux_l2_in_1_/S
+ mem_left_track_15.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__084__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_150 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_107_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_7_110 vpwr vgnd scs8hd_fill_2
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_11_172 vpwr vgnd scs8hd_fill_2
X_038_ _038_/HI _038_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_2.mux_l2_in_2__A0 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_1_ _033_/HI left_top_grid_pin_42_ mux_left_track_9.mux_l2_in_0_/S
+ mux_left_track_9.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_40_267 vgnd vpwr scs8hd_decap_8
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_3__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_38_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_4__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_1__A0 mux_top_track_2.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_201 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_0_171 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_2__S mux_bottom_track_17.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_175 vpwr vgnd scs8hd_fill_2
XFILLER_39_142 vpwr vgnd scs8hd_fill_2
XFILLER_39_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_19.mux_l2_in_0__S mux_left_track_19.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_40_46 vgnd vpwr scs8hd_decap_6
XANTENNA__092__A _092_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l2_in_2_ chanx_left_in[6] chany_bottom_in[13] mux_top_track_2.mux_l2_in_1_/S
+ mux_top_track_2.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
Xmem_bottom_track_17.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_17.mux_l2_in_0_/S
+ mux_bottom_track_17.mux_l3_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0__A0 chany_bottom_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_10_16 vgnd vpwr scs8hd_fill_1
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_10_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_3__A0 _046_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l4_in_0__A0 mux_top_track_2.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_3
XANTENNA__087__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
X_071_ _071_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_2_233 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_18_123 vgnd vpwr scs8hd_fill_1
XFILLER_41_181 vpwr vgnd scs8hd_fill_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_9.mux_l1_in_0__S mux_left_track_9.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_2.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l4_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ mux_left_track_17.mux_l2_in_0_/S mux_left_track_17.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l1_in_3__A0 _048_/HI vgnd vpwr scs8hd_diode_2
XFILLER_23_170 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_6__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_148 vpwr vgnd scs8hd_fill_2
X_054_ chany_top_in[1] chanx_left_out[19] vgnd vpwr scs8hd_buf_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_3
XFILLER_38_218 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_3.mux_l2_in_0__A0 mux_left_track_3.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.scs8hd_buf_4_0_ mux_top_track_4.mux_l4_in_0_/X _111_/A vgnd vpwr
+ scs8hd_buf_1
Xmux_top_track_24.mux_l1_in_1_ chany_bottom_in[18] chany_bottom_in[9] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 top_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XFILLER_14_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
Xmem_left_track_15.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_13.mux_l3_in_0_/S mux_left_track_15.mux_l1_in_0_/S
+ mem_left_track_15.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_12_107 vpwr vgnd scs8hd_fill_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_3_ _041_/HI chanx_left_in[15] mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
X_106_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
Xmux_left_track_17.mux_l1_in_1_ _052_/HI left_top_grid_pin_46_ mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_037_ _037_/HI _037_/LO vgnd vpwr scs8hd_conb_1
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.mux_l2_in_0_ chany_bottom_in[8] mux_left_track_9.mux_l1_in_0_/X
+ mux_left_track_9.mux_l2_in_0_/S mux_left_track_9.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_2__A1 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_21.mux_l1_in_1__A0 _027_/HI vgnd vpwr scs8hd_diode_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A chany_bottom_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_4_103 vpwr vgnd scs8hd_fill_2
XFILLER_4_29 vpwr vgnd scs8hd_fill_2
XFILLER_4_158 vgnd vpwr scs8hd_decap_4
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_13_16 vpwr vgnd scs8hd_fill_2
XFILLER_1_106 vpwr vgnd scs8hd_fill_2
XFILLER_38_24 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_5.mux_l1_in_4__A1 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_1__A1 mux_top_track_2.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_21.mux_l2_in_0__A0 mux_left_track_21.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l3_in_0__S mux_left_track_7.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D mux_bottom_track_25.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_154 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ mux_bottom_track_1.mux_l4_in_0_/S mux_bottom_track_1.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l2_in_1_ chany_bottom_in[4] top_left_grid_pin_41_ mux_top_track_2.mux_l2_in_1_/S
+ mux_top_track_2.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_80 vgnd vpwr scs8hd_decap_6
XFILLER_36_146 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_17.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_17.mux_l1_in_3_/S
+ mux_bottom_track_17.mux_l2_in_0_/S mem_bottom_track_17.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l2_in_0__A1 mux_left_track_13.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_3__A1 mux_bottom_track_5.mux_l1_in_6_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l4_in_0__A1 mux_top_track_2.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
X_070_ _070_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_245 vgnd vpwr scs8hd_decap_12
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_18_168 vpwr vgnd scs8hd_fill_2
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_91 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_2.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_2.mux_l2_in_1_/S mux_top_track_2.mux_l3_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_2_84 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S mux_bottom_track_1.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_13.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D mux_bottom_track_33.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_3__A1 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_15_116 vgnd vpwr scs8hd_decap_4
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
X_053_ _053_/HI _053_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_23.mux_l1_in_0__S mux_left_track_23.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l2_in_0__A1 mux_left_track_3.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_24.mux_l1_in_0_ top_left_grid_pin_40_ top_left_grid_pin_36_ mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vpwr vgnd scs8hd_fill_2
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
X_105_ _105_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_1.mux_l2_in_2_ chanx_left_in[8] chanx_left_in[1] mux_bottom_track_1.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_11_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_24.mux_l3_in_0__S mux_top_track_24.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_ chany_bottom_in[13] chany_top_in[13] mux_left_track_17.mux_l1_in_1_/S
+ mux_left_track_17.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A0 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
X_036_ _036_/HI _036_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_8_50 vgnd vpwr scs8hd_decap_3
XFILLER_8_72 vpwr vgnd scs8hd_fill_2
XFILLER_8_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_21.mux_l1_in_1__A1 left_top_grid_pin_48_ vgnd vpwr scs8hd_diode_2
XFILLER_4_137 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_16_200 vgnd vpwr scs8hd_decap_12
XFILLER_17_81 vpwr vgnd scs8hd_fill_2
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_91 vpwr vgnd scs8hd_fill_2
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_38_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A0 mux_bottom_track_17.mux_l1_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l1_in_0_ chany_bottom_in[7] chany_top_in[8] mux_left_track_9.mux_l1_in_0_/S
+ mux_left_track_9.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l3_in_0_/S
+ mem_left_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_21.mux_l2_in_0__A1 mux_left_track_21.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.scs8hd_buf_4_0__A mux_left_track_11.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_40 vpwr vgnd scs8hd_fill_2
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_39_166 vgnd vpwr scs8hd_fill_1
XFILLER_39_188 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_4__A0 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l2_in_0_ top_left_grid_pin_39_ mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S mux_top_track_2.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_14_71 vpwr vgnd scs8hd_fill_2
XFILLER_5_210 vpwr vgnd scs8hd_fill_2
XFILLER_5_221 vpwr vgnd scs8hd_fill_2
XFILLER_5_243 vgnd vpwr scs8hd_fill_1
XFILLER_39_7 vpwr vgnd scs8hd_fill_2
XFILLER_36_125 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_17.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_9.mux_l4_in_0_/S
+ mux_bottom_track_17.mux_l1_in_3_/S mem_bottom_track_17.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A0 mux_bottom_track_17.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_27_103 vgnd vpwr scs8hd_decap_6
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_35_37 vpwr vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_11.scs8hd_dfxbp_1_0__D mux_left_track_9.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 top_left_grid_pin_36_ vgnd vpwr scs8hd_diode_2
XFILLER_2_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0__S mux_left_track_15.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_136 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_2.mux_l1_in_0_/S mux_top_track_2.mux_l2_in_1_/S
+ mem_top_track_2.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_4.mux_l2_in_3__A0 _039_/HI vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S mux_bottom_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_24_139 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_21_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A0 chanx_left_in[13] vgnd vpwr scs8hd_diode_2
X_052_ _052_/HI _052_/LO vgnd vpwr scs8hd_conb_1
XFILLER_36_91 vgnd vpwr scs8hd_fill_1
XFILLER_21_109 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__S mux_left_track_5.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_231 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
X_104_ chany_bottom_in[8] chany_top_out[9] vgnd vpwr scs8hd_buf_2
XFILLER_22_82 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_1_ bottom_left_grid_pin_41_ mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_168 vgnd vpwr scs8hd_decap_3
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
X_035_ _035_/HI _035_/LO vgnd vpwr scs8hd_conb_1
XFILLER_11_197 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l1_in_0__A0 chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A1 chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XFILLER_27_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 _043_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_2__D mux_left_track_3.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_4_149 vpwr vgnd scs8hd_fill_2
XFILLER_4_116 vpwr vgnd scs8hd_fill_2
XFILLER_16_212 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_193 vpwr vgnd scs8hd_fill_2
XFILLER_3_160 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l2_in_1__A0 _051_/HI vgnd vpwr scs8hd_diode_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_39_ bottom_left_grid_pin_37_
+ mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A1 mux_bottom_track_17.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_1__A0 mux_bottom_track_9.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
Xmem_left_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_5.mux_l1_in_3_/S mux_left_track_5.mux_l2_in_1_/S
+ mem_left_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_left_track_23.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_23.mux_l1_in_1_/S mux_left_track_23.mux_l2_in_0_/S
+ mem_left_track_23.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.scs8hd_buf_4_0__A mux_top_track_16.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_85 vpwr vgnd scs8hd_fill_2
XFILLER_24_39 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_4.mux_l1_in_4__A1 top_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 top_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XFILLER_14_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A0 mux_left_track_5.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l3_in_0__A0 mux_left_track_15.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_233 vpwr vgnd scs8hd_fill_2
XFILLER_36_115 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 chany_bottom_in[18] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_3__S mux_left_track_5.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A1 mux_bottom_track_17.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l3_in_0__S mux_left_track_3.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_33.mux_l1_in_2__A0 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l4_in_0__A0 mux_bottom_track_9.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_4.mux_l1_in_5__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XFILLER_33_118 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_18_126 vgnd vpwr scs8hd_fill_1
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__S mux_left_track_9.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_2.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_0.mux_l4_in_0_/S mux_top_track_2.mux_l1_in_0_/S
+ mem_top_track_2.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_top_track_16.mux_l1_in_3__A0 _035_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l2_in_3__A1 mux_top_track_4.mux_l1_in_6_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_97 vgnd vpwr scs8hd_fill_1
XFILLER_2_20 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_ top_left_grid_pin_37_ top_left_grid_pin_35_ mux_top_track_2.mux_l1_in_0_/S
+ mux_top_track_2.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 chany_top_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_21_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D mux_left_track_5.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l3_in_0__A0 mux_left_track_5.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_3__S mux_top_track_8.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
X_051_ _051_/HI _051_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_23_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_2__A1 chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_2__D mux_top_track_24.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_81 vgnd vpwr scs8hd_decap_4
XFILLER_36_70 vpwr vgnd scs8hd_fill_2
XFILLER_14_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_33.mux_l2_in_1__A0 _045_/HI vgnd vpwr scs8hd_diode_2
XFILLER_37_243 vgnd vpwr scs8hd_fill_1
XFILLER_20_110 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S mem_bottom_track_25.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ chany_bottom_in[9] chany_top_out[10] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_left_track_13.scs8hd_dfxbp_1_2__D mux_left_track_13.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_0_/S mux_bottom_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_7_136 vgnd vpwr scs8hd_decap_4
XFILLER_11_176 vgnd vpwr scs8hd_decap_4
X_034_ _034_/HI _034_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A1 chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_243 vgnd vpwr scs8hd_fill_1
XFILLER_8_41 vgnd vpwr scs8hd_decap_3
XFILLER_27_39 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 mux_bottom_track_25.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_1__S mux_bottom_track_33.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_1.scs8hd_buf_4_0_ mux_left_track_1.mux_l3_in_0_/X _073_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_33.mux_l3_in_0__A0 mux_bottom_track_33.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l2_in_1__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_38_16 vpwr vgnd scs8hd_fill_2
XFILLER_38_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_19.scs8hd_buf_4_0__A mux_left_track_19.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_ bottom_left_grid_pin_35_ bottom_right_grid_pin_1_
+ mux_bottom_track_1.mux_l1_in_1_/S mux_bottom_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_205 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_1__A1 mux_bottom_track_9.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_left_track_23.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_21.mux_l2_in_0_/S mux_left_track_23.mux_l1_in_1_/S
+ mem_left_track_23.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_2__D mux_top_track_0.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_3.mux_l3_in_0_/S mux_left_track_5.mux_l1_in_3_/S
+ mem_left_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_20 vgnd vpwr scs8hd_decap_4
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_39_179 vpwr vgnd scs8hd_fill_2
XFILLER_39_146 vpwr vgnd scs8hd_fill_2
XFILLER_39_135 vgnd vpwr scs8hd_fill_1
XFILLER_39_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__D mux_left_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_1__A1 mux_left_track_5.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l3_in_0__A1 mux_left_track_15.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_40 vgnd vpwr scs8hd_fill_1
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_30_50 vgnd vpwr scs8hd_decap_4
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l1_in_3__A0 _037_/HI vgnd vpwr scs8hd_diode_2
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l4_in_0__A1 mux_bottom_track_9.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_2__A1 chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vpwr vgnd scs8hd_fill_2
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XFILLER_41_71 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.scs8hd_dfxbp_1_1__D mux_left_track_15.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_43 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_3__A1 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
XFILLER_17_160 vpwr vgnd scs8hd_fill_2
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_5.mux_l3_in_0__A1 mux_left_track_5.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_108 vpwr vgnd scs8hd_fill_2
X_050_ _050_/HI _050_/LO vgnd vpwr scs8hd_conb_1
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_11_30 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_33.mux_l2_in_1__A1 mux_bottom_track_33.mux_l1_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0__S mux_left_track_11.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_200 vgnd vpwr scs8hd_decap_12
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_25.mux_l1_in_2_/S
+ mux_bottom_track_25.mux_l2_in_1_/S mem_bottom_track_25.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_17.mux_l1_in_1__S mux_left_track_17.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
X_102_ chany_bottom_in[10] chany_top_out[11] vgnd vpwr scs8hd_buf_2
X_033_ _033_/HI _033_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_1__D mux_top_track_2.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D mux_top_track_32.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_2__A0 chanx_left_in[11] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l3_in_0__A1 mux_bottom_track_33.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_50 vpwr vgnd scs8hd_fill_2
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XFILLER_38_28 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_13_217 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_0_165 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.scs8hd_buf_4_0__A mux_left_track_3.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_23.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_0__D mux_left_track_15.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_210 vgnd vpwr scs8hd_fill_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_114 vpwr vgnd scs8hd_fill_2
XFILLER_39_169 vpwr vgnd scs8hd_fill_2
XFILLER_39_158 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_19.mux_l1_in_1__A0 _053_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_1__A0 mux_top_track_8.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l1_in_3__A1 chanx_left_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_35_161 vpwr vgnd scs8hd_fill_2
XFILLER_27_128 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.scs8hd_buf_4_0_ mux_left_track_11.mux_l3_in_0_/X _068_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_9.mux_l4_in_0__S mux_bottom_track_9.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_7 vgnd vpwr scs8hd_decap_4
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
XFILLER_18_106 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_19.mux_l2_in_0__A0 mux_left_track_19.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_41_83 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _112_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l4_in_0__A0 mux_top_track_8.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D mux_top_track_2.mux_l4_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_131 vpwr vgnd scs8hd_fill_2
XFILLER_2_88 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_3__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_3__D mux_bottom_track_1.mux_l3_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__D mux_left_track_9.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vgnd vpwr scs8hd_fill_1
XFILLER_36_50 vgnd vpwr scs8hd_decap_4
XFILLER_14_120 vgnd vpwr scs8hd_decap_3
XANTENNA__107__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_7.mux_l1_in_3__A0 _032_/HI vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_212 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_5.mux_l2_in_1__S mux_left_track_5.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_167 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_25.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_17.mux_l3_in_0_/S
+ mux_bottom_track_25.mux_l1_in_2_/S mem_bottom_track_25.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
X_101_ _101_/A chany_top_out[12] vgnd vpwr scs8hd_buf_2
XFILLER_11_101 vpwr vgnd scs8hd_fill_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_4.mux_l2_in_3__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
X_032_ _032_/HI _032_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_85 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l4_in_0__S mux_top_track_2.mux_l4_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_3_ _031_/HI left_top_grid_pin_48_ mux_left_track_5.mux_l1_in_3_/S
+ mux_left_track_5.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_76 vpwr vgnd scs8hd_fill_2
XFILLER_8_87 vgnd vpwr scs8hd_decap_3
XFILLER_40_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l3_in_1__S mux_top_track_8.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l3_in_0_ mux_left_track_13.mux_l2_in_1_/X mux_left_track_13.mux_l2_in_0_/X
+ mux_left_track_13.mux_l3_in_0_/S mux_left_track_13.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_2__A1 chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_52 vgnd vpwr scs8hd_decap_3
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_4
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XFILLER_13_229 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_3__D mux_top_track_4.mux_l3_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_19.mux_l1_in_1__A1 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_1_ _050_/HI left_top_grid_pin_44_ mux_left_track_13.mux_l2_in_1_/S
+ mux_left_track_13.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_8.mux_l3_in_1__A1 mux_top_track_8.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_170 vgnd vpwr scs8hd_decap_3
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ mux_left_track_5.mux_l3_in_0_/S mux_left_track_5.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_20 vgnd vpwr scs8hd_fill_1
XFILLER_30_63 vpwr vgnd scs8hd_fill_2
XFILLER_5_214 vpwr vgnd scs8hd_fill_2
XFILLER_5_225 vpwr vgnd scs8hd_fill_2
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_29_181 vpwr vgnd scs8hd_fill_2
XFILLER_27_118 vgnd vpwr scs8hd_decap_4
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_165 vpwr vgnd scs8hd_fill_2
XPHY_74 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_19.mux_l2_in_0__A1 mux_left_track_19.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XFILLER_25_85 vgnd vpwr scs8hd_decap_4
XFILLER_25_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_95 vgnd vpwr scs8hd_decap_12
XFILLER_41_62 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_8.mux_l4_in_0__A1 mux_top_track_8.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_121 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_24.scs8hd_buf_4_0__A mux_top_track_24.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_10 vgnd vpwr scs8hd_decap_4
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XFILLER_14_198 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l1_in_3__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_20_146 vgnd vpwr scs8hd_decap_4
XFILLER_28_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0__A1 mux_left_track_9.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
X_100_ chany_bottom_in[12] chany_top_out[13] vgnd vpwr scs8hd_buf_2
X_031_ _031_/HI _031_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_16.scs8hd_buf_4_0_ mux_top_track_16.mux_l3_in_0_/X _105_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l1_in_2_ left_top_grid_pin_46_ left_top_grid_pin_44_ mux_left_track_5.mux_l1_in_3_/S
+ mux_left_track_5.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 bottom_right_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_40_219 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A mux_bottom_track_1.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_6_/S
+ vgnd vpwr scs8hd_diode_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_42 vgnd vpwr scs8hd_decap_4
XFILLER_3_197 vpwr vgnd scs8hd_fill_2
XFILLER_3_153 vgnd vpwr scs8hd_fill_1
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_19.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_0_178 vpwr vgnd scs8hd_fill_2
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S mux_top_track_32.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_28_52 vpwr vgnd scs8hd_fill_2
XFILLER_28_41 vpwr vgnd scs8hd_fill_2
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_12 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_33.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_33.mux_l2_in_1_/S
+ mux_bottom_track_33.mux_l3_in_0_/S mem_bottom_track_33.scs8hd_dfxbp_1_2_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_39_127 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_3_ _040_/HI chanx_left_in[18] mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_13.mux_l2_in_0_ chany_bottom_in[15] mux_left_track_13.mux_l1_in_0_/X
+ mux_left_track_13.mux_l2_in_1_/S mux_left_track_13.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_left_track_13.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_13.mux_l2_in_1_/S mux_left_track_13.mux_l3_in_0_/S
+ mem_left_track_13.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_54 vpwr vgnd scs8hd_fill_2
XFILLER_5_237 vgnd vpwr scs8hd_decap_4
XFILLER_39_51 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
Xmux_top_track_32.mux_l2_in_1_ _038_/HI mux_top_track_32.mux_l1_in_2_/X mux_top_track_32.mux_l2_in_1_/S
+ mux_top_track_32.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_163 vgnd vpwr scs8hd_decap_12
XFILLER_26_152 vgnd vpwr scs8hd_fill_1
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_18_119 vgnd vpwr scs8hd_decap_4
XFILLER_41_41 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_24 vpwr vgnd scs8hd_fill_2
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_144 vpwr vgnd scs8hd_fill_2
XFILLER_17_174 vpwr vgnd scs8hd_fill_2
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D mux_top_track_8.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S mux_left_track_5.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_111 vpwr vgnd scs8hd_fill_2
XFILLER_23_166 vpwr vgnd scs8hd_fill_2
Xmux_top_track_24.scs8hd_buf_4_0_ mux_top_track_24.mux_l3_in_0_/X _101_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_bottom_track_5.mux_l4_in_0__S mux_bottom_track_5.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ mux_top_track_8.mux_l4_in_0_/S mux_top_track_8.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XFILLER_42_7 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l1_in_2_ chanx_left_in[15] chanx_left_in[8] mux_top_track_32.mux_l1_in_2_/S
+ mux_top_track_32.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_114 vpwr vgnd scs8hd_fill_2
XFILLER_20_125 vpwr vgnd scs8hd_fill_2
XFILLER_9_181 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
X_030_ _030_/HI _030_/LO vgnd vpwr scs8hd_conb_1
XFILLER_22_10 vpwr vgnd scs8hd_fill_2
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_34_206 vgnd vpwr scs8hd_decap_8
Xmux_left_track_5.mux_l1_in_1_ left_top_grid_pin_42_ chany_bottom_in[5] mux_left_track_5.mux_l1_in_3_/S
+ mux_left_track_5.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_19_203 vgnd vpwr scs8hd_decap_12
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XFILLER_6_162 vgnd vpwr scs8hd_decap_4
XFILLER_6_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_21.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_1.mux_l2_in_1__S mux_left_track_1.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_20 vgnd vpwr scs8hd_decap_3
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l2_in_3__S mux_top_track_0.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_2__S mux_left_track_7.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_3.scs8hd_buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X _092_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_21_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l3_in_1__S mux_top_track_4.mux_l3_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_28_97 vgnd vpwr scs8hd_fill_1
XFILLER_8_202 vpwr vgnd scs8hd_fill_2
XFILLER_8_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_24 vgnd vpwr scs8hd_fill_1
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_33.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l2_in_1_/S mem_bottom_track_33.scs8hd_dfxbp_1_1_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_39_106 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l2_in_2_ chanx_left_in[11] chanx_left_in[4] mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 mux_top_track_0.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_13.mux_l1_in_0_/S mux_left_track_13.mux_l2_in_1_/S
+ mem_left_track_13.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_2_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XFILLER_39_85 vpwr vgnd scs8hd_fill_2
XFILLER_29_161 vgnd vpwr scs8hd_decap_12
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_32.scs8hd_buf_4_0_ mux_top_track_32.mux_l3_in_0_/X _097_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_175 vgnd vpwr scs8hd_decap_12
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_53 vgnd vpwr scs8hd_decap_8
Xmux_left_track_13.mux_l1_in_0_ chany_bottom_in[10] chany_top_in[10] mux_left_track_13.mux_l1_in_0_/S
+ mux_left_track_13.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_36 vgnd vpwr scs8hd_fill_1
XFILLER_17_164 vpwr vgnd scs8hd_fill_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XFILLER_32_101 vgnd vpwr scs8hd_fill_1
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ ccff_tail mux_left_track_25.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_123 vpwr vgnd scs8hd_fill_2
XFILLER_11_78 vpwr vgnd scs8hd_fill_2
XFILLER_14_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_2__S mux_top_track_24.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_7 vgnd vpwr scs8hd_decap_3
XFILLER_28_6 vpwr vgnd scs8hd_fill_2
Xmux_top_track_32.mux_l1_in_1_ chanx_left_in[1] chany_bottom_in[10] mux_top_track_32.mux_l1_in_2_/S
+ mux_top_track_32.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_9_171 vgnd vpwr scs8hd_decap_4
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_16.mux_l2_in_0_/S mux_top_track_16.mux_l3_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_2__D mux_top_track_32.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_55 vpwr vgnd scs8hd_fill_2
XFILLER_11_148 vgnd vpwr scs8hd_decap_4
XFILLER_11_159 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_ chany_bottom_in[1] chany_top_in[5] mux_left_track_5.mux_l1_in_3_/S
+ mux_left_track_5.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_19_215 vgnd vpwr scs8hd_decap_12
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A mux_bottom_track_9.mux_l4_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_1_ _029_/HI left_top_grid_pin_42_ mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
X_089_ _089_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_10_192 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA__060__A left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XFILLER_17_11 vpwr vgnd scs8hd_fill_2
XFILLER_17_99 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 top_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_87 vpwr vgnd scs8hd_fill_2
XFILLER_33_54 vpwr vgnd scs8hd_fill_2
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_3_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_3__A0 _041_/HI vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.scs8hd_buf_4_0_ mux_left_track_7.mux_l3_in_0_/X _070_/A vgnd vpwr
+ scs8hd_buf_1
Xmem_top_track_0.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l4_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__055__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_21_232 vgnd vpwr scs8hd_decap_12
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_28_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_28_87 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_36 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_33.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_33.mux_l1_in_1_/S mem_bottom_track_33.scs8hd_dfxbp_1_0_/QN vgnd
+ vpwr scs8hd_dfxbp_1
XFILLER_39_118 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_1_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_0.scs8hd_buf_4_0_ mux_top_track_0.mux_l4_in_0_/X _113_/A vgnd vpwr
+ scs8hd_buf_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_11.mux_l3_in_0_/S mux_left_track_13.mux_l1_in_0_/S
+ mem_left_track_13.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_33.mux_l3_in_0__S mux_bottom_track_33.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_11 vpwr vgnd scs8hd_fill_2
XFILLER_14_12 vpwr vgnd scs8hd_fill_2
XFILLER_14_23 vpwr vgnd scs8hd_fill_2
XFILLER_14_67 vpwr vgnd scs8hd_fill_2
XFILLER_39_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_25.mux_l2_in_0__S ccff_tail vgnd vpwr scs8hd_diode_2
XFILLER_30_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_39_97 vgnd vpwr scs8hd_fill_1
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_173 vgnd vpwr scs8hd_decap_8
XFILLER_35_165 vgnd vpwr scs8hd_decap_12
XFILLER_35_132 vpwr vgnd scs8hd_fill_2
XFILLER_2_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_19.mux_l1_in_0__S mux_left_track_19.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_187 vgnd vpwr scs8hd_decap_12
XFILLER_25_11 vgnd vpwr scs8hd_fill_1
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_1_253 vgnd vpwr scs8hd_decap_12
XFILLER_1_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_143 vpwr vgnd scs8hd_fill_2
XFILLER_23_135 vpwr vgnd scs8hd_fill_2
XFILLER_23_102 vgnd vpwr scs8hd_decap_3
XANTENNA__063__A _063_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_87 vgnd vpwr scs8hd_decap_4
XFILLER_36_54 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_23.scs8hd_dfxbp_1_1__D mux_left_track_23.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_32.mux_l1_in_0_ top_left_grid_pin_41_ top_left_grid_pin_37_ mux_top_track_32.mux_l1_in_2_/S
+ mux_top_track_32.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_16.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_16.mux_l1_in_0_/S mux_top_track_16.mux_l2_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XANTENNA__058__A chany_top_in[15] vgnd vpwr scs8hd_diode_2
XFILLER_22_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_11_105 vgnd vpwr scs8hd_decap_4
XFILLER_22_89 vgnd vpwr scs8hd_fill_1
XFILLER_22_78 vgnd vpwr scs8hd_decap_4
XFILLER_19_227 vgnd vpwr scs8hd_decap_12
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.scs8hd_buf_4_0__A mux_top_track_4.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l2_in_3__S mux_bottom_track_3.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_25.mux_l1_in_0_ chany_bottom_in[18] chany_top_in[18] mux_left_track_25.mux_l1_in_0_/S
+ mux_left_track_25.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_10_160 vpwr vgnd scs8hd_fill_2
XFILLER_10_171 vpwr vgnd scs8hd_fill_2
XFILLER_40_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l4_in_0__S mux_bottom_track_1.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
X_088_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_15.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_89 vgnd vpwr scs8hd_decap_4
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_44 vgnd vpwr scs8hd_decap_4
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_156 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_3__A1 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.scs8hd_buf_4_0__A mux_top_track_32.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_241 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_0.mux_l2_in_1_/S mux_top_track_0.mux_l3_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_top_track_16.scs8hd_dfxbp_1_0__D mux_top_track_8.mux_l4_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA__071__A _071_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_200 vgnd vpwr scs8hd_decap_12
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_2_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_ top_right_grid_pin_1_ mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_2__S mux_left_track_3.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__066__A _066_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XFILLER_5_229 vpwr vgnd scs8hd_fill_2
XFILLER_30_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D mux_left_track_23.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l3_in_1__S mux_top_track_0.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0__S mux_left_track_7.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_177 vgnd vpwr scs8hd_decap_6
XFILLER_35_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 top_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_6_80 vgnd vpwr scs8hd_fill_1
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_169 vgnd vpwr scs8hd_decap_12
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XFILLER_41_11 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_199 vgnd vpwr scs8hd_decap_12
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_1_210 vpwr vgnd scs8hd_fill_2
XFILLER_2_16 vpwr vgnd scs8hd_fill_2
XFILLER_1_265 vgnd vpwr scs8hd_decap_12
XFILLER_1_243 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.scs8hd_buf_4_0_ mux_left_track_17.mux_l2_in_0_/X _065_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_32_125 vgnd vpwr scs8hd_decap_4
XFILLER_23_158 vpwr vgnd scs8hd_fill_2
XFILLER_11_14 vgnd vpwr scs8hd_fill_1
XFILLER_36_99 vgnd vpwr scs8hd_fill_1
XFILLER_36_77 vpwr vgnd scs8hd_fill_2
XFILLER_36_66 vpwr vgnd scs8hd_fill_2
XFILLER_36_22 vgnd vpwr scs8hd_decap_3
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
XFILLER_14_136 vpwr vgnd scs8hd_fill_2
XFILLER_14_158 vpwr vgnd scs8hd_fill_2
Xmem_left_track_3.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_3.mux_l2_in_1_/S mux_left_track_3.mux_l3_in_0_/S
+ mem_left_track_3.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_37_217 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_8.mux_l4_in_0_/S mux_top_track_16.mux_l1_in_0_/S
+ mem_top_track_16.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_20_106 vpwr vgnd scs8hd_fill_2
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.scs8hd_dfxbp_1_3_ prog_clk mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l4_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA__074__A chany_top_in[18] vgnd vpwr scs8hd_diode_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_239 vgnd vpwr scs8hd_decap_4
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_087_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_154 vpwr vgnd scs8hd_fill_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _069_/A vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_12 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_8.scs8hd_dfxbp_1_3_ prog_clk mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l4_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_3_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_3_102 vgnd vpwr scs8hd_fill_1
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_0.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_0.mux_l1_in_0_/S mux_top_track_0.mux_l2_in_1_/S
+ mem_top_track_0.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_9_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_3__A0 _034_/HI vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_32.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_138 vgnd vpwr scs8hd_decap_3
XFILLER_28_56 vpwr vgnd scs8hd_fill_2
XFILLER_28_45 vpwr vgnd scs8hd_fill_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l1_in_0__A0 chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_12_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_5_16 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_142 vpwr vgnd scs8hd_fill_2
XFILLER_38_120 vgnd vpwr scs8hd_decap_4
XFILLER_14_36 vpwr vgnd scs8hd_fill_2
XFILLER_30_46 vpwr vgnd scs8hd_fill_2
XANTENNA__082__A chany_top_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_39_55 vpwr vgnd scs8hd_fill_2
Xmux_left_track_25.scs8hd_buf_4_0_ mux_left_track_25.mux_l2_in_0_/X _061_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_2__A0 mux_bottom_track_5.mux_l1_in_5_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_26_134 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vpwr vgnd scs8hd_fill_2
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_25_46 vpwr vgnd scs8hd_fill_2
XFILLER_1_222 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l1_in_0_ top_left_grid_pin_38_ top_left_grid_pin_34_ mux_top_track_8.mux_l1_in_0_/S
+ mux_top_track_8.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_2_39 vpwr vgnd scs8hd_fill_2
XFILLER_2_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_32_148 vgnd vpwr scs8hd_decap_4
XFILLER_17_123 vgnd vpwr scs8hd_fill_1
XFILLER_17_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_21.mux_l2_in_0__S mux_left_track_21.mux_l2_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_31_181 vpwr vgnd scs8hd_fill_2
XFILLER_23_115 vgnd vpwr scs8hd_decap_4
XFILLER_11_26 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 left_top_grid_pin_46_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_1__A0 _049_/HI vgnd vpwr scs8hd_diode_2
XFILLER_14_148 vgnd vpwr scs8hd_decap_3
Xmem_left_track_21.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_21.mux_l1_in_0_/S mux_left_track_21.mux_l2_in_0_/S
+ mem_left_track_21.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_left_track_3.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_3.mux_l1_in_1_/S mux_left_track_3.mux_l2_in_1_/S
+ mem_left_track_3.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_15.mux_l1_in_0__S mux_left_track_15.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_1__A0 mux_bottom_track_5.mux_l2_in_3_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_129 vpwr vgnd scs8hd_fill_2
XFILLER_3_71 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.scs8hd_dfxbp_1_2_ prog_clk mux_bottom_track_5.mux_l2_in_3_/S mux_bottom_track_5.mux_l3_in_0_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l3_in_0__S mux_top_track_16.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
X_086_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_33_7 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_1__A0 mux_left_track_1.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l3_in_0__A0 mux_left_track_11.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l3_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _085_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l4_in_0__A0 mux_bottom_track_5.mux_l3_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.scs8hd_dfxbp_1_0_ prog_clk ccff_head mux_top_track_0.mux_l1_in_0_/S
+ mem_top_track_0.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
X_069_ _069_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l2_in_3__A1 chanx_left_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_28_79 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l1_in_0__A1 chany_top_in[10] vgnd vpwr scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l3_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_8_206 vgnd vpwr scs8hd_decap_4
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l3_in_0__A0 mux_left_track_1.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_3__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_4__S mux_bottom_track_5.mux_l1_in_6_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_1__S mux_bottom_track_3.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_6_ chanx_left_in[19] chanx_left_in[12] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_6_/X vgnd vpwr scs8hd_mux2_1
XFILLER_30_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l2_in_2__S mux_bottom_track_9.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_89 vgnd vpwr scs8hd_decap_8
XFILLER_29_132 vpwr vgnd scs8hd_fill_2
XFILLER_29_110 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l3_in_0__S mux_left_track_13.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_3__S mux_bottom_track_17.mux_l1_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_2__A1 mux_bottom_track_5.mux_l1_in_4_/X vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_146 vgnd vpwr scs8hd_decap_6
XFILLER_26_113 vpwr vgnd scs8hd_fill_2
XFILLER_25_14 vpwr vgnd scs8hd_fill_2
XPHY_47 vgnd vpwr scs8hd_decap_3
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_41_68 vgnd vpwr scs8hd_fill_1
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_171 vgnd vpwr scs8hd_decap_8
XFILLER_15_91 vpwr vgnd scs8hd_fill_2
XFILLER_17_168 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_3_ _048_/HI left_top_grid_pin_48_ mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_23_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0__S mux_left_track_3.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.scs8hd_buf_4_0__A mux_left_track_17.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 left_top_grid_pin_44_ vgnd vpwr scs8hd_diode_2
XFILLER_36_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l2_in_1__A1 left_top_grid_pin_43_ vgnd vpwr scs8hd_diode_2
XANTENNA__088__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_116 vpwr vgnd scs8hd_fill_2
Xmem_left_track_3.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_1.mux_l3_in_0_/S mux_left_track_3.mux_l1_in_1_/S
+ mem_left_track_3.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
Xmem_left_track_21.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_19.mux_l2_in_0_/S mux_left_track_21.mux_l1_in_0_/S
+ mem_left_track_21.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_13.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_2__S mux_top_track_2.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_1__A1 mux_bottom_track_5.mux_l2_in_2_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.scs8hd_dfxbp_1_1_ prog_clk mux_bottom_track_5.mux_l1_in_6_/S mux_bottom_track_5.mux_l2_in_3_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_10_141 vpwr vgnd scs8hd_fill_2
X_085_ _085_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 bottom_left_grid_pin_38_ vgnd vpwr scs8hd_diode_2
XFILLER_6_112 vpwr vgnd scs8hd_fill_2
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_6_189 vgnd vpwr scs8hd_decap_4
XFILLER_10_196 vgnd vpwr scs8hd_decap_4
XFILLER_26_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_1__A1 mux_left_track_1.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l3_in_0__A1 mux_left_track_11.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_21.mux_l1_in_0__A1 chany_top_in[16] vgnd vpwr scs8hd_diode_2
XFILLER_24_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_17_15 vpwr vgnd scs8hd_fill_2
XFILLER_17_48 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_8.mux_l1_in_0_/S mux_top_track_8.mux_l2_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ mux_left_track_1.mux_l3_in_0_/S mux_left_track_1.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_58 vgnd vpwr scs8hd_decap_3
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_5.mux_l4_in_0__A1 mux_bottom_track_5.mux_l3_in_0_/X vgnd
+ vpwr scs8hd_diode_2
X_068_ _068_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_192 vpwr vgnd scs8hd_fill_2
XFILLER_0_51 vpwr vgnd scs8hd_fill_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_71 vgnd vpwr scs8hd_decap_4
XFILLER_0_107 vgnd vpwr scs8hd_decap_3
XANTENNA__096__A chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_1.mux_l3_in_0__A1 mux_left_track_1.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_1__S mux_top_track_32.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_9.scs8hd_buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X _089_/A vgnd
+ vpwr scs8hd_buf_1
Xmux_top_track_4.mux_l1_in_5_ chanx_left_in[5] chany_bottom_in[14] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_5_/X vgnd vpwr scs8hd_mux2_1
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_38_188 vgnd vpwr scs8hd_decap_12
XFILLER_38_177 vgnd vpwr scs8hd_decap_8
XFILLER_14_16 vgnd vpwr scs8hd_decap_4
XFILLER_14_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_3__A0 top_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
XFILLER_39_24 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_136 vgnd vpwr scs8hd_decap_4
XFILLER_35_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_72 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_37 vpwr vgnd scs8hd_fill_2
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XFILLER_41_25 vpwr vgnd scs8hd_fill_2
XFILLER_1_235 vgnd vpwr scs8hd_decap_8
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_147 vpwr vgnd scs8hd_fill_2
XFILLER_40_183 vgnd vpwr scs8hd_decap_8
XFILLER_25_180 vgnd vpwr scs8hd_decap_3
Xmux_left_track_1.mux_l1_in_2_ left_top_grid_pin_46_ left_top_grid_pin_44_ mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_31_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l2_in_2__A0 mux_top_track_4.mux_l1_in_5_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_161 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.scs8hd_buf_4_0__A mux_left_track_1.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 bottom_left_grid_pin_39_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_132 vpwr vgnd scs8hd_fill_2
XFILLER_9_154 vpwr vgnd scs8hd_fill_2
XFILLER_13_161 vgnd vpwr scs8hd_fill_1
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
Xmem_bottom_track_5.scs8hd_dfxbp_1_0_ prog_clk mux_bottom_track_3.mux_l4_in_0_/S mux_bottom_track_5.mux_l1_in_6_/S
+ mem_bottom_track_5.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D mux_left_track_1.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_27 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A chany_bottom_in[13] vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l3_in_1__A0 mux_top_track_4.mux_l2_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_131 vgnd vpwr scs8hd_fill_1
XFILLER_10_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_23.mux_l1_in_1__S mux_left_track_23.mux_l1_in_1_/S vgnd vpwr
+ scs8hd_diode_2
X_084_ chany_top_in[8] chany_bottom_out[9] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 bottom_left_grid_pin_34_ vgnd vpwr scs8hd_diode_2
XFILLER_6_168 vpwr vgnd scs8hd_fill_2
XFILLER_12_60 vpwr vgnd scs8hd_fill_2
XFILLER_19_7 vgnd vpwr scs8hd_fill_1
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0__S mux_left_track_11.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 bottom_left_grid_pin_41_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_3_ _039_/HI mux_top_track_4.mux_l1_in_6_/X mux_top_track_4.mux_l2_in_1_/S
+ mux_top_track_4.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 mux_bottom_track_25.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__S mux_bottom_track_25.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_track_8.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_4.mux_l4_in_0_/S mux_top_track_8.mux_l1_in_0_/S
+ mem_top_track_8.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_17_38 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_149 vgnd vpwr scs8hd_decap_4
XFILLER_3_105 vpwr vgnd scs8hd_fill_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_6__A0 chanx_left_in[17] vgnd vpwr scs8hd_diode_2
X_067_ _067_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 left_top_grid_pin_42_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l2_in_0__A0 chany_bottom_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l4_in_0__A0 mux_top_track_4.mux_l3_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_24.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_16.mux_l3_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ mem_top_track_24.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l1_in_4_ chany_bottom_in[5] top_right_grid_pin_1_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_4_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_0_/S mux_left_track_1.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_3__A1 top_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_3__A0 _030_/HI vgnd vpwr scs8hd_diode_2
XFILLER_30_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ mux_top_track_4.mux_l4_in_0_/S mux_top_track_4.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l2_in_0__A0 mux_left_track_5.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_104 vgnd vpwr scs8hd_fill_1
XFILLER_6_51 vpwr vgnd scs8hd_fill_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_41_107 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.scs8hd_dfxbp_1_0__D mux_left_track_1.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_170 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A0 chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_1_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_2__S mux_bottom_track_5.mux_l2_in_3_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_195 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_1_ left_top_grid_pin_42_ chany_bottom_in[2] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_2__A1 mux_top_track_4.mux_l1_in_4_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2__A0 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XFILLER_23_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_23.mux_l1_in_1__A0 _028_/HI vgnd vpwr scs8hd_diode_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_173 vgnd vpwr scs8hd_decap_8
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_1_/S mux_top_track_4.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A1 bottom_left_grid_pin_35_ vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_1__S mux_left_track_15.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_11.scs8hd_dfxbp_1_1__D mux_left_track_11.mux_l1_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 mux_bottom_track_33.mux_l1_in_1_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_177 vpwr vgnd scs8hd_fill_2
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l2_in_1__S mux_bottom_track_17.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l3_in_1__A1 mux_top_track_4.mux_l2_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A0 mux_top_track_16.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
X_083_ chany_top_in[9] chany_bottom_out[10] vgnd vpwr scs8hd_buf_2
XFILLER_10_154 vgnd vpwr scs8hd_decap_4
XFILLER_12_72 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_23.mux_l2_in_0__A0 mux_left_track_23.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_210 vgnd vpwr scs8hd_decap_4
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 bottom_left_grid_pin_37_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_2_ mux_top_track_4.mux_l1_in_5_/X mux_top_track_4.mux_l1_in_4_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_5.mux_l1_in_1__S mux_left_track_5.mux_l1_in_3_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_16 vpwr vgnd scs8hd_fill_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_4.mux_l1_in_3__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_30_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_6__A1 chanx_left_in[10] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
X_066_ _066_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_7 vpwr vgnd scs8hd_fill_2
XFILLER_24_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l2_in_0__A1 mux_left_track_15.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_4.mux_l4_in_0__A1 mux_top_track_4.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l3_in_0__A0 mux_top_track_16.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_19.mux_l2_in_0_ mux_left_track_19.mux_l1_in_1_/X mux_left_track_19.mux_l1_in_0_/X
+ mux_left_track_19.mux_l2_in_0_/S mux_left_track_19.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D mux_top_track_16.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_82 vgnd vpwr scs8hd_decap_4
Xmux_top_track_4.mux_l1_in_3_ top_left_grid_pin_41_ top_left_grid_pin_40_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_7_220 vpwr vgnd scs8hd_fill_2
X_049_ _049_/HI _049_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_146 vgnd vpwr scs8hd_decap_6
Xmux_left_track_21.mux_l2_in_0_ mux_left_track_21.mux_l1_in_1_/X mux_left_track_21.mux_l1_in_0_/X
+ mux_left_track_21.mux_l2_in_0_/S mux_left_track_21.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_3__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
XFILLER_39_59 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_2__D mux_bottom_track_17.mux_l2_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0__A1 mux_left_track_5.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_13.scs8hd_dfxbp_1_0__D mux_left_track_11.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_4_223 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l1_in_2__A0 chanx_left_in[9] vgnd vpwr scs8hd_diode_2
XFILLER_20_72 vgnd vpwr scs8hd_decap_3
XFILLER_28_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_11.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_26_105 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A1 bottom_left_grid_pin_40_ vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_119 vgnd vpwr scs8hd_decap_3
XFILLER_34_182 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_3_ _044_/HI chanx_left_in[16] mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l2_in_3_/X vgnd vpwr scs8hd_mux2_1
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_left_track_19.mux_l1_in_1_ _053_/HI left_top_grid_pin_47_ mux_left_track_19.mux_l1_in_0_/S
+ mux_left_track_19.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_25_160 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_ chany_top_in[2] chany_top_in[0] mux_left_track_1.mux_l1_in_0_/S
+ mux_left_track_1.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
Xmem_top_track_32.scs8hd_dfxbp_1_2_ prog_clk mux_top_track_32.mux_l2_in_1_/S mux_top_track_32.mux_l3_in_0_/S
+ mem_top_track_32.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
Xmux_left_track_21.mux_l1_in_1_ _027_/HI left_top_grid_pin_48_ mux_left_track_21.mux_l1_in_0_/S
+ mux_left_track_21.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_2__A1 chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.scs8hd_buf_4_0__A mux_left_track_9.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_23_119 vgnd vpwr scs8hd_fill_1
XFILLER_16_171 vpwr vgnd scs8hd_fill_2
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_23.mux_l1_in_1__A1 left_top_grid_pin_49_ vgnd vpwr scs8hd_diode_2
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_1_/S mux_top_track_4.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_36_27 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_24.mux_l2_in_1__A0 mux_top_track_24.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_4.mux_l1_in_6__S mux_top_track_4.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
XFILLER_26_93 vgnd vpwr scs8hd_decap_3
XFILLER_13_174 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D ccff_head vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_145 vpwr vgnd scs8hd_fill_2
XFILLER_9_167 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.scs8hd_dfxbp_1_2_ prog_clk mux_left_track_11.mux_l2_in_1_/S mux_left_track_11.mux_l3_in_0_/S
+ mem_left_track_11.scs8hd_dfxbp_1_2_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mem_left_track_5.scs8hd_dfxbp_1_2__D mux_left_track_5.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A1 mux_top_track_16.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
X_082_ chany_top_in[10] chany_bottom_out[11] vgnd vpwr scs8hd_buf_2
XFILLER_10_111 vpwr vgnd scs8hd_fill_2
XFILLER_10_188 vpwr vgnd scs8hd_fill_2
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_23.mux_l2_in_0__A1 mux_left_track_23.mux_l1_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_92 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ mux_bottom_track_3.mux_l4_in_0_/S mux_bottom_track_3.mux_l4_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_24.mux_l3_in_0__A0 mux_top_track_24.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 chany_bottom_in[16] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_25.scs8hd_buf_4_0__A mux_left_track_25.mux_l2_in_0_/X vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
X_065_ _065_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_2_162 vgnd vpwr scs8hd_decap_4
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_9_41 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_33.mux_l1_in_2__S mux_bottom_track_33.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l3_in_0__A1 mux_top_track_16.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_6__A0 chanx_left_in[19] vgnd vpwr scs8hd_diode_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_32.mux_l1_in_2__A0 chanx_left_in[15] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_1_/X vgnd vpwr scs8hd_mux2_1
Xmux_top_track_4.mux_l1_in_2_ top_left_grid_pin_39_ top_left_grid_pin_38_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_34_82 vgnd vpwr scs8hd_decap_3
XFILLER_7_243 vgnd vpwr scs8hd_fill_1
X_048_ _048_/HI _048_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_158 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 chany_bottom_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_136 vpwr vgnd scs8hd_fill_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_37_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_3_ _042_/HI chanx_left_in[19] mux_bottom_track_17.mux_l1_in_3_/S
+ mux_bottom_track_17.mux_l1_in_3_/X vgnd vpwr scs8hd_mux2_1
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_24.mux_l1_in_2__A1 chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_62 vgnd vpwr scs8hd_decap_4
XFILLER_20_84 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.scs8hd_dfxbp_1_3__D mux_top_track_0.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_7.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l2_in_1__A0 _038_/HI vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
Xmux_left_track_19.mux_l1_in_0_ chany_bottom_in[14] chany_top_in[14] mux_left_track_19.mux_l1_in_0_/S
+ mux_left_track_19.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_194 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_3.mux_l2_in_2_ chanx_left_in[9] chanx_left_in[2] mux_bottom_track_3.mux_l2_in_0_/S
+ mux_bottom_track_3.mux_l2_in_2_/X vgnd vpwr scs8hd_mux2_1
XFILLER_1_249 vpwr vgnd scs8hd_fill_2
XFILLER_1_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_7.scs8hd_dfxbp_1_1__D mux_left_track_7.mux_l1_in_2_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_15_95 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A chany_bottom_in[10] vgnd vpwr scs8hd_diode_2
Xmux_left_track_21.mux_l1_in_0_ chany_bottom_in[16] chany_top_in[16] mux_left_track_21.mux_l1_in_0_/S
+ mux_left_track_21.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_0_/S vgnd vpwr scs8hd_diode_2
Xmem_top_track_32.scs8hd_dfxbp_1_1_ prog_clk mux_top_track_32.mux_l1_in_2_/S mux_top_track_32.mux_l2_in_1_/S
+ mem_top_track_32.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_39_253 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_24.mux_l2_in_1__A1 mux_top_track_24.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_22_175 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_32.mux_l3_in_0__A0 mux_top_track_32.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_83 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_15.scs8hd_dfxbp_1_2__D mux_left_track_15.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_13_164 vgnd vpwr scs8hd_fill_1
XFILLER_13_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l1_in_2__A0 left_top_grid_pin_47_ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_2__S mux_bottom_track_1.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_3_98 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S mux_bottom_track_17.mux_l3_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
Xmem_left_track_11.scs8hd_dfxbp_1_1_ prog_clk mux_left_track_11.mux_l1_in_0_/S mux_left_track_11.mux_l2_in_1_/S
+ mem_left_track_11.scs8hd_dfxbp_1_1_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_2__CLK prog_clk vgnd vpwr scs8hd_diode_2
X_081_ _081_/A chany_bottom_out[12] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_116 vpwr vgnd scs8hd_fill_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_37_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 chany_top_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_24.mux_l3_in_0__A1 mux_top_track_24.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_left_track_11.mux_l2_in_1__S mux_left_track_11.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_160 vgnd vpwr scs8hd_decap_4
XFILLER_5_193 vpwr vgnd scs8hd_fill_2
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_1__A0 mux_left_track_7.mux_l1_in_3_/X vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
X_064_ _064_/A chanx_left_out[9] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_17.mux_l2_in_1_ mux_bottom_track_17.mux_l1_in_3_/X mux_bottom_track_17.mux_l1_in_2_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mem_top_track_2.scs8hd_dfxbp_1_2__D mux_top_track_2.mux_l2_in_1_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XANTENNA__110__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_0_55 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_1_/S
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_4.mux_l1_in_6__A1 chanx_left_in[12] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__S mux_left_track_1.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_32.mux_l1_in_2__A1 chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D mux_left_track_7.mux_l3_in_0_/S vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_40 vpwr vgnd scs8hd_fill_2
Xmux_top_track_4.mux_l1_in_1_ top_left_grid_pin_37_ top_left_grid_pin_36_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_1_/X vgnd vpwr scs8hd_mux2_1
XFILLER_34_61 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_233 vpwr vgnd scs8hd_fill_2
X_047_ _047_/HI _047_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A1 chany_top_in[14] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l3_in_0__A0 mux_left_track_7.mux_l2_in_1_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_39_28 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_2_ chanx_left_in[12] chanx_left_in[5] mux_bottom_track_17.mux_l1_in_3_/S
+ mux_bottom_track_17.mux_l1_in_2_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_1_/S vgnd vpwr scs8hd_diode_2
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_29_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.scs8hd_dfxbp_1_1__D mux_left_track_17.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_6_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l2_in_1__A1 mux_top_track_32.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_3.mux_l2_in_1_ bottom_left_grid_pin_40_ bottom_left_grid_pin_38_
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_1_/X vgnd vpwr scs8hd_mux2_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_41_29 vgnd vpwr scs8hd_decap_12
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_84 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vpwr vgnd scs8hd_fill_2
Xmem_top_track_32.scs8hd_dfxbp_1_0_ prog_clk mux_top_track_24.mux_l3_in_0_/S mux_top_track_32.mux_l1_in_2_/S
+ mem_top_track_32.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_184 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_3.scs8hd_buf_4_0_ mux_left_track_3.mux_l3_in_0_/X _072_/A vgnd vpwr
+ scs8hd_buf_1
XFILLER_39_265 vgnd vpwr scs8hd_decap_12
XFILLER_22_187 vgnd vpwr scs8hd_decap_12
XFILLER_26_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_32.mux_l3_in_0__A1 mux_top_track_32.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l1_in_2__A1 left_top_grid_pin_45_ vgnd vpwr scs8hd_diode_2
XFILLER_3_22 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D mux_top_track_4.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_213 vgnd vpwr scs8hd_fill_1
Xmem_left_track_11.scs8hd_dfxbp_1_0_ prog_clk mux_left_track_9.mux_l3_in_0_/S mux_left_track_11.mux_l1_in_0_/S
+ mem_left_track_11.scs8hd_dfxbp_1_0_/QN vgnd vpwr scs8hd_dfxbp_1
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D mux_bottom_track_1.mux_l4_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ chany_top_in[12] chany_bottom_out[13] vgnd vpwr scs8hd_buf_2
XFILLER_10_102 vgnd vpwr scs8hd_decap_3
XFILLER_10_124 vgnd vpwr scs8hd_decap_4
XFILLER_6_139 vgnd vpwr scs8hd_decap_4
XFILLER_12_64 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chany_top_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.scs8hd_buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X _085_/A vgnd
+ vpwr scs8hd_buf_1
XFILLER_38_3 vpwr vgnd scs8hd_fill_2
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XFILLER_3_109 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_7.mux_l2_in_1__A1 mux_left_track_7.mux_l1_in_2_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_15_205 vgnd vpwr scs8hd_decap_12
X_063_ _063_/A chanx_left_out[10] vgnd vpwr scs8hd_buf_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_0_/S mux_bottom_track_17.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_left_track_9.mux_l3_in_0__S mux_left_track_9.mux_l3_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__D mux_left_track_17.mux_l2_in_0_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_208 vgnd vpwr scs8hd_decap_12
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_20_263 vgnd vpwr scs8hd_decap_12
Xmux_top_track_4.mux_l1_in_0_ top_left_grid_pin_35_ top_left_grid_pin_34_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X vgnd vpwr scs8hd_mux2_1
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_19.scs8hd_dfxbp_1_0__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_11_241 vgnd vpwr scs8hd_decap_3
X_046_ _046_/HI _046_/LO vgnd vpwr scs8hd_conb_1
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_38_127 vgnd vpwr scs8hd_decap_8
XFILLER_22_6 vpwr vgnd scs8hd_fill_2
XFILLER_38_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l3_in_0__A1 mux_left_track_7.mux_l2_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_149 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_1_ bottom_left_grid_pin_38_ bottom_left_grid_pin_34_
+ mux_bottom_track_17.mux_l1_in_3_/S mux_bottom_track_17.mux_l1_in_1_/X vgnd vpwr
+ scs8hd_mux2_1
XANTENNA_mux_top_track_2.scs8hd_buf_4_0__A mux_top_track_2.mux_l4_in_0_/X vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_1_/S vgnd
+ vpwr scs8hd_diode_2
X_029_ _029_/HI _029_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_22 vgnd vpwr scs8hd_decap_4
XFILLER_6_55 vpwr vgnd scs8hd_fill_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XFILLER_34_152 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_0_/S mux_bottom_track_3.mux_l2_in_0_/X vgnd vpwr scs8hd_mux2_1
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S mux_bottom_track_33.mux_l2_in_1_/S vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__D mux_bottom_track_3.mux_l3_in_0_/S
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_166 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_25.mux_l1_in_0__S mux_left_track_25.mux_l1_in_0_/S vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_3__CLK prog_clk vgnd vpwr scs8hd_diode_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_16_141 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK prog_clk vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

