

module fpga_core
( prog_clk, Test_en, IO_ISOL_N, clk, gfpga_pad_EMBEDDED_IO_HD_SOC_IN, gfpga_pad_EMBEDDED_IO_HD_SOC_OUT, gfpga_pad_EMBEDDED_IO_HD_SOC_DIR, ccff_head, ccff_tail, sc_head, sc_tail ); 
  input [0:0] prog_clk;
  input [0:0] Test_en;
  input [0:0] IO_ISOL_N;
  input [0:0] clk;
  input [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;
  output [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
  output [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;
  input [0:0] ccff_head;
  output [0:0] ccff_tail;
  input sc_head;
  output sc_tail;

  wire [0:0] cbx_1__0__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__0_ccff_tail;
  wire [0:19] cbx_1__0__0_chanx_left_out;
  wire [0:19] cbx_1__0__0_chanx_right_out;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__1_ccff_tail;
  wire [0:19] cbx_1__0__1_chanx_left_out;
  wire [0:19] cbx_1__0__1_chanx_right_out;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__2_ccff_tail;
  wire [0:19] cbx_1__0__2_chanx_left_out;
  wire [0:19] cbx_1__0__2_chanx_right_out;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__3_ccff_tail;
  wire [0:19] cbx_1__0__3_chanx_left_out;
  wire [0:19] cbx_1__0__3_chanx_right_out;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__4_ccff_tail;
  wire [0:19] cbx_1__0__4_chanx_left_out;
  wire [0:19] cbx_1__0__4_chanx_right_out;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__5_ccff_tail;
  wire [0:19] cbx_1__0__5_chanx_left_out;
  wire [0:19] cbx_1__0__5_chanx_right_out;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__6_ccff_tail;
  wire [0:19] cbx_1__0__6_chanx_left_out;
  wire [0:19] cbx_1__0__6_chanx_right_out;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_16_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__0__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__0__7_ccff_tail;
  wire [0:19] cbx_1__0__7_chanx_left_out;
  wire [0:19] cbx_1__0__7_chanx_right_out;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__0_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__0_ccff_tail;
  wire [0:19] cbx_1__1__0_chanx_left_out;
  wire [0:19] cbx_1__1__0_chanx_right_out;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__10_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__10_ccff_tail;
  wire [0:19] cbx_1__1__10_chanx_left_out;
  wire [0:19] cbx_1__1__10_chanx_right_out;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__11_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__11_ccff_tail;
  wire [0:19] cbx_1__1__11_chanx_left_out;
  wire [0:19] cbx_1__1__11_chanx_right_out;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__12_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__12_ccff_tail;
  wire [0:19] cbx_1__1__12_chanx_left_out;
  wire [0:19] cbx_1__1__12_chanx_right_out;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__13_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__13_ccff_tail;
  wire [0:19] cbx_1__1__13_chanx_left_out;
  wire [0:19] cbx_1__1__13_chanx_right_out;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__14_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__14_ccff_tail;
  wire [0:19] cbx_1__1__14_chanx_left_out;
  wire [0:19] cbx_1__1__14_chanx_right_out;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__15_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__15_ccff_tail;
  wire [0:19] cbx_1__1__15_chanx_left_out;
  wire [0:19] cbx_1__1__15_chanx_right_out;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__16_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__16_ccff_tail;
  wire [0:19] cbx_1__1__16_chanx_left_out;
  wire [0:19] cbx_1__1__16_chanx_right_out;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__17_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__17_ccff_tail;
  wire [0:19] cbx_1__1__17_chanx_left_out;
  wire [0:19] cbx_1__1__17_chanx_right_out;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__18_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__18_ccff_tail;
  wire [0:19] cbx_1__1__18_chanx_left_out;
  wire [0:19] cbx_1__1__18_chanx_right_out;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__19_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__19_ccff_tail;
  wire [0:19] cbx_1__1__19_chanx_left_out;
  wire [0:19] cbx_1__1__19_chanx_right_out;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__1_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__1_ccff_tail;
  wire [0:19] cbx_1__1__1_chanx_left_out;
  wire [0:19] cbx_1__1__1_chanx_right_out;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__20_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__20_ccff_tail;
  wire [0:19] cbx_1__1__20_chanx_left_out;
  wire [0:19] cbx_1__1__20_chanx_right_out;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__21_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__21_ccff_tail;
  wire [0:19] cbx_1__1__21_chanx_left_out;
  wire [0:19] cbx_1__1__21_chanx_right_out;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__22_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__22_ccff_tail;
  wire [0:19] cbx_1__1__22_chanx_left_out;
  wire [0:19] cbx_1__1__22_chanx_right_out;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__23_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__23_ccff_tail;
  wire [0:19] cbx_1__1__23_chanx_left_out;
  wire [0:19] cbx_1__1__23_chanx_right_out;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__24_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__24_ccff_tail;
  wire [0:19] cbx_1__1__24_chanx_left_out;
  wire [0:19] cbx_1__1__24_chanx_right_out;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__25_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__25_ccff_tail;
  wire [0:19] cbx_1__1__25_chanx_left_out;
  wire [0:19] cbx_1__1__25_chanx_right_out;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__26_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__26_ccff_tail;
  wire [0:19] cbx_1__1__26_chanx_left_out;
  wire [0:19] cbx_1__1__26_chanx_right_out;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__27_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__27_ccff_tail;
  wire [0:19] cbx_1__1__27_chanx_left_out;
  wire [0:19] cbx_1__1__27_chanx_right_out;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__28_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__28_ccff_tail;
  wire [0:19] cbx_1__1__28_chanx_left_out;
  wire [0:19] cbx_1__1__28_chanx_right_out;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__29_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__29_ccff_tail;
  wire [0:19] cbx_1__1__29_chanx_left_out;
  wire [0:19] cbx_1__1__29_chanx_right_out;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__2_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__2_ccff_tail;
  wire [0:19] cbx_1__1__2_chanx_left_out;
  wire [0:19] cbx_1__1__2_chanx_right_out;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__30_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__30_ccff_tail;
  wire [0:19] cbx_1__1__30_chanx_left_out;
  wire [0:19] cbx_1__1__30_chanx_right_out;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__31_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__31_ccff_tail;
  wire [0:19] cbx_1__1__31_chanx_left_out;
  wire [0:19] cbx_1__1__31_chanx_right_out;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__32_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__32_ccff_tail;
  wire [0:19] cbx_1__1__32_chanx_left_out;
  wire [0:19] cbx_1__1__32_chanx_right_out;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__33_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__33_ccff_tail;
  wire [0:19] cbx_1__1__33_chanx_left_out;
  wire [0:19] cbx_1__1__33_chanx_right_out;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__34_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__34_ccff_tail;
  wire [0:19] cbx_1__1__34_chanx_left_out;
  wire [0:19] cbx_1__1__34_chanx_right_out;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__35_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__35_ccff_tail;
  wire [0:19] cbx_1__1__35_chanx_left_out;
  wire [0:19] cbx_1__1__35_chanx_right_out;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__36_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__36_ccff_tail;
  wire [0:19] cbx_1__1__36_chanx_left_out;
  wire [0:19] cbx_1__1__36_chanx_right_out;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__37_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__37_ccff_tail;
  wire [0:19] cbx_1__1__37_chanx_left_out;
  wire [0:19] cbx_1__1__37_chanx_right_out;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__38_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__38_ccff_tail;
  wire [0:19] cbx_1__1__38_chanx_left_out;
  wire [0:19] cbx_1__1__38_chanx_right_out;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__39_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__39_ccff_tail;
  wire [0:19] cbx_1__1__39_chanx_left_out;
  wire [0:19] cbx_1__1__39_chanx_right_out;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__3_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__3_ccff_tail;
  wire [0:19] cbx_1__1__3_chanx_left_out;
  wire [0:19] cbx_1__1__3_chanx_right_out;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__40_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__40_ccff_tail;
  wire [0:19] cbx_1__1__40_chanx_left_out;
  wire [0:19] cbx_1__1__40_chanx_right_out;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__41_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__41_ccff_tail;
  wire [0:19] cbx_1__1__41_chanx_left_out;
  wire [0:19] cbx_1__1__41_chanx_right_out;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__42_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__42_ccff_tail;
  wire [0:19] cbx_1__1__42_chanx_left_out;
  wire [0:19] cbx_1__1__42_chanx_right_out;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__43_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__43_ccff_tail;
  wire [0:19] cbx_1__1__43_chanx_left_out;
  wire [0:19] cbx_1__1__43_chanx_right_out;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__44_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__44_ccff_tail;
  wire [0:19] cbx_1__1__44_chanx_left_out;
  wire [0:19] cbx_1__1__44_chanx_right_out;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__45_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__45_ccff_tail;
  wire [0:19] cbx_1__1__45_chanx_left_out;
  wire [0:19] cbx_1__1__45_chanx_right_out;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__46_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__46_ccff_tail;
  wire [0:19] cbx_1__1__46_chanx_left_out;
  wire [0:19] cbx_1__1__46_chanx_right_out;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__47_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__47_ccff_tail;
  wire [0:19] cbx_1__1__47_chanx_left_out;
  wire [0:19] cbx_1__1__47_chanx_right_out;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__48_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__48_ccff_tail;
  wire [0:19] cbx_1__1__48_chanx_left_out;
  wire [0:19] cbx_1__1__48_chanx_right_out;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__49_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__49_ccff_tail;
  wire [0:19] cbx_1__1__49_chanx_left_out;
  wire [0:19] cbx_1__1__49_chanx_right_out;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__4_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__4_ccff_tail;
  wire [0:19] cbx_1__1__4_chanx_left_out;
  wire [0:19] cbx_1__1__4_chanx_right_out;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__50_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__50_ccff_tail;
  wire [0:19] cbx_1__1__50_chanx_left_out;
  wire [0:19] cbx_1__1__50_chanx_right_out;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__51_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__51_ccff_tail;
  wire [0:19] cbx_1__1__51_chanx_left_out;
  wire [0:19] cbx_1__1__51_chanx_right_out;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__52_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__52_ccff_tail;
  wire [0:19] cbx_1__1__52_chanx_left_out;
  wire [0:19] cbx_1__1__52_chanx_right_out;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__53_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__53_ccff_tail;
  wire [0:19] cbx_1__1__53_chanx_left_out;
  wire [0:19] cbx_1__1__53_chanx_right_out;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__54_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__54_ccff_tail;
  wire [0:19] cbx_1__1__54_chanx_left_out;
  wire [0:19] cbx_1__1__54_chanx_right_out;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__55_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__55_ccff_tail;
  wire [0:19] cbx_1__1__55_chanx_left_out;
  wire [0:19] cbx_1__1__55_chanx_right_out;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__5_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__5_ccff_tail;
  wire [0:19] cbx_1__1__5_chanx_left_out;
  wire [0:19] cbx_1__1__5_chanx_right_out;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__6_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__6_ccff_tail;
  wire [0:19] cbx_1__1__6_chanx_left_out;
  wire [0:19] cbx_1__1__6_chanx_right_out;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__7_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__7_ccff_tail;
  wire [0:19] cbx_1__1__7_chanx_left_out;
  wire [0:19] cbx_1__1__7_chanx_right_out;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__8_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__8_ccff_tail;
  wire [0:19] cbx_1__1__8_chanx_left_out;
  wire [0:19] cbx_1__1__8_chanx_right_out;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_0_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_10_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_11_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_12_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_13_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_14_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_15_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_1_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_2_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_3_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_4_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_5_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_6_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_7_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_8_;
  wire [0:0] cbx_1__1__9_bottom_grid_pin_9_;
  wire [0:0] cbx_1__1__9_ccff_tail;
  wire [0:19] cbx_1__1__9_chanx_left_out;
  wire [0:19] cbx_1__1__9_chanx_right_out;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__0_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__0_ccff_tail;
  wire [0:19] cbx_1__8__0_chanx_left_out;
  wire [0:19] cbx_1__8__0_chanx_right_out;
  wire [0:0] cbx_1__8__0_top_grid_pin_0_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__1_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__1_ccff_tail;
  wire [0:19] cbx_1__8__1_chanx_left_out;
  wire [0:19] cbx_1__8__1_chanx_right_out;
  wire [0:0] cbx_1__8__1_top_grid_pin_0_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__2_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__2_ccff_tail;
  wire [0:19] cbx_1__8__2_chanx_left_out;
  wire [0:19] cbx_1__8__2_chanx_right_out;
  wire [0:0] cbx_1__8__2_top_grid_pin_0_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__3_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__3_ccff_tail;
  wire [0:19] cbx_1__8__3_chanx_left_out;
  wire [0:19] cbx_1__8__3_chanx_right_out;
  wire [0:0] cbx_1__8__3_top_grid_pin_0_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__4_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__4_ccff_tail;
  wire [0:19] cbx_1__8__4_chanx_left_out;
  wire [0:19] cbx_1__8__4_chanx_right_out;
  wire [0:0] cbx_1__8__4_top_grid_pin_0_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__5_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__5_ccff_tail;
  wire [0:19] cbx_1__8__5_chanx_left_out;
  wire [0:19] cbx_1__8__5_chanx_right_out;
  wire [0:0] cbx_1__8__5_top_grid_pin_0_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__6_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__6_ccff_tail;
  wire [0:19] cbx_1__8__6_chanx_left_out;
  wire [0:19] cbx_1__8__6_chanx_right_out;
  wire [0:0] cbx_1__8__6_top_grid_pin_0_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_0_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_10_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_11_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_12_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_13_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_14_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_15_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_1_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_2_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_3_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_4_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_5_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_6_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_7_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_8_;
  wire [0:0] cbx_1__8__7_bottom_grid_pin_9_;
  wire [0:0] cbx_1__8__7_ccff_tail;
  wire [0:19] cbx_1__8__7_chanx_left_out;
  wire [0:19] cbx_1__8__7_chanx_right_out;
  wire [0:0] cbx_1__8__7_top_grid_pin_0_;
  wire [0:0] cby_0__1__0_ccff_tail;
  wire [0:19] cby_0__1__0_chany_bottom_out;
  wire [0:19] cby_0__1__0_chany_top_out;
  wire [0:0] cby_0__1__0_left_grid_pin_0_;
  wire [0:0] cby_0__1__1_ccff_tail;
  wire [0:19] cby_0__1__1_chany_bottom_out;
  wire [0:19] cby_0__1__1_chany_top_out;
  wire [0:0] cby_0__1__1_left_grid_pin_0_;
  wire [0:0] cby_0__1__2_ccff_tail;
  wire [0:19] cby_0__1__2_chany_bottom_out;
  wire [0:19] cby_0__1__2_chany_top_out;
  wire [0:0] cby_0__1__2_left_grid_pin_0_;
  wire [0:0] cby_0__1__3_ccff_tail;
  wire [0:19] cby_0__1__3_chany_bottom_out;
  wire [0:19] cby_0__1__3_chany_top_out;
  wire [0:0] cby_0__1__3_left_grid_pin_0_;
  wire [0:0] cby_0__1__4_ccff_tail;
  wire [0:19] cby_0__1__4_chany_bottom_out;
  wire [0:19] cby_0__1__4_chany_top_out;
  wire [0:0] cby_0__1__4_left_grid_pin_0_;
  wire [0:0] cby_0__1__5_ccff_tail;
  wire [0:19] cby_0__1__5_chany_bottom_out;
  wire [0:19] cby_0__1__5_chany_top_out;
  wire [0:0] cby_0__1__5_left_grid_pin_0_;
  wire [0:0] cby_0__1__6_ccff_tail;
  wire [0:19] cby_0__1__6_chany_bottom_out;
  wire [0:19] cby_0__1__6_chany_top_out;
  wire [0:0] cby_0__1__6_left_grid_pin_0_;
  wire [0:0] cby_0__1__7_ccff_tail;
  wire [0:19] cby_0__1__7_chany_bottom_out;
  wire [0:19] cby_0__1__7_chany_top_out;
  wire [0:0] cby_0__1__7_left_grid_pin_0_;
  wire [0:0] cby_1__1__0_ccff_tail;
  wire [0:19] cby_1__1__0_chany_bottom_out;
  wire [0:19] cby_1__1__0_chany_top_out;
  wire [0:0] cby_1__1__0_left_grid_pin_16_;
  wire [0:0] cby_1__1__0_left_grid_pin_17_;
  wire [0:0] cby_1__1__0_left_grid_pin_18_;
  wire [0:0] cby_1__1__0_left_grid_pin_19_;
  wire [0:0] cby_1__1__0_left_grid_pin_20_;
  wire [0:0] cby_1__1__0_left_grid_pin_21_;
  wire [0:0] cby_1__1__0_left_grid_pin_22_;
  wire [0:0] cby_1__1__0_left_grid_pin_23_;
  wire [0:0] cby_1__1__0_left_grid_pin_24_;
  wire [0:0] cby_1__1__0_left_grid_pin_25_;
  wire [0:0] cby_1__1__0_left_grid_pin_26_;
  wire [0:0] cby_1__1__0_left_grid_pin_27_;
  wire [0:0] cby_1__1__0_left_grid_pin_28_;
  wire [0:0] cby_1__1__0_left_grid_pin_29_;
  wire [0:0] cby_1__1__0_left_grid_pin_30_;
  wire [0:0] cby_1__1__0_left_grid_pin_31_;
  wire [0:0] cby_1__1__10_ccff_tail;
  wire [0:19] cby_1__1__10_chany_bottom_out;
  wire [0:19] cby_1__1__10_chany_top_out;
  wire [0:0] cby_1__1__10_left_grid_pin_16_;
  wire [0:0] cby_1__1__10_left_grid_pin_17_;
  wire [0:0] cby_1__1__10_left_grid_pin_18_;
  wire [0:0] cby_1__1__10_left_grid_pin_19_;
  wire [0:0] cby_1__1__10_left_grid_pin_20_;
  wire [0:0] cby_1__1__10_left_grid_pin_21_;
  wire [0:0] cby_1__1__10_left_grid_pin_22_;
  wire [0:0] cby_1__1__10_left_grid_pin_23_;
  wire [0:0] cby_1__1__10_left_grid_pin_24_;
  wire [0:0] cby_1__1__10_left_grid_pin_25_;
  wire [0:0] cby_1__1__10_left_grid_pin_26_;
  wire [0:0] cby_1__1__10_left_grid_pin_27_;
  wire [0:0] cby_1__1__10_left_grid_pin_28_;
  wire [0:0] cby_1__1__10_left_grid_pin_29_;
  wire [0:0] cby_1__1__10_left_grid_pin_30_;
  wire [0:0] cby_1__1__10_left_grid_pin_31_;
  wire [0:0] cby_1__1__11_ccff_tail;
  wire [0:19] cby_1__1__11_chany_bottom_out;
  wire [0:19] cby_1__1__11_chany_top_out;
  wire [0:0] cby_1__1__11_left_grid_pin_16_;
  wire [0:0] cby_1__1__11_left_grid_pin_17_;
  wire [0:0] cby_1__1__11_left_grid_pin_18_;
  wire [0:0] cby_1__1__11_left_grid_pin_19_;
  wire [0:0] cby_1__1__11_left_grid_pin_20_;
  wire [0:0] cby_1__1__11_left_grid_pin_21_;
  wire [0:0] cby_1__1__11_left_grid_pin_22_;
  wire [0:0] cby_1__1__11_left_grid_pin_23_;
  wire [0:0] cby_1__1__11_left_grid_pin_24_;
  wire [0:0] cby_1__1__11_left_grid_pin_25_;
  wire [0:0] cby_1__1__11_left_grid_pin_26_;
  wire [0:0] cby_1__1__11_left_grid_pin_27_;
  wire [0:0] cby_1__1__11_left_grid_pin_28_;
  wire [0:0] cby_1__1__11_left_grid_pin_29_;
  wire [0:0] cby_1__1__11_left_grid_pin_30_;
  wire [0:0] cby_1__1__11_left_grid_pin_31_;
  wire [0:0] cby_1__1__12_ccff_tail;
  wire [0:19] cby_1__1__12_chany_bottom_out;
  wire [0:19] cby_1__1__12_chany_top_out;
  wire [0:0] cby_1__1__12_left_grid_pin_16_;
  wire [0:0] cby_1__1__12_left_grid_pin_17_;
  wire [0:0] cby_1__1__12_left_grid_pin_18_;
  wire [0:0] cby_1__1__12_left_grid_pin_19_;
  wire [0:0] cby_1__1__12_left_grid_pin_20_;
  wire [0:0] cby_1__1__12_left_grid_pin_21_;
  wire [0:0] cby_1__1__12_left_grid_pin_22_;
  wire [0:0] cby_1__1__12_left_grid_pin_23_;
  wire [0:0] cby_1__1__12_left_grid_pin_24_;
  wire [0:0] cby_1__1__12_left_grid_pin_25_;
  wire [0:0] cby_1__1__12_left_grid_pin_26_;
  wire [0:0] cby_1__1__12_left_grid_pin_27_;
  wire [0:0] cby_1__1__12_left_grid_pin_28_;
  wire [0:0] cby_1__1__12_left_grid_pin_29_;
  wire [0:0] cby_1__1__12_left_grid_pin_30_;
  wire [0:0] cby_1__1__12_left_grid_pin_31_;
  wire [0:0] cby_1__1__13_ccff_tail;
  wire [0:19] cby_1__1__13_chany_bottom_out;
  wire [0:19] cby_1__1__13_chany_top_out;
  wire [0:0] cby_1__1__13_left_grid_pin_16_;
  wire [0:0] cby_1__1__13_left_grid_pin_17_;
  wire [0:0] cby_1__1__13_left_grid_pin_18_;
  wire [0:0] cby_1__1__13_left_grid_pin_19_;
  wire [0:0] cby_1__1__13_left_grid_pin_20_;
  wire [0:0] cby_1__1__13_left_grid_pin_21_;
  wire [0:0] cby_1__1__13_left_grid_pin_22_;
  wire [0:0] cby_1__1__13_left_grid_pin_23_;
  wire [0:0] cby_1__1__13_left_grid_pin_24_;
  wire [0:0] cby_1__1__13_left_grid_pin_25_;
  wire [0:0] cby_1__1__13_left_grid_pin_26_;
  wire [0:0] cby_1__1__13_left_grid_pin_27_;
  wire [0:0] cby_1__1__13_left_grid_pin_28_;
  wire [0:0] cby_1__1__13_left_grid_pin_29_;
  wire [0:0] cby_1__1__13_left_grid_pin_30_;
  wire [0:0] cby_1__1__13_left_grid_pin_31_;
  wire [0:0] cby_1__1__14_ccff_tail;
  wire [0:19] cby_1__1__14_chany_bottom_out;
  wire [0:19] cby_1__1__14_chany_top_out;
  wire [0:0] cby_1__1__14_left_grid_pin_16_;
  wire [0:0] cby_1__1__14_left_grid_pin_17_;
  wire [0:0] cby_1__1__14_left_grid_pin_18_;
  wire [0:0] cby_1__1__14_left_grid_pin_19_;
  wire [0:0] cby_1__1__14_left_grid_pin_20_;
  wire [0:0] cby_1__1__14_left_grid_pin_21_;
  wire [0:0] cby_1__1__14_left_grid_pin_22_;
  wire [0:0] cby_1__1__14_left_grid_pin_23_;
  wire [0:0] cby_1__1__14_left_grid_pin_24_;
  wire [0:0] cby_1__1__14_left_grid_pin_25_;
  wire [0:0] cby_1__1__14_left_grid_pin_26_;
  wire [0:0] cby_1__1__14_left_grid_pin_27_;
  wire [0:0] cby_1__1__14_left_grid_pin_28_;
  wire [0:0] cby_1__1__14_left_grid_pin_29_;
  wire [0:0] cby_1__1__14_left_grid_pin_30_;
  wire [0:0] cby_1__1__14_left_grid_pin_31_;
  wire [0:0] cby_1__1__15_ccff_tail;
  wire [0:19] cby_1__1__15_chany_bottom_out;
  wire [0:19] cby_1__1__15_chany_top_out;
  wire [0:0] cby_1__1__15_left_grid_pin_16_;
  wire [0:0] cby_1__1__15_left_grid_pin_17_;
  wire [0:0] cby_1__1__15_left_grid_pin_18_;
  wire [0:0] cby_1__1__15_left_grid_pin_19_;
  wire [0:0] cby_1__1__15_left_grid_pin_20_;
  wire [0:0] cby_1__1__15_left_grid_pin_21_;
  wire [0:0] cby_1__1__15_left_grid_pin_22_;
  wire [0:0] cby_1__1__15_left_grid_pin_23_;
  wire [0:0] cby_1__1__15_left_grid_pin_24_;
  wire [0:0] cby_1__1__15_left_grid_pin_25_;
  wire [0:0] cby_1__1__15_left_grid_pin_26_;
  wire [0:0] cby_1__1__15_left_grid_pin_27_;
  wire [0:0] cby_1__1__15_left_grid_pin_28_;
  wire [0:0] cby_1__1__15_left_grid_pin_29_;
  wire [0:0] cby_1__1__15_left_grid_pin_30_;
  wire [0:0] cby_1__1__15_left_grid_pin_31_;
  wire [0:0] cby_1__1__16_ccff_tail;
  wire [0:19] cby_1__1__16_chany_bottom_out;
  wire [0:19] cby_1__1__16_chany_top_out;
  wire [0:0] cby_1__1__16_left_grid_pin_16_;
  wire [0:0] cby_1__1__16_left_grid_pin_17_;
  wire [0:0] cby_1__1__16_left_grid_pin_18_;
  wire [0:0] cby_1__1__16_left_grid_pin_19_;
  wire [0:0] cby_1__1__16_left_grid_pin_20_;
  wire [0:0] cby_1__1__16_left_grid_pin_21_;
  wire [0:0] cby_1__1__16_left_grid_pin_22_;
  wire [0:0] cby_1__1__16_left_grid_pin_23_;
  wire [0:0] cby_1__1__16_left_grid_pin_24_;
  wire [0:0] cby_1__1__16_left_grid_pin_25_;
  wire [0:0] cby_1__1__16_left_grid_pin_26_;
  wire [0:0] cby_1__1__16_left_grid_pin_27_;
  wire [0:0] cby_1__1__16_left_grid_pin_28_;
  wire [0:0] cby_1__1__16_left_grid_pin_29_;
  wire [0:0] cby_1__1__16_left_grid_pin_30_;
  wire [0:0] cby_1__1__16_left_grid_pin_31_;
  wire [0:0] cby_1__1__17_ccff_tail;
  wire [0:19] cby_1__1__17_chany_bottom_out;
  wire [0:19] cby_1__1__17_chany_top_out;
  wire [0:0] cby_1__1__17_left_grid_pin_16_;
  wire [0:0] cby_1__1__17_left_grid_pin_17_;
  wire [0:0] cby_1__1__17_left_grid_pin_18_;
  wire [0:0] cby_1__1__17_left_grid_pin_19_;
  wire [0:0] cby_1__1__17_left_grid_pin_20_;
  wire [0:0] cby_1__1__17_left_grid_pin_21_;
  wire [0:0] cby_1__1__17_left_grid_pin_22_;
  wire [0:0] cby_1__1__17_left_grid_pin_23_;
  wire [0:0] cby_1__1__17_left_grid_pin_24_;
  wire [0:0] cby_1__1__17_left_grid_pin_25_;
  wire [0:0] cby_1__1__17_left_grid_pin_26_;
  wire [0:0] cby_1__1__17_left_grid_pin_27_;
  wire [0:0] cby_1__1__17_left_grid_pin_28_;
  wire [0:0] cby_1__1__17_left_grid_pin_29_;
  wire [0:0] cby_1__1__17_left_grid_pin_30_;
  wire [0:0] cby_1__1__17_left_grid_pin_31_;
  wire [0:0] cby_1__1__18_ccff_tail;
  wire [0:19] cby_1__1__18_chany_bottom_out;
  wire [0:19] cby_1__1__18_chany_top_out;
  wire [0:0] cby_1__1__18_left_grid_pin_16_;
  wire [0:0] cby_1__1__18_left_grid_pin_17_;
  wire [0:0] cby_1__1__18_left_grid_pin_18_;
  wire [0:0] cby_1__1__18_left_grid_pin_19_;
  wire [0:0] cby_1__1__18_left_grid_pin_20_;
  wire [0:0] cby_1__1__18_left_grid_pin_21_;
  wire [0:0] cby_1__1__18_left_grid_pin_22_;
  wire [0:0] cby_1__1__18_left_grid_pin_23_;
  wire [0:0] cby_1__1__18_left_grid_pin_24_;
  wire [0:0] cby_1__1__18_left_grid_pin_25_;
  wire [0:0] cby_1__1__18_left_grid_pin_26_;
  wire [0:0] cby_1__1__18_left_grid_pin_27_;
  wire [0:0] cby_1__1__18_left_grid_pin_28_;
  wire [0:0] cby_1__1__18_left_grid_pin_29_;
  wire [0:0] cby_1__1__18_left_grid_pin_30_;
  wire [0:0] cby_1__1__18_left_grid_pin_31_;
  wire [0:0] cby_1__1__19_ccff_tail;
  wire [0:19] cby_1__1__19_chany_bottom_out;
  wire [0:19] cby_1__1__19_chany_top_out;
  wire [0:0] cby_1__1__19_left_grid_pin_16_;
  wire [0:0] cby_1__1__19_left_grid_pin_17_;
  wire [0:0] cby_1__1__19_left_grid_pin_18_;
  wire [0:0] cby_1__1__19_left_grid_pin_19_;
  wire [0:0] cby_1__1__19_left_grid_pin_20_;
  wire [0:0] cby_1__1__19_left_grid_pin_21_;
  wire [0:0] cby_1__1__19_left_grid_pin_22_;
  wire [0:0] cby_1__1__19_left_grid_pin_23_;
  wire [0:0] cby_1__1__19_left_grid_pin_24_;
  wire [0:0] cby_1__1__19_left_grid_pin_25_;
  wire [0:0] cby_1__1__19_left_grid_pin_26_;
  wire [0:0] cby_1__1__19_left_grid_pin_27_;
  wire [0:0] cby_1__1__19_left_grid_pin_28_;
  wire [0:0] cby_1__1__19_left_grid_pin_29_;
  wire [0:0] cby_1__1__19_left_grid_pin_30_;
  wire [0:0] cby_1__1__19_left_grid_pin_31_;
  wire [0:0] cby_1__1__1_ccff_tail;
  wire [0:19] cby_1__1__1_chany_bottom_out;
  wire [0:19] cby_1__1__1_chany_top_out;
  wire [0:0] cby_1__1__1_left_grid_pin_16_;
  wire [0:0] cby_1__1__1_left_grid_pin_17_;
  wire [0:0] cby_1__1__1_left_grid_pin_18_;
  wire [0:0] cby_1__1__1_left_grid_pin_19_;
  wire [0:0] cby_1__1__1_left_grid_pin_20_;
  wire [0:0] cby_1__1__1_left_grid_pin_21_;
  wire [0:0] cby_1__1__1_left_grid_pin_22_;
  wire [0:0] cby_1__1__1_left_grid_pin_23_;
  wire [0:0] cby_1__1__1_left_grid_pin_24_;
  wire [0:0] cby_1__1__1_left_grid_pin_25_;
  wire [0:0] cby_1__1__1_left_grid_pin_26_;
  wire [0:0] cby_1__1__1_left_grid_pin_27_;
  wire [0:0] cby_1__1__1_left_grid_pin_28_;
  wire [0:0] cby_1__1__1_left_grid_pin_29_;
  wire [0:0] cby_1__1__1_left_grid_pin_30_;
  wire [0:0] cby_1__1__1_left_grid_pin_31_;
  wire [0:0] cby_1__1__20_ccff_tail;
  wire [0:19] cby_1__1__20_chany_bottom_out;
  wire [0:19] cby_1__1__20_chany_top_out;
  wire [0:0] cby_1__1__20_left_grid_pin_16_;
  wire [0:0] cby_1__1__20_left_grid_pin_17_;
  wire [0:0] cby_1__1__20_left_grid_pin_18_;
  wire [0:0] cby_1__1__20_left_grid_pin_19_;
  wire [0:0] cby_1__1__20_left_grid_pin_20_;
  wire [0:0] cby_1__1__20_left_grid_pin_21_;
  wire [0:0] cby_1__1__20_left_grid_pin_22_;
  wire [0:0] cby_1__1__20_left_grid_pin_23_;
  wire [0:0] cby_1__1__20_left_grid_pin_24_;
  wire [0:0] cby_1__1__20_left_grid_pin_25_;
  wire [0:0] cby_1__1__20_left_grid_pin_26_;
  wire [0:0] cby_1__1__20_left_grid_pin_27_;
  wire [0:0] cby_1__1__20_left_grid_pin_28_;
  wire [0:0] cby_1__1__20_left_grid_pin_29_;
  wire [0:0] cby_1__1__20_left_grid_pin_30_;
  wire [0:0] cby_1__1__20_left_grid_pin_31_;
  wire [0:0] cby_1__1__21_ccff_tail;
  wire [0:19] cby_1__1__21_chany_bottom_out;
  wire [0:19] cby_1__1__21_chany_top_out;
  wire [0:0] cby_1__1__21_left_grid_pin_16_;
  wire [0:0] cby_1__1__21_left_grid_pin_17_;
  wire [0:0] cby_1__1__21_left_grid_pin_18_;
  wire [0:0] cby_1__1__21_left_grid_pin_19_;
  wire [0:0] cby_1__1__21_left_grid_pin_20_;
  wire [0:0] cby_1__1__21_left_grid_pin_21_;
  wire [0:0] cby_1__1__21_left_grid_pin_22_;
  wire [0:0] cby_1__1__21_left_grid_pin_23_;
  wire [0:0] cby_1__1__21_left_grid_pin_24_;
  wire [0:0] cby_1__1__21_left_grid_pin_25_;
  wire [0:0] cby_1__1__21_left_grid_pin_26_;
  wire [0:0] cby_1__1__21_left_grid_pin_27_;
  wire [0:0] cby_1__1__21_left_grid_pin_28_;
  wire [0:0] cby_1__1__21_left_grid_pin_29_;
  wire [0:0] cby_1__1__21_left_grid_pin_30_;
  wire [0:0] cby_1__1__21_left_grid_pin_31_;
  wire [0:0] cby_1__1__22_ccff_tail;
  wire [0:19] cby_1__1__22_chany_bottom_out;
  wire [0:19] cby_1__1__22_chany_top_out;
  wire [0:0] cby_1__1__22_left_grid_pin_16_;
  wire [0:0] cby_1__1__22_left_grid_pin_17_;
  wire [0:0] cby_1__1__22_left_grid_pin_18_;
  wire [0:0] cby_1__1__22_left_grid_pin_19_;
  wire [0:0] cby_1__1__22_left_grid_pin_20_;
  wire [0:0] cby_1__1__22_left_grid_pin_21_;
  wire [0:0] cby_1__1__22_left_grid_pin_22_;
  wire [0:0] cby_1__1__22_left_grid_pin_23_;
  wire [0:0] cby_1__1__22_left_grid_pin_24_;
  wire [0:0] cby_1__1__22_left_grid_pin_25_;
  wire [0:0] cby_1__1__22_left_grid_pin_26_;
  wire [0:0] cby_1__1__22_left_grid_pin_27_;
  wire [0:0] cby_1__1__22_left_grid_pin_28_;
  wire [0:0] cby_1__1__22_left_grid_pin_29_;
  wire [0:0] cby_1__1__22_left_grid_pin_30_;
  wire [0:0] cby_1__1__22_left_grid_pin_31_;
  wire [0:0] cby_1__1__23_ccff_tail;
  wire [0:19] cby_1__1__23_chany_bottom_out;
  wire [0:19] cby_1__1__23_chany_top_out;
  wire [0:0] cby_1__1__23_left_grid_pin_16_;
  wire [0:0] cby_1__1__23_left_grid_pin_17_;
  wire [0:0] cby_1__1__23_left_grid_pin_18_;
  wire [0:0] cby_1__1__23_left_grid_pin_19_;
  wire [0:0] cby_1__1__23_left_grid_pin_20_;
  wire [0:0] cby_1__1__23_left_grid_pin_21_;
  wire [0:0] cby_1__1__23_left_grid_pin_22_;
  wire [0:0] cby_1__1__23_left_grid_pin_23_;
  wire [0:0] cby_1__1__23_left_grid_pin_24_;
  wire [0:0] cby_1__1__23_left_grid_pin_25_;
  wire [0:0] cby_1__1__23_left_grid_pin_26_;
  wire [0:0] cby_1__1__23_left_grid_pin_27_;
  wire [0:0] cby_1__1__23_left_grid_pin_28_;
  wire [0:0] cby_1__1__23_left_grid_pin_29_;
  wire [0:0] cby_1__1__23_left_grid_pin_30_;
  wire [0:0] cby_1__1__23_left_grid_pin_31_;
  wire [0:0] cby_1__1__24_ccff_tail;
  wire [0:19] cby_1__1__24_chany_bottom_out;
  wire [0:19] cby_1__1__24_chany_top_out;
  wire [0:0] cby_1__1__24_left_grid_pin_16_;
  wire [0:0] cby_1__1__24_left_grid_pin_17_;
  wire [0:0] cby_1__1__24_left_grid_pin_18_;
  wire [0:0] cby_1__1__24_left_grid_pin_19_;
  wire [0:0] cby_1__1__24_left_grid_pin_20_;
  wire [0:0] cby_1__1__24_left_grid_pin_21_;
  wire [0:0] cby_1__1__24_left_grid_pin_22_;
  wire [0:0] cby_1__1__24_left_grid_pin_23_;
  wire [0:0] cby_1__1__24_left_grid_pin_24_;
  wire [0:0] cby_1__1__24_left_grid_pin_25_;
  wire [0:0] cby_1__1__24_left_grid_pin_26_;
  wire [0:0] cby_1__1__24_left_grid_pin_27_;
  wire [0:0] cby_1__1__24_left_grid_pin_28_;
  wire [0:0] cby_1__1__24_left_grid_pin_29_;
  wire [0:0] cby_1__1__24_left_grid_pin_30_;
  wire [0:0] cby_1__1__24_left_grid_pin_31_;
  wire [0:0] cby_1__1__25_ccff_tail;
  wire [0:19] cby_1__1__25_chany_bottom_out;
  wire [0:19] cby_1__1__25_chany_top_out;
  wire [0:0] cby_1__1__25_left_grid_pin_16_;
  wire [0:0] cby_1__1__25_left_grid_pin_17_;
  wire [0:0] cby_1__1__25_left_grid_pin_18_;
  wire [0:0] cby_1__1__25_left_grid_pin_19_;
  wire [0:0] cby_1__1__25_left_grid_pin_20_;
  wire [0:0] cby_1__1__25_left_grid_pin_21_;
  wire [0:0] cby_1__1__25_left_grid_pin_22_;
  wire [0:0] cby_1__1__25_left_grid_pin_23_;
  wire [0:0] cby_1__1__25_left_grid_pin_24_;
  wire [0:0] cby_1__1__25_left_grid_pin_25_;
  wire [0:0] cby_1__1__25_left_grid_pin_26_;
  wire [0:0] cby_1__1__25_left_grid_pin_27_;
  wire [0:0] cby_1__1__25_left_grid_pin_28_;
  wire [0:0] cby_1__1__25_left_grid_pin_29_;
  wire [0:0] cby_1__1__25_left_grid_pin_30_;
  wire [0:0] cby_1__1__25_left_grid_pin_31_;
  wire [0:0] cby_1__1__26_ccff_tail;
  wire [0:19] cby_1__1__26_chany_bottom_out;
  wire [0:19] cby_1__1__26_chany_top_out;
  wire [0:0] cby_1__1__26_left_grid_pin_16_;
  wire [0:0] cby_1__1__26_left_grid_pin_17_;
  wire [0:0] cby_1__1__26_left_grid_pin_18_;
  wire [0:0] cby_1__1__26_left_grid_pin_19_;
  wire [0:0] cby_1__1__26_left_grid_pin_20_;
  wire [0:0] cby_1__1__26_left_grid_pin_21_;
  wire [0:0] cby_1__1__26_left_grid_pin_22_;
  wire [0:0] cby_1__1__26_left_grid_pin_23_;
  wire [0:0] cby_1__1__26_left_grid_pin_24_;
  wire [0:0] cby_1__1__26_left_grid_pin_25_;
  wire [0:0] cby_1__1__26_left_grid_pin_26_;
  wire [0:0] cby_1__1__26_left_grid_pin_27_;
  wire [0:0] cby_1__1__26_left_grid_pin_28_;
  wire [0:0] cby_1__1__26_left_grid_pin_29_;
  wire [0:0] cby_1__1__26_left_grid_pin_30_;
  wire [0:0] cby_1__1__26_left_grid_pin_31_;
  wire [0:0] cby_1__1__27_ccff_tail;
  wire [0:19] cby_1__1__27_chany_bottom_out;
  wire [0:19] cby_1__1__27_chany_top_out;
  wire [0:0] cby_1__1__27_left_grid_pin_16_;
  wire [0:0] cby_1__1__27_left_grid_pin_17_;
  wire [0:0] cby_1__1__27_left_grid_pin_18_;
  wire [0:0] cby_1__1__27_left_grid_pin_19_;
  wire [0:0] cby_1__1__27_left_grid_pin_20_;
  wire [0:0] cby_1__1__27_left_grid_pin_21_;
  wire [0:0] cby_1__1__27_left_grid_pin_22_;
  wire [0:0] cby_1__1__27_left_grid_pin_23_;
  wire [0:0] cby_1__1__27_left_grid_pin_24_;
  wire [0:0] cby_1__1__27_left_grid_pin_25_;
  wire [0:0] cby_1__1__27_left_grid_pin_26_;
  wire [0:0] cby_1__1__27_left_grid_pin_27_;
  wire [0:0] cby_1__1__27_left_grid_pin_28_;
  wire [0:0] cby_1__1__27_left_grid_pin_29_;
  wire [0:0] cby_1__1__27_left_grid_pin_30_;
  wire [0:0] cby_1__1__27_left_grid_pin_31_;
  wire [0:0] cby_1__1__28_ccff_tail;
  wire [0:19] cby_1__1__28_chany_bottom_out;
  wire [0:19] cby_1__1__28_chany_top_out;
  wire [0:0] cby_1__1__28_left_grid_pin_16_;
  wire [0:0] cby_1__1__28_left_grid_pin_17_;
  wire [0:0] cby_1__1__28_left_grid_pin_18_;
  wire [0:0] cby_1__1__28_left_grid_pin_19_;
  wire [0:0] cby_1__1__28_left_grid_pin_20_;
  wire [0:0] cby_1__1__28_left_grid_pin_21_;
  wire [0:0] cby_1__1__28_left_grid_pin_22_;
  wire [0:0] cby_1__1__28_left_grid_pin_23_;
  wire [0:0] cby_1__1__28_left_grid_pin_24_;
  wire [0:0] cby_1__1__28_left_grid_pin_25_;
  wire [0:0] cby_1__1__28_left_grid_pin_26_;
  wire [0:0] cby_1__1__28_left_grid_pin_27_;
  wire [0:0] cby_1__1__28_left_grid_pin_28_;
  wire [0:0] cby_1__1__28_left_grid_pin_29_;
  wire [0:0] cby_1__1__28_left_grid_pin_30_;
  wire [0:0] cby_1__1__28_left_grid_pin_31_;
  wire [0:0] cby_1__1__29_ccff_tail;
  wire [0:19] cby_1__1__29_chany_bottom_out;
  wire [0:19] cby_1__1__29_chany_top_out;
  wire [0:0] cby_1__1__29_left_grid_pin_16_;
  wire [0:0] cby_1__1__29_left_grid_pin_17_;
  wire [0:0] cby_1__1__29_left_grid_pin_18_;
  wire [0:0] cby_1__1__29_left_grid_pin_19_;
  wire [0:0] cby_1__1__29_left_grid_pin_20_;
  wire [0:0] cby_1__1__29_left_grid_pin_21_;
  wire [0:0] cby_1__1__29_left_grid_pin_22_;
  wire [0:0] cby_1__1__29_left_grid_pin_23_;
  wire [0:0] cby_1__1__29_left_grid_pin_24_;
  wire [0:0] cby_1__1__29_left_grid_pin_25_;
  wire [0:0] cby_1__1__29_left_grid_pin_26_;
  wire [0:0] cby_1__1__29_left_grid_pin_27_;
  wire [0:0] cby_1__1__29_left_grid_pin_28_;
  wire [0:0] cby_1__1__29_left_grid_pin_29_;
  wire [0:0] cby_1__1__29_left_grid_pin_30_;
  wire [0:0] cby_1__1__29_left_grid_pin_31_;
  wire [0:0] cby_1__1__2_ccff_tail;
  wire [0:19] cby_1__1__2_chany_bottom_out;
  wire [0:19] cby_1__1__2_chany_top_out;
  wire [0:0] cby_1__1__2_left_grid_pin_16_;
  wire [0:0] cby_1__1__2_left_grid_pin_17_;
  wire [0:0] cby_1__1__2_left_grid_pin_18_;
  wire [0:0] cby_1__1__2_left_grid_pin_19_;
  wire [0:0] cby_1__1__2_left_grid_pin_20_;
  wire [0:0] cby_1__1__2_left_grid_pin_21_;
  wire [0:0] cby_1__1__2_left_grid_pin_22_;
  wire [0:0] cby_1__1__2_left_grid_pin_23_;
  wire [0:0] cby_1__1__2_left_grid_pin_24_;
  wire [0:0] cby_1__1__2_left_grid_pin_25_;
  wire [0:0] cby_1__1__2_left_grid_pin_26_;
  wire [0:0] cby_1__1__2_left_grid_pin_27_;
  wire [0:0] cby_1__1__2_left_grid_pin_28_;
  wire [0:0] cby_1__1__2_left_grid_pin_29_;
  wire [0:0] cby_1__1__2_left_grid_pin_30_;
  wire [0:0] cby_1__1__2_left_grid_pin_31_;
  wire [0:0] cby_1__1__30_ccff_tail;
  wire [0:19] cby_1__1__30_chany_bottom_out;
  wire [0:19] cby_1__1__30_chany_top_out;
  wire [0:0] cby_1__1__30_left_grid_pin_16_;
  wire [0:0] cby_1__1__30_left_grid_pin_17_;
  wire [0:0] cby_1__1__30_left_grid_pin_18_;
  wire [0:0] cby_1__1__30_left_grid_pin_19_;
  wire [0:0] cby_1__1__30_left_grid_pin_20_;
  wire [0:0] cby_1__1__30_left_grid_pin_21_;
  wire [0:0] cby_1__1__30_left_grid_pin_22_;
  wire [0:0] cby_1__1__30_left_grid_pin_23_;
  wire [0:0] cby_1__1__30_left_grid_pin_24_;
  wire [0:0] cby_1__1__30_left_grid_pin_25_;
  wire [0:0] cby_1__1__30_left_grid_pin_26_;
  wire [0:0] cby_1__1__30_left_grid_pin_27_;
  wire [0:0] cby_1__1__30_left_grid_pin_28_;
  wire [0:0] cby_1__1__30_left_grid_pin_29_;
  wire [0:0] cby_1__1__30_left_grid_pin_30_;
  wire [0:0] cby_1__1__30_left_grid_pin_31_;
  wire [0:0] cby_1__1__31_ccff_tail;
  wire [0:19] cby_1__1__31_chany_bottom_out;
  wire [0:19] cby_1__1__31_chany_top_out;
  wire [0:0] cby_1__1__31_left_grid_pin_16_;
  wire [0:0] cby_1__1__31_left_grid_pin_17_;
  wire [0:0] cby_1__1__31_left_grid_pin_18_;
  wire [0:0] cby_1__1__31_left_grid_pin_19_;
  wire [0:0] cby_1__1__31_left_grid_pin_20_;
  wire [0:0] cby_1__1__31_left_grid_pin_21_;
  wire [0:0] cby_1__1__31_left_grid_pin_22_;
  wire [0:0] cby_1__1__31_left_grid_pin_23_;
  wire [0:0] cby_1__1__31_left_grid_pin_24_;
  wire [0:0] cby_1__1__31_left_grid_pin_25_;
  wire [0:0] cby_1__1__31_left_grid_pin_26_;
  wire [0:0] cby_1__1__31_left_grid_pin_27_;
  wire [0:0] cby_1__1__31_left_grid_pin_28_;
  wire [0:0] cby_1__1__31_left_grid_pin_29_;
  wire [0:0] cby_1__1__31_left_grid_pin_30_;
  wire [0:0] cby_1__1__31_left_grid_pin_31_;
  wire [0:0] cby_1__1__32_ccff_tail;
  wire [0:19] cby_1__1__32_chany_bottom_out;
  wire [0:19] cby_1__1__32_chany_top_out;
  wire [0:0] cby_1__1__32_left_grid_pin_16_;
  wire [0:0] cby_1__1__32_left_grid_pin_17_;
  wire [0:0] cby_1__1__32_left_grid_pin_18_;
  wire [0:0] cby_1__1__32_left_grid_pin_19_;
  wire [0:0] cby_1__1__32_left_grid_pin_20_;
  wire [0:0] cby_1__1__32_left_grid_pin_21_;
  wire [0:0] cby_1__1__32_left_grid_pin_22_;
  wire [0:0] cby_1__1__32_left_grid_pin_23_;
  wire [0:0] cby_1__1__32_left_grid_pin_24_;
  wire [0:0] cby_1__1__32_left_grid_pin_25_;
  wire [0:0] cby_1__1__32_left_grid_pin_26_;
  wire [0:0] cby_1__1__32_left_grid_pin_27_;
  wire [0:0] cby_1__1__32_left_grid_pin_28_;
  wire [0:0] cby_1__1__32_left_grid_pin_29_;
  wire [0:0] cby_1__1__32_left_grid_pin_30_;
  wire [0:0] cby_1__1__32_left_grid_pin_31_;
  wire [0:0] cby_1__1__33_ccff_tail;
  wire [0:19] cby_1__1__33_chany_bottom_out;
  wire [0:19] cby_1__1__33_chany_top_out;
  wire [0:0] cby_1__1__33_left_grid_pin_16_;
  wire [0:0] cby_1__1__33_left_grid_pin_17_;
  wire [0:0] cby_1__1__33_left_grid_pin_18_;
  wire [0:0] cby_1__1__33_left_grid_pin_19_;
  wire [0:0] cby_1__1__33_left_grid_pin_20_;
  wire [0:0] cby_1__1__33_left_grid_pin_21_;
  wire [0:0] cby_1__1__33_left_grid_pin_22_;
  wire [0:0] cby_1__1__33_left_grid_pin_23_;
  wire [0:0] cby_1__1__33_left_grid_pin_24_;
  wire [0:0] cby_1__1__33_left_grid_pin_25_;
  wire [0:0] cby_1__1__33_left_grid_pin_26_;
  wire [0:0] cby_1__1__33_left_grid_pin_27_;
  wire [0:0] cby_1__1__33_left_grid_pin_28_;
  wire [0:0] cby_1__1__33_left_grid_pin_29_;
  wire [0:0] cby_1__1__33_left_grid_pin_30_;
  wire [0:0] cby_1__1__33_left_grid_pin_31_;
  wire [0:0] cby_1__1__34_ccff_tail;
  wire [0:19] cby_1__1__34_chany_bottom_out;
  wire [0:19] cby_1__1__34_chany_top_out;
  wire [0:0] cby_1__1__34_left_grid_pin_16_;
  wire [0:0] cby_1__1__34_left_grid_pin_17_;
  wire [0:0] cby_1__1__34_left_grid_pin_18_;
  wire [0:0] cby_1__1__34_left_grid_pin_19_;
  wire [0:0] cby_1__1__34_left_grid_pin_20_;
  wire [0:0] cby_1__1__34_left_grid_pin_21_;
  wire [0:0] cby_1__1__34_left_grid_pin_22_;
  wire [0:0] cby_1__1__34_left_grid_pin_23_;
  wire [0:0] cby_1__1__34_left_grid_pin_24_;
  wire [0:0] cby_1__1__34_left_grid_pin_25_;
  wire [0:0] cby_1__1__34_left_grid_pin_26_;
  wire [0:0] cby_1__1__34_left_grid_pin_27_;
  wire [0:0] cby_1__1__34_left_grid_pin_28_;
  wire [0:0] cby_1__1__34_left_grid_pin_29_;
  wire [0:0] cby_1__1__34_left_grid_pin_30_;
  wire [0:0] cby_1__1__34_left_grid_pin_31_;
  wire [0:0] cby_1__1__35_ccff_tail;
  wire [0:19] cby_1__1__35_chany_bottom_out;
  wire [0:19] cby_1__1__35_chany_top_out;
  wire [0:0] cby_1__1__35_left_grid_pin_16_;
  wire [0:0] cby_1__1__35_left_grid_pin_17_;
  wire [0:0] cby_1__1__35_left_grid_pin_18_;
  wire [0:0] cby_1__1__35_left_grid_pin_19_;
  wire [0:0] cby_1__1__35_left_grid_pin_20_;
  wire [0:0] cby_1__1__35_left_grid_pin_21_;
  wire [0:0] cby_1__1__35_left_grid_pin_22_;
  wire [0:0] cby_1__1__35_left_grid_pin_23_;
  wire [0:0] cby_1__1__35_left_grid_pin_24_;
  wire [0:0] cby_1__1__35_left_grid_pin_25_;
  wire [0:0] cby_1__1__35_left_grid_pin_26_;
  wire [0:0] cby_1__1__35_left_grid_pin_27_;
  wire [0:0] cby_1__1__35_left_grid_pin_28_;
  wire [0:0] cby_1__1__35_left_grid_pin_29_;
  wire [0:0] cby_1__1__35_left_grid_pin_30_;
  wire [0:0] cby_1__1__35_left_grid_pin_31_;
  wire [0:0] cby_1__1__36_ccff_tail;
  wire [0:19] cby_1__1__36_chany_bottom_out;
  wire [0:19] cby_1__1__36_chany_top_out;
  wire [0:0] cby_1__1__36_left_grid_pin_16_;
  wire [0:0] cby_1__1__36_left_grid_pin_17_;
  wire [0:0] cby_1__1__36_left_grid_pin_18_;
  wire [0:0] cby_1__1__36_left_grid_pin_19_;
  wire [0:0] cby_1__1__36_left_grid_pin_20_;
  wire [0:0] cby_1__1__36_left_grid_pin_21_;
  wire [0:0] cby_1__1__36_left_grid_pin_22_;
  wire [0:0] cby_1__1__36_left_grid_pin_23_;
  wire [0:0] cby_1__1__36_left_grid_pin_24_;
  wire [0:0] cby_1__1__36_left_grid_pin_25_;
  wire [0:0] cby_1__1__36_left_grid_pin_26_;
  wire [0:0] cby_1__1__36_left_grid_pin_27_;
  wire [0:0] cby_1__1__36_left_grid_pin_28_;
  wire [0:0] cby_1__1__36_left_grid_pin_29_;
  wire [0:0] cby_1__1__36_left_grid_pin_30_;
  wire [0:0] cby_1__1__36_left_grid_pin_31_;
  wire [0:0] cby_1__1__37_ccff_tail;
  wire [0:19] cby_1__1__37_chany_bottom_out;
  wire [0:19] cby_1__1__37_chany_top_out;
  wire [0:0] cby_1__1__37_left_grid_pin_16_;
  wire [0:0] cby_1__1__37_left_grid_pin_17_;
  wire [0:0] cby_1__1__37_left_grid_pin_18_;
  wire [0:0] cby_1__1__37_left_grid_pin_19_;
  wire [0:0] cby_1__1__37_left_grid_pin_20_;
  wire [0:0] cby_1__1__37_left_grid_pin_21_;
  wire [0:0] cby_1__1__37_left_grid_pin_22_;
  wire [0:0] cby_1__1__37_left_grid_pin_23_;
  wire [0:0] cby_1__1__37_left_grid_pin_24_;
  wire [0:0] cby_1__1__37_left_grid_pin_25_;
  wire [0:0] cby_1__1__37_left_grid_pin_26_;
  wire [0:0] cby_1__1__37_left_grid_pin_27_;
  wire [0:0] cby_1__1__37_left_grid_pin_28_;
  wire [0:0] cby_1__1__37_left_grid_pin_29_;
  wire [0:0] cby_1__1__37_left_grid_pin_30_;
  wire [0:0] cby_1__1__37_left_grid_pin_31_;
  wire [0:0] cby_1__1__38_ccff_tail;
  wire [0:19] cby_1__1__38_chany_bottom_out;
  wire [0:19] cby_1__1__38_chany_top_out;
  wire [0:0] cby_1__1__38_left_grid_pin_16_;
  wire [0:0] cby_1__1__38_left_grid_pin_17_;
  wire [0:0] cby_1__1__38_left_grid_pin_18_;
  wire [0:0] cby_1__1__38_left_grid_pin_19_;
  wire [0:0] cby_1__1__38_left_grid_pin_20_;
  wire [0:0] cby_1__1__38_left_grid_pin_21_;
  wire [0:0] cby_1__1__38_left_grid_pin_22_;
  wire [0:0] cby_1__1__38_left_grid_pin_23_;
  wire [0:0] cby_1__1__38_left_grid_pin_24_;
  wire [0:0] cby_1__1__38_left_grid_pin_25_;
  wire [0:0] cby_1__1__38_left_grid_pin_26_;
  wire [0:0] cby_1__1__38_left_grid_pin_27_;
  wire [0:0] cby_1__1__38_left_grid_pin_28_;
  wire [0:0] cby_1__1__38_left_grid_pin_29_;
  wire [0:0] cby_1__1__38_left_grid_pin_30_;
  wire [0:0] cby_1__1__38_left_grid_pin_31_;
  wire [0:0] cby_1__1__39_ccff_tail;
  wire [0:19] cby_1__1__39_chany_bottom_out;
  wire [0:19] cby_1__1__39_chany_top_out;
  wire [0:0] cby_1__1__39_left_grid_pin_16_;
  wire [0:0] cby_1__1__39_left_grid_pin_17_;
  wire [0:0] cby_1__1__39_left_grid_pin_18_;
  wire [0:0] cby_1__1__39_left_grid_pin_19_;
  wire [0:0] cby_1__1__39_left_grid_pin_20_;
  wire [0:0] cby_1__1__39_left_grid_pin_21_;
  wire [0:0] cby_1__1__39_left_grid_pin_22_;
  wire [0:0] cby_1__1__39_left_grid_pin_23_;
  wire [0:0] cby_1__1__39_left_grid_pin_24_;
  wire [0:0] cby_1__1__39_left_grid_pin_25_;
  wire [0:0] cby_1__1__39_left_grid_pin_26_;
  wire [0:0] cby_1__1__39_left_grid_pin_27_;
  wire [0:0] cby_1__1__39_left_grid_pin_28_;
  wire [0:0] cby_1__1__39_left_grid_pin_29_;
  wire [0:0] cby_1__1__39_left_grid_pin_30_;
  wire [0:0] cby_1__1__39_left_grid_pin_31_;
  wire [0:0] cby_1__1__3_ccff_tail;
  wire [0:19] cby_1__1__3_chany_bottom_out;
  wire [0:19] cby_1__1__3_chany_top_out;
  wire [0:0] cby_1__1__3_left_grid_pin_16_;
  wire [0:0] cby_1__1__3_left_grid_pin_17_;
  wire [0:0] cby_1__1__3_left_grid_pin_18_;
  wire [0:0] cby_1__1__3_left_grid_pin_19_;
  wire [0:0] cby_1__1__3_left_grid_pin_20_;
  wire [0:0] cby_1__1__3_left_grid_pin_21_;
  wire [0:0] cby_1__1__3_left_grid_pin_22_;
  wire [0:0] cby_1__1__3_left_grid_pin_23_;
  wire [0:0] cby_1__1__3_left_grid_pin_24_;
  wire [0:0] cby_1__1__3_left_grid_pin_25_;
  wire [0:0] cby_1__1__3_left_grid_pin_26_;
  wire [0:0] cby_1__1__3_left_grid_pin_27_;
  wire [0:0] cby_1__1__3_left_grid_pin_28_;
  wire [0:0] cby_1__1__3_left_grid_pin_29_;
  wire [0:0] cby_1__1__3_left_grid_pin_30_;
  wire [0:0] cby_1__1__3_left_grid_pin_31_;
  wire [0:0] cby_1__1__40_ccff_tail;
  wire [0:19] cby_1__1__40_chany_bottom_out;
  wire [0:19] cby_1__1__40_chany_top_out;
  wire [0:0] cby_1__1__40_left_grid_pin_16_;
  wire [0:0] cby_1__1__40_left_grid_pin_17_;
  wire [0:0] cby_1__1__40_left_grid_pin_18_;
  wire [0:0] cby_1__1__40_left_grid_pin_19_;
  wire [0:0] cby_1__1__40_left_grid_pin_20_;
  wire [0:0] cby_1__1__40_left_grid_pin_21_;
  wire [0:0] cby_1__1__40_left_grid_pin_22_;
  wire [0:0] cby_1__1__40_left_grid_pin_23_;
  wire [0:0] cby_1__1__40_left_grid_pin_24_;
  wire [0:0] cby_1__1__40_left_grid_pin_25_;
  wire [0:0] cby_1__1__40_left_grid_pin_26_;
  wire [0:0] cby_1__1__40_left_grid_pin_27_;
  wire [0:0] cby_1__1__40_left_grid_pin_28_;
  wire [0:0] cby_1__1__40_left_grid_pin_29_;
  wire [0:0] cby_1__1__40_left_grid_pin_30_;
  wire [0:0] cby_1__1__40_left_grid_pin_31_;
  wire [0:0] cby_1__1__41_ccff_tail;
  wire [0:19] cby_1__1__41_chany_bottom_out;
  wire [0:19] cby_1__1__41_chany_top_out;
  wire [0:0] cby_1__1__41_left_grid_pin_16_;
  wire [0:0] cby_1__1__41_left_grid_pin_17_;
  wire [0:0] cby_1__1__41_left_grid_pin_18_;
  wire [0:0] cby_1__1__41_left_grid_pin_19_;
  wire [0:0] cby_1__1__41_left_grid_pin_20_;
  wire [0:0] cby_1__1__41_left_grid_pin_21_;
  wire [0:0] cby_1__1__41_left_grid_pin_22_;
  wire [0:0] cby_1__1__41_left_grid_pin_23_;
  wire [0:0] cby_1__1__41_left_grid_pin_24_;
  wire [0:0] cby_1__1__41_left_grid_pin_25_;
  wire [0:0] cby_1__1__41_left_grid_pin_26_;
  wire [0:0] cby_1__1__41_left_grid_pin_27_;
  wire [0:0] cby_1__1__41_left_grid_pin_28_;
  wire [0:0] cby_1__1__41_left_grid_pin_29_;
  wire [0:0] cby_1__1__41_left_grid_pin_30_;
  wire [0:0] cby_1__1__41_left_grid_pin_31_;
  wire [0:0] cby_1__1__42_ccff_tail;
  wire [0:19] cby_1__1__42_chany_bottom_out;
  wire [0:19] cby_1__1__42_chany_top_out;
  wire [0:0] cby_1__1__42_left_grid_pin_16_;
  wire [0:0] cby_1__1__42_left_grid_pin_17_;
  wire [0:0] cby_1__1__42_left_grid_pin_18_;
  wire [0:0] cby_1__1__42_left_grid_pin_19_;
  wire [0:0] cby_1__1__42_left_grid_pin_20_;
  wire [0:0] cby_1__1__42_left_grid_pin_21_;
  wire [0:0] cby_1__1__42_left_grid_pin_22_;
  wire [0:0] cby_1__1__42_left_grid_pin_23_;
  wire [0:0] cby_1__1__42_left_grid_pin_24_;
  wire [0:0] cby_1__1__42_left_grid_pin_25_;
  wire [0:0] cby_1__1__42_left_grid_pin_26_;
  wire [0:0] cby_1__1__42_left_grid_pin_27_;
  wire [0:0] cby_1__1__42_left_grid_pin_28_;
  wire [0:0] cby_1__1__42_left_grid_pin_29_;
  wire [0:0] cby_1__1__42_left_grid_pin_30_;
  wire [0:0] cby_1__1__42_left_grid_pin_31_;
  wire [0:0] cby_1__1__43_ccff_tail;
  wire [0:19] cby_1__1__43_chany_bottom_out;
  wire [0:19] cby_1__1__43_chany_top_out;
  wire [0:0] cby_1__1__43_left_grid_pin_16_;
  wire [0:0] cby_1__1__43_left_grid_pin_17_;
  wire [0:0] cby_1__1__43_left_grid_pin_18_;
  wire [0:0] cby_1__1__43_left_grid_pin_19_;
  wire [0:0] cby_1__1__43_left_grid_pin_20_;
  wire [0:0] cby_1__1__43_left_grid_pin_21_;
  wire [0:0] cby_1__1__43_left_grid_pin_22_;
  wire [0:0] cby_1__1__43_left_grid_pin_23_;
  wire [0:0] cby_1__1__43_left_grid_pin_24_;
  wire [0:0] cby_1__1__43_left_grid_pin_25_;
  wire [0:0] cby_1__1__43_left_grid_pin_26_;
  wire [0:0] cby_1__1__43_left_grid_pin_27_;
  wire [0:0] cby_1__1__43_left_grid_pin_28_;
  wire [0:0] cby_1__1__43_left_grid_pin_29_;
  wire [0:0] cby_1__1__43_left_grid_pin_30_;
  wire [0:0] cby_1__1__43_left_grid_pin_31_;
  wire [0:0] cby_1__1__44_ccff_tail;
  wire [0:19] cby_1__1__44_chany_bottom_out;
  wire [0:19] cby_1__1__44_chany_top_out;
  wire [0:0] cby_1__1__44_left_grid_pin_16_;
  wire [0:0] cby_1__1__44_left_grid_pin_17_;
  wire [0:0] cby_1__1__44_left_grid_pin_18_;
  wire [0:0] cby_1__1__44_left_grid_pin_19_;
  wire [0:0] cby_1__1__44_left_grid_pin_20_;
  wire [0:0] cby_1__1__44_left_grid_pin_21_;
  wire [0:0] cby_1__1__44_left_grid_pin_22_;
  wire [0:0] cby_1__1__44_left_grid_pin_23_;
  wire [0:0] cby_1__1__44_left_grid_pin_24_;
  wire [0:0] cby_1__1__44_left_grid_pin_25_;
  wire [0:0] cby_1__1__44_left_grid_pin_26_;
  wire [0:0] cby_1__1__44_left_grid_pin_27_;
  wire [0:0] cby_1__1__44_left_grid_pin_28_;
  wire [0:0] cby_1__1__44_left_grid_pin_29_;
  wire [0:0] cby_1__1__44_left_grid_pin_30_;
  wire [0:0] cby_1__1__44_left_grid_pin_31_;
  wire [0:0] cby_1__1__45_ccff_tail;
  wire [0:19] cby_1__1__45_chany_bottom_out;
  wire [0:19] cby_1__1__45_chany_top_out;
  wire [0:0] cby_1__1__45_left_grid_pin_16_;
  wire [0:0] cby_1__1__45_left_grid_pin_17_;
  wire [0:0] cby_1__1__45_left_grid_pin_18_;
  wire [0:0] cby_1__1__45_left_grid_pin_19_;
  wire [0:0] cby_1__1__45_left_grid_pin_20_;
  wire [0:0] cby_1__1__45_left_grid_pin_21_;
  wire [0:0] cby_1__1__45_left_grid_pin_22_;
  wire [0:0] cby_1__1__45_left_grid_pin_23_;
  wire [0:0] cby_1__1__45_left_grid_pin_24_;
  wire [0:0] cby_1__1__45_left_grid_pin_25_;
  wire [0:0] cby_1__1__45_left_grid_pin_26_;
  wire [0:0] cby_1__1__45_left_grid_pin_27_;
  wire [0:0] cby_1__1__45_left_grid_pin_28_;
  wire [0:0] cby_1__1__45_left_grid_pin_29_;
  wire [0:0] cby_1__1__45_left_grid_pin_30_;
  wire [0:0] cby_1__1__45_left_grid_pin_31_;
  wire [0:0] cby_1__1__46_ccff_tail;
  wire [0:19] cby_1__1__46_chany_bottom_out;
  wire [0:19] cby_1__1__46_chany_top_out;
  wire [0:0] cby_1__1__46_left_grid_pin_16_;
  wire [0:0] cby_1__1__46_left_grid_pin_17_;
  wire [0:0] cby_1__1__46_left_grid_pin_18_;
  wire [0:0] cby_1__1__46_left_grid_pin_19_;
  wire [0:0] cby_1__1__46_left_grid_pin_20_;
  wire [0:0] cby_1__1__46_left_grid_pin_21_;
  wire [0:0] cby_1__1__46_left_grid_pin_22_;
  wire [0:0] cby_1__1__46_left_grid_pin_23_;
  wire [0:0] cby_1__1__46_left_grid_pin_24_;
  wire [0:0] cby_1__1__46_left_grid_pin_25_;
  wire [0:0] cby_1__1__46_left_grid_pin_26_;
  wire [0:0] cby_1__1__46_left_grid_pin_27_;
  wire [0:0] cby_1__1__46_left_grid_pin_28_;
  wire [0:0] cby_1__1__46_left_grid_pin_29_;
  wire [0:0] cby_1__1__46_left_grid_pin_30_;
  wire [0:0] cby_1__1__46_left_grid_pin_31_;
  wire [0:0] cby_1__1__47_ccff_tail;
  wire [0:19] cby_1__1__47_chany_bottom_out;
  wire [0:19] cby_1__1__47_chany_top_out;
  wire [0:0] cby_1__1__47_left_grid_pin_16_;
  wire [0:0] cby_1__1__47_left_grid_pin_17_;
  wire [0:0] cby_1__1__47_left_grid_pin_18_;
  wire [0:0] cby_1__1__47_left_grid_pin_19_;
  wire [0:0] cby_1__1__47_left_grid_pin_20_;
  wire [0:0] cby_1__1__47_left_grid_pin_21_;
  wire [0:0] cby_1__1__47_left_grid_pin_22_;
  wire [0:0] cby_1__1__47_left_grid_pin_23_;
  wire [0:0] cby_1__1__47_left_grid_pin_24_;
  wire [0:0] cby_1__1__47_left_grid_pin_25_;
  wire [0:0] cby_1__1__47_left_grid_pin_26_;
  wire [0:0] cby_1__1__47_left_grid_pin_27_;
  wire [0:0] cby_1__1__47_left_grid_pin_28_;
  wire [0:0] cby_1__1__47_left_grid_pin_29_;
  wire [0:0] cby_1__1__47_left_grid_pin_30_;
  wire [0:0] cby_1__1__47_left_grid_pin_31_;
  wire [0:0] cby_1__1__48_ccff_tail;
  wire [0:19] cby_1__1__48_chany_bottom_out;
  wire [0:19] cby_1__1__48_chany_top_out;
  wire [0:0] cby_1__1__48_left_grid_pin_16_;
  wire [0:0] cby_1__1__48_left_grid_pin_17_;
  wire [0:0] cby_1__1__48_left_grid_pin_18_;
  wire [0:0] cby_1__1__48_left_grid_pin_19_;
  wire [0:0] cby_1__1__48_left_grid_pin_20_;
  wire [0:0] cby_1__1__48_left_grid_pin_21_;
  wire [0:0] cby_1__1__48_left_grid_pin_22_;
  wire [0:0] cby_1__1__48_left_grid_pin_23_;
  wire [0:0] cby_1__1__48_left_grid_pin_24_;
  wire [0:0] cby_1__1__48_left_grid_pin_25_;
  wire [0:0] cby_1__1__48_left_grid_pin_26_;
  wire [0:0] cby_1__1__48_left_grid_pin_27_;
  wire [0:0] cby_1__1__48_left_grid_pin_28_;
  wire [0:0] cby_1__1__48_left_grid_pin_29_;
  wire [0:0] cby_1__1__48_left_grid_pin_30_;
  wire [0:0] cby_1__1__48_left_grid_pin_31_;
  wire [0:0] cby_1__1__49_ccff_tail;
  wire [0:19] cby_1__1__49_chany_bottom_out;
  wire [0:19] cby_1__1__49_chany_top_out;
  wire [0:0] cby_1__1__49_left_grid_pin_16_;
  wire [0:0] cby_1__1__49_left_grid_pin_17_;
  wire [0:0] cby_1__1__49_left_grid_pin_18_;
  wire [0:0] cby_1__1__49_left_grid_pin_19_;
  wire [0:0] cby_1__1__49_left_grid_pin_20_;
  wire [0:0] cby_1__1__49_left_grid_pin_21_;
  wire [0:0] cby_1__1__49_left_grid_pin_22_;
  wire [0:0] cby_1__1__49_left_grid_pin_23_;
  wire [0:0] cby_1__1__49_left_grid_pin_24_;
  wire [0:0] cby_1__1__49_left_grid_pin_25_;
  wire [0:0] cby_1__1__49_left_grid_pin_26_;
  wire [0:0] cby_1__1__49_left_grid_pin_27_;
  wire [0:0] cby_1__1__49_left_grid_pin_28_;
  wire [0:0] cby_1__1__49_left_grid_pin_29_;
  wire [0:0] cby_1__1__49_left_grid_pin_30_;
  wire [0:0] cby_1__1__49_left_grid_pin_31_;
  wire [0:0] cby_1__1__4_ccff_tail;
  wire [0:19] cby_1__1__4_chany_bottom_out;
  wire [0:19] cby_1__1__4_chany_top_out;
  wire [0:0] cby_1__1__4_left_grid_pin_16_;
  wire [0:0] cby_1__1__4_left_grid_pin_17_;
  wire [0:0] cby_1__1__4_left_grid_pin_18_;
  wire [0:0] cby_1__1__4_left_grid_pin_19_;
  wire [0:0] cby_1__1__4_left_grid_pin_20_;
  wire [0:0] cby_1__1__4_left_grid_pin_21_;
  wire [0:0] cby_1__1__4_left_grid_pin_22_;
  wire [0:0] cby_1__1__4_left_grid_pin_23_;
  wire [0:0] cby_1__1__4_left_grid_pin_24_;
  wire [0:0] cby_1__1__4_left_grid_pin_25_;
  wire [0:0] cby_1__1__4_left_grid_pin_26_;
  wire [0:0] cby_1__1__4_left_grid_pin_27_;
  wire [0:0] cby_1__1__4_left_grid_pin_28_;
  wire [0:0] cby_1__1__4_left_grid_pin_29_;
  wire [0:0] cby_1__1__4_left_grid_pin_30_;
  wire [0:0] cby_1__1__4_left_grid_pin_31_;
  wire [0:0] cby_1__1__50_ccff_tail;
  wire [0:19] cby_1__1__50_chany_bottom_out;
  wire [0:19] cby_1__1__50_chany_top_out;
  wire [0:0] cby_1__1__50_left_grid_pin_16_;
  wire [0:0] cby_1__1__50_left_grid_pin_17_;
  wire [0:0] cby_1__1__50_left_grid_pin_18_;
  wire [0:0] cby_1__1__50_left_grid_pin_19_;
  wire [0:0] cby_1__1__50_left_grid_pin_20_;
  wire [0:0] cby_1__1__50_left_grid_pin_21_;
  wire [0:0] cby_1__1__50_left_grid_pin_22_;
  wire [0:0] cby_1__1__50_left_grid_pin_23_;
  wire [0:0] cby_1__1__50_left_grid_pin_24_;
  wire [0:0] cby_1__1__50_left_grid_pin_25_;
  wire [0:0] cby_1__1__50_left_grid_pin_26_;
  wire [0:0] cby_1__1__50_left_grid_pin_27_;
  wire [0:0] cby_1__1__50_left_grid_pin_28_;
  wire [0:0] cby_1__1__50_left_grid_pin_29_;
  wire [0:0] cby_1__1__50_left_grid_pin_30_;
  wire [0:0] cby_1__1__50_left_grid_pin_31_;
  wire [0:0] cby_1__1__51_ccff_tail;
  wire [0:19] cby_1__1__51_chany_bottom_out;
  wire [0:19] cby_1__1__51_chany_top_out;
  wire [0:0] cby_1__1__51_left_grid_pin_16_;
  wire [0:0] cby_1__1__51_left_grid_pin_17_;
  wire [0:0] cby_1__1__51_left_grid_pin_18_;
  wire [0:0] cby_1__1__51_left_grid_pin_19_;
  wire [0:0] cby_1__1__51_left_grid_pin_20_;
  wire [0:0] cby_1__1__51_left_grid_pin_21_;
  wire [0:0] cby_1__1__51_left_grid_pin_22_;
  wire [0:0] cby_1__1__51_left_grid_pin_23_;
  wire [0:0] cby_1__1__51_left_grid_pin_24_;
  wire [0:0] cby_1__1__51_left_grid_pin_25_;
  wire [0:0] cby_1__1__51_left_grid_pin_26_;
  wire [0:0] cby_1__1__51_left_grid_pin_27_;
  wire [0:0] cby_1__1__51_left_grid_pin_28_;
  wire [0:0] cby_1__1__51_left_grid_pin_29_;
  wire [0:0] cby_1__1__51_left_grid_pin_30_;
  wire [0:0] cby_1__1__51_left_grid_pin_31_;
  wire [0:0] cby_1__1__52_ccff_tail;
  wire [0:19] cby_1__1__52_chany_bottom_out;
  wire [0:19] cby_1__1__52_chany_top_out;
  wire [0:0] cby_1__1__52_left_grid_pin_16_;
  wire [0:0] cby_1__1__52_left_grid_pin_17_;
  wire [0:0] cby_1__1__52_left_grid_pin_18_;
  wire [0:0] cby_1__1__52_left_grid_pin_19_;
  wire [0:0] cby_1__1__52_left_grid_pin_20_;
  wire [0:0] cby_1__1__52_left_grid_pin_21_;
  wire [0:0] cby_1__1__52_left_grid_pin_22_;
  wire [0:0] cby_1__1__52_left_grid_pin_23_;
  wire [0:0] cby_1__1__52_left_grid_pin_24_;
  wire [0:0] cby_1__1__52_left_grid_pin_25_;
  wire [0:0] cby_1__1__52_left_grid_pin_26_;
  wire [0:0] cby_1__1__52_left_grid_pin_27_;
  wire [0:0] cby_1__1__52_left_grid_pin_28_;
  wire [0:0] cby_1__1__52_left_grid_pin_29_;
  wire [0:0] cby_1__1__52_left_grid_pin_30_;
  wire [0:0] cby_1__1__52_left_grid_pin_31_;
  wire [0:0] cby_1__1__53_ccff_tail;
  wire [0:19] cby_1__1__53_chany_bottom_out;
  wire [0:19] cby_1__1__53_chany_top_out;
  wire [0:0] cby_1__1__53_left_grid_pin_16_;
  wire [0:0] cby_1__1__53_left_grid_pin_17_;
  wire [0:0] cby_1__1__53_left_grid_pin_18_;
  wire [0:0] cby_1__1__53_left_grid_pin_19_;
  wire [0:0] cby_1__1__53_left_grid_pin_20_;
  wire [0:0] cby_1__1__53_left_grid_pin_21_;
  wire [0:0] cby_1__1__53_left_grid_pin_22_;
  wire [0:0] cby_1__1__53_left_grid_pin_23_;
  wire [0:0] cby_1__1__53_left_grid_pin_24_;
  wire [0:0] cby_1__1__53_left_grid_pin_25_;
  wire [0:0] cby_1__1__53_left_grid_pin_26_;
  wire [0:0] cby_1__1__53_left_grid_pin_27_;
  wire [0:0] cby_1__1__53_left_grid_pin_28_;
  wire [0:0] cby_1__1__53_left_grid_pin_29_;
  wire [0:0] cby_1__1__53_left_grid_pin_30_;
  wire [0:0] cby_1__1__53_left_grid_pin_31_;
  wire [0:0] cby_1__1__54_ccff_tail;
  wire [0:19] cby_1__1__54_chany_bottom_out;
  wire [0:19] cby_1__1__54_chany_top_out;
  wire [0:0] cby_1__1__54_left_grid_pin_16_;
  wire [0:0] cby_1__1__54_left_grid_pin_17_;
  wire [0:0] cby_1__1__54_left_grid_pin_18_;
  wire [0:0] cby_1__1__54_left_grid_pin_19_;
  wire [0:0] cby_1__1__54_left_grid_pin_20_;
  wire [0:0] cby_1__1__54_left_grid_pin_21_;
  wire [0:0] cby_1__1__54_left_grid_pin_22_;
  wire [0:0] cby_1__1__54_left_grid_pin_23_;
  wire [0:0] cby_1__1__54_left_grid_pin_24_;
  wire [0:0] cby_1__1__54_left_grid_pin_25_;
  wire [0:0] cby_1__1__54_left_grid_pin_26_;
  wire [0:0] cby_1__1__54_left_grid_pin_27_;
  wire [0:0] cby_1__1__54_left_grid_pin_28_;
  wire [0:0] cby_1__1__54_left_grid_pin_29_;
  wire [0:0] cby_1__1__54_left_grid_pin_30_;
  wire [0:0] cby_1__1__54_left_grid_pin_31_;
  wire [0:0] cby_1__1__55_ccff_tail;
  wire [0:19] cby_1__1__55_chany_bottom_out;
  wire [0:19] cby_1__1__55_chany_top_out;
  wire [0:0] cby_1__1__55_left_grid_pin_16_;
  wire [0:0] cby_1__1__55_left_grid_pin_17_;
  wire [0:0] cby_1__1__55_left_grid_pin_18_;
  wire [0:0] cby_1__1__55_left_grid_pin_19_;
  wire [0:0] cby_1__1__55_left_grid_pin_20_;
  wire [0:0] cby_1__1__55_left_grid_pin_21_;
  wire [0:0] cby_1__1__55_left_grid_pin_22_;
  wire [0:0] cby_1__1__55_left_grid_pin_23_;
  wire [0:0] cby_1__1__55_left_grid_pin_24_;
  wire [0:0] cby_1__1__55_left_grid_pin_25_;
  wire [0:0] cby_1__1__55_left_grid_pin_26_;
  wire [0:0] cby_1__1__55_left_grid_pin_27_;
  wire [0:0] cby_1__1__55_left_grid_pin_28_;
  wire [0:0] cby_1__1__55_left_grid_pin_29_;
  wire [0:0] cby_1__1__55_left_grid_pin_30_;
  wire [0:0] cby_1__1__55_left_grid_pin_31_;
  wire [0:0] cby_1__1__5_ccff_tail;
  wire [0:19] cby_1__1__5_chany_bottom_out;
  wire [0:19] cby_1__1__5_chany_top_out;
  wire [0:0] cby_1__1__5_left_grid_pin_16_;
  wire [0:0] cby_1__1__5_left_grid_pin_17_;
  wire [0:0] cby_1__1__5_left_grid_pin_18_;
  wire [0:0] cby_1__1__5_left_grid_pin_19_;
  wire [0:0] cby_1__1__5_left_grid_pin_20_;
  wire [0:0] cby_1__1__5_left_grid_pin_21_;
  wire [0:0] cby_1__1__5_left_grid_pin_22_;
  wire [0:0] cby_1__1__5_left_grid_pin_23_;
  wire [0:0] cby_1__1__5_left_grid_pin_24_;
  wire [0:0] cby_1__1__5_left_grid_pin_25_;
  wire [0:0] cby_1__1__5_left_grid_pin_26_;
  wire [0:0] cby_1__1__5_left_grid_pin_27_;
  wire [0:0] cby_1__1__5_left_grid_pin_28_;
  wire [0:0] cby_1__1__5_left_grid_pin_29_;
  wire [0:0] cby_1__1__5_left_grid_pin_30_;
  wire [0:0] cby_1__1__5_left_grid_pin_31_;
  wire [0:0] cby_1__1__6_ccff_tail;
  wire [0:19] cby_1__1__6_chany_bottom_out;
  wire [0:19] cby_1__1__6_chany_top_out;
  wire [0:0] cby_1__1__6_left_grid_pin_16_;
  wire [0:0] cby_1__1__6_left_grid_pin_17_;
  wire [0:0] cby_1__1__6_left_grid_pin_18_;
  wire [0:0] cby_1__1__6_left_grid_pin_19_;
  wire [0:0] cby_1__1__6_left_grid_pin_20_;
  wire [0:0] cby_1__1__6_left_grid_pin_21_;
  wire [0:0] cby_1__1__6_left_grid_pin_22_;
  wire [0:0] cby_1__1__6_left_grid_pin_23_;
  wire [0:0] cby_1__1__6_left_grid_pin_24_;
  wire [0:0] cby_1__1__6_left_grid_pin_25_;
  wire [0:0] cby_1__1__6_left_grid_pin_26_;
  wire [0:0] cby_1__1__6_left_grid_pin_27_;
  wire [0:0] cby_1__1__6_left_grid_pin_28_;
  wire [0:0] cby_1__1__6_left_grid_pin_29_;
  wire [0:0] cby_1__1__6_left_grid_pin_30_;
  wire [0:0] cby_1__1__6_left_grid_pin_31_;
  wire [0:0] cby_1__1__7_ccff_tail;
  wire [0:19] cby_1__1__7_chany_bottom_out;
  wire [0:19] cby_1__1__7_chany_top_out;
  wire [0:0] cby_1__1__7_left_grid_pin_16_;
  wire [0:0] cby_1__1__7_left_grid_pin_17_;
  wire [0:0] cby_1__1__7_left_grid_pin_18_;
  wire [0:0] cby_1__1__7_left_grid_pin_19_;
  wire [0:0] cby_1__1__7_left_grid_pin_20_;
  wire [0:0] cby_1__1__7_left_grid_pin_21_;
  wire [0:0] cby_1__1__7_left_grid_pin_22_;
  wire [0:0] cby_1__1__7_left_grid_pin_23_;
  wire [0:0] cby_1__1__7_left_grid_pin_24_;
  wire [0:0] cby_1__1__7_left_grid_pin_25_;
  wire [0:0] cby_1__1__7_left_grid_pin_26_;
  wire [0:0] cby_1__1__7_left_grid_pin_27_;
  wire [0:0] cby_1__1__7_left_grid_pin_28_;
  wire [0:0] cby_1__1__7_left_grid_pin_29_;
  wire [0:0] cby_1__1__7_left_grid_pin_30_;
  wire [0:0] cby_1__1__7_left_grid_pin_31_;
  wire [0:0] cby_1__1__8_ccff_tail;
  wire [0:19] cby_1__1__8_chany_bottom_out;
  wire [0:19] cby_1__1__8_chany_top_out;
  wire [0:0] cby_1__1__8_left_grid_pin_16_;
  wire [0:0] cby_1__1__8_left_grid_pin_17_;
  wire [0:0] cby_1__1__8_left_grid_pin_18_;
  wire [0:0] cby_1__1__8_left_grid_pin_19_;
  wire [0:0] cby_1__1__8_left_grid_pin_20_;
  wire [0:0] cby_1__1__8_left_grid_pin_21_;
  wire [0:0] cby_1__1__8_left_grid_pin_22_;
  wire [0:0] cby_1__1__8_left_grid_pin_23_;
  wire [0:0] cby_1__1__8_left_grid_pin_24_;
  wire [0:0] cby_1__1__8_left_grid_pin_25_;
  wire [0:0] cby_1__1__8_left_grid_pin_26_;
  wire [0:0] cby_1__1__8_left_grid_pin_27_;
  wire [0:0] cby_1__1__8_left_grid_pin_28_;
  wire [0:0] cby_1__1__8_left_grid_pin_29_;
  wire [0:0] cby_1__1__8_left_grid_pin_30_;
  wire [0:0] cby_1__1__8_left_grid_pin_31_;
  wire [0:0] cby_1__1__9_ccff_tail;
  wire [0:19] cby_1__1__9_chany_bottom_out;
  wire [0:19] cby_1__1__9_chany_top_out;
  wire [0:0] cby_1__1__9_left_grid_pin_16_;
  wire [0:0] cby_1__1__9_left_grid_pin_17_;
  wire [0:0] cby_1__1__9_left_grid_pin_18_;
  wire [0:0] cby_1__1__9_left_grid_pin_19_;
  wire [0:0] cby_1__1__9_left_grid_pin_20_;
  wire [0:0] cby_1__1__9_left_grid_pin_21_;
  wire [0:0] cby_1__1__9_left_grid_pin_22_;
  wire [0:0] cby_1__1__9_left_grid_pin_23_;
  wire [0:0] cby_1__1__9_left_grid_pin_24_;
  wire [0:0] cby_1__1__9_left_grid_pin_25_;
  wire [0:0] cby_1__1__9_left_grid_pin_26_;
  wire [0:0] cby_1__1__9_left_grid_pin_27_;
  wire [0:0] cby_1__1__9_left_grid_pin_28_;
  wire [0:0] cby_1__1__9_left_grid_pin_29_;
  wire [0:0] cby_1__1__9_left_grid_pin_30_;
  wire [0:0] cby_1__1__9_left_grid_pin_31_;
  wire [0:0] cby_8__1__0_ccff_tail;
  wire [0:19] cby_8__1__0_chany_bottom_out;
  wire [0:19] cby_8__1__0_chany_top_out;
  wire [0:0] cby_8__1__0_left_grid_pin_16_;
  wire [0:0] cby_8__1__0_left_grid_pin_17_;
  wire [0:0] cby_8__1__0_left_grid_pin_18_;
  wire [0:0] cby_8__1__0_left_grid_pin_19_;
  wire [0:0] cby_8__1__0_left_grid_pin_20_;
  wire [0:0] cby_8__1__0_left_grid_pin_21_;
  wire [0:0] cby_8__1__0_left_grid_pin_22_;
  wire [0:0] cby_8__1__0_left_grid_pin_23_;
  wire [0:0] cby_8__1__0_left_grid_pin_24_;
  wire [0:0] cby_8__1__0_left_grid_pin_25_;
  wire [0:0] cby_8__1__0_left_grid_pin_26_;
  wire [0:0] cby_8__1__0_left_grid_pin_27_;
  wire [0:0] cby_8__1__0_left_grid_pin_28_;
  wire [0:0] cby_8__1__0_left_grid_pin_29_;
  wire [0:0] cby_8__1__0_left_grid_pin_30_;
  wire [0:0] cby_8__1__0_left_grid_pin_31_;
  wire [0:0] cby_8__1__0_right_grid_pin_0_;
  wire [0:0] cby_8__1__1_ccff_tail;
  wire [0:19] cby_8__1__1_chany_bottom_out;
  wire [0:19] cby_8__1__1_chany_top_out;
  wire [0:0] cby_8__1__1_left_grid_pin_16_;
  wire [0:0] cby_8__1__1_left_grid_pin_17_;
  wire [0:0] cby_8__1__1_left_grid_pin_18_;
  wire [0:0] cby_8__1__1_left_grid_pin_19_;
  wire [0:0] cby_8__1__1_left_grid_pin_20_;
  wire [0:0] cby_8__1__1_left_grid_pin_21_;
  wire [0:0] cby_8__1__1_left_grid_pin_22_;
  wire [0:0] cby_8__1__1_left_grid_pin_23_;
  wire [0:0] cby_8__1__1_left_grid_pin_24_;
  wire [0:0] cby_8__1__1_left_grid_pin_25_;
  wire [0:0] cby_8__1__1_left_grid_pin_26_;
  wire [0:0] cby_8__1__1_left_grid_pin_27_;
  wire [0:0] cby_8__1__1_left_grid_pin_28_;
  wire [0:0] cby_8__1__1_left_grid_pin_29_;
  wire [0:0] cby_8__1__1_left_grid_pin_30_;
  wire [0:0] cby_8__1__1_left_grid_pin_31_;
  wire [0:0] cby_8__1__1_right_grid_pin_0_;
  wire [0:0] cby_8__1__2_ccff_tail;
  wire [0:19] cby_8__1__2_chany_bottom_out;
  wire [0:19] cby_8__1__2_chany_top_out;
  wire [0:0] cby_8__1__2_left_grid_pin_16_;
  wire [0:0] cby_8__1__2_left_grid_pin_17_;
  wire [0:0] cby_8__1__2_left_grid_pin_18_;
  wire [0:0] cby_8__1__2_left_grid_pin_19_;
  wire [0:0] cby_8__1__2_left_grid_pin_20_;
  wire [0:0] cby_8__1__2_left_grid_pin_21_;
  wire [0:0] cby_8__1__2_left_grid_pin_22_;
  wire [0:0] cby_8__1__2_left_grid_pin_23_;
  wire [0:0] cby_8__1__2_left_grid_pin_24_;
  wire [0:0] cby_8__1__2_left_grid_pin_25_;
  wire [0:0] cby_8__1__2_left_grid_pin_26_;
  wire [0:0] cby_8__1__2_left_grid_pin_27_;
  wire [0:0] cby_8__1__2_left_grid_pin_28_;
  wire [0:0] cby_8__1__2_left_grid_pin_29_;
  wire [0:0] cby_8__1__2_left_grid_pin_30_;
  wire [0:0] cby_8__1__2_left_grid_pin_31_;
  wire [0:0] cby_8__1__2_right_grid_pin_0_;
  wire [0:0] cby_8__1__3_ccff_tail;
  wire [0:19] cby_8__1__3_chany_bottom_out;
  wire [0:19] cby_8__1__3_chany_top_out;
  wire [0:0] cby_8__1__3_left_grid_pin_16_;
  wire [0:0] cby_8__1__3_left_grid_pin_17_;
  wire [0:0] cby_8__1__3_left_grid_pin_18_;
  wire [0:0] cby_8__1__3_left_grid_pin_19_;
  wire [0:0] cby_8__1__3_left_grid_pin_20_;
  wire [0:0] cby_8__1__3_left_grid_pin_21_;
  wire [0:0] cby_8__1__3_left_grid_pin_22_;
  wire [0:0] cby_8__1__3_left_grid_pin_23_;
  wire [0:0] cby_8__1__3_left_grid_pin_24_;
  wire [0:0] cby_8__1__3_left_grid_pin_25_;
  wire [0:0] cby_8__1__3_left_grid_pin_26_;
  wire [0:0] cby_8__1__3_left_grid_pin_27_;
  wire [0:0] cby_8__1__3_left_grid_pin_28_;
  wire [0:0] cby_8__1__3_left_grid_pin_29_;
  wire [0:0] cby_8__1__3_left_grid_pin_30_;
  wire [0:0] cby_8__1__3_left_grid_pin_31_;
  wire [0:0] cby_8__1__3_right_grid_pin_0_;
  wire [0:0] cby_8__1__4_ccff_tail;
  wire [0:19] cby_8__1__4_chany_bottom_out;
  wire [0:19] cby_8__1__4_chany_top_out;
  wire [0:0] cby_8__1__4_left_grid_pin_16_;
  wire [0:0] cby_8__1__4_left_grid_pin_17_;
  wire [0:0] cby_8__1__4_left_grid_pin_18_;
  wire [0:0] cby_8__1__4_left_grid_pin_19_;
  wire [0:0] cby_8__1__4_left_grid_pin_20_;
  wire [0:0] cby_8__1__4_left_grid_pin_21_;
  wire [0:0] cby_8__1__4_left_grid_pin_22_;
  wire [0:0] cby_8__1__4_left_grid_pin_23_;
  wire [0:0] cby_8__1__4_left_grid_pin_24_;
  wire [0:0] cby_8__1__4_left_grid_pin_25_;
  wire [0:0] cby_8__1__4_left_grid_pin_26_;
  wire [0:0] cby_8__1__4_left_grid_pin_27_;
  wire [0:0] cby_8__1__4_left_grid_pin_28_;
  wire [0:0] cby_8__1__4_left_grid_pin_29_;
  wire [0:0] cby_8__1__4_left_grid_pin_30_;
  wire [0:0] cby_8__1__4_left_grid_pin_31_;
  wire [0:0] cby_8__1__4_right_grid_pin_0_;
  wire [0:0] cby_8__1__5_ccff_tail;
  wire [0:19] cby_8__1__5_chany_bottom_out;
  wire [0:19] cby_8__1__5_chany_top_out;
  wire [0:0] cby_8__1__5_left_grid_pin_16_;
  wire [0:0] cby_8__1__5_left_grid_pin_17_;
  wire [0:0] cby_8__1__5_left_grid_pin_18_;
  wire [0:0] cby_8__1__5_left_grid_pin_19_;
  wire [0:0] cby_8__1__5_left_grid_pin_20_;
  wire [0:0] cby_8__1__5_left_grid_pin_21_;
  wire [0:0] cby_8__1__5_left_grid_pin_22_;
  wire [0:0] cby_8__1__5_left_grid_pin_23_;
  wire [0:0] cby_8__1__5_left_grid_pin_24_;
  wire [0:0] cby_8__1__5_left_grid_pin_25_;
  wire [0:0] cby_8__1__5_left_grid_pin_26_;
  wire [0:0] cby_8__1__5_left_grid_pin_27_;
  wire [0:0] cby_8__1__5_left_grid_pin_28_;
  wire [0:0] cby_8__1__5_left_grid_pin_29_;
  wire [0:0] cby_8__1__5_left_grid_pin_30_;
  wire [0:0] cby_8__1__5_left_grid_pin_31_;
  wire [0:0] cby_8__1__5_right_grid_pin_0_;
  wire [0:0] cby_8__1__6_ccff_tail;
  wire [0:19] cby_8__1__6_chany_bottom_out;
  wire [0:19] cby_8__1__6_chany_top_out;
  wire [0:0] cby_8__1__6_left_grid_pin_16_;
  wire [0:0] cby_8__1__6_left_grid_pin_17_;
  wire [0:0] cby_8__1__6_left_grid_pin_18_;
  wire [0:0] cby_8__1__6_left_grid_pin_19_;
  wire [0:0] cby_8__1__6_left_grid_pin_20_;
  wire [0:0] cby_8__1__6_left_grid_pin_21_;
  wire [0:0] cby_8__1__6_left_grid_pin_22_;
  wire [0:0] cby_8__1__6_left_grid_pin_23_;
  wire [0:0] cby_8__1__6_left_grid_pin_24_;
  wire [0:0] cby_8__1__6_left_grid_pin_25_;
  wire [0:0] cby_8__1__6_left_grid_pin_26_;
  wire [0:0] cby_8__1__6_left_grid_pin_27_;
  wire [0:0] cby_8__1__6_left_grid_pin_28_;
  wire [0:0] cby_8__1__6_left_grid_pin_29_;
  wire [0:0] cby_8__1__6_left_grid_pin_30_;
  wire [0:0] cby_8__1__6_left_grid_pin_31_;
  wire [0:0] cby_8__1__6_right_grid_pin_0_;
  wire [0:0] cby_8__1__7_ccff_tail;
  wire [0:19] cby_8__1__7_chany_bottom_out;
  wire [0:19] cby_8__1__7_chany_top_out;
  wire [0:0] cby_8__1__7_left_grid_pin_16_;
  wire [0:0] cby_8__1__7_left_grid_pin_17_;
  wire [0:0] cby_8__1__7_left_grid_pin_18_;
  wire [0:0] cby_8__1__7_left_grid_pin_19_;
  wire [0:0] cby_8__1__7_left_grid_pin_20_;
  wire [0:0] cby_8__1__7_left_grid_pin_21_;
  wire [0:0] cby_8__1__7_left_grid_pin_22_;
  wire [0:0] cby_8__1__7_left_grid_pin_23_;
  wire [0:0] cby_8__1__7_left_grid_pin_24_;
  wire [0:0] cby_8__1__7_left_grid_pin_25_;
  wire [0:0] cby_8__1__7_left_grid_pin_26_;
  wire [0:0] cby_8__1__7_left_grid_pin_27_;
  wire [0:0] cby_8__1__7_left_grid_pin_28_;
  wire [0:0] cby_8__1__7_left_grid_pin_29_;
  wire [0:0] cby_8__1__7_left_grid_pin_30_;
  wire [0:0] cby_8__1__7_left_grid_pin_31_;
  wire [0:0] cby_8__1__7_right_grid_pin_0_;
  wire [0:0] direct_interc_0_out;
  wire [0:0] direct_interc_100_out;
  wire [0:0] direct_interc_101_out;
  wire [0:0] direct_interc_102_out;
  wire [0:0] direct_interc_103_out;
  wire [0:0] direct_interc_104_out;
  wire [0:0] direct_interc_105_out;
  wire [0:0] direct_interc_106_out;
  wire [0:0] direct_interc_107_out;
  wire [0:0] direct_interc_108_out;
  wire [0:0] direct_interc_109_out;
  wire [0:0] direct_interc_10_out;
  wire [0:0] direct_interc_110_out;
  wire [0:0] direct_interc_111_out;
  wire [0:0] direct_interc_112_out;
  wire [0:0] direct_interc_113_out;
  wire [0:0] direct_interc_114_out;
  wire [0:0] direct_interc_115_out;
  wire [0:0] direct_interc_116_out;
  wire [0:0] direct_interc_117_out;
  wire [0:0] direct_interc_118_out;
  wire [0:0] direct_interc_11_out;
  wire [0:0] direct_interc_12_out;
  wire [0:0] direct_interc_13_out;
  wire [0:0] direct_interc_14_out;
  wire [0:0] direct_interc_15_out;
  wire [0:0] direct_interc_16_out;
  wire [0:0] direct_interc_17_out;
  wire [0:0] direct_interc_18_out;
  wire [0:0] direct_interc_19_out;
  wire [0:0] direct_interc_1_out;
  wire [0:0] direct_interc_20_out;
  wire [0:0] direct_interc_21_out;
  wire [0:0] direct_interc_22_out;
  wire [0:0] direct_interc_23_out;
  wire [0:0] direct_interc_24_out;
  wire [0:0] direct_interc_25_out;
  wire [0:0] direct_interc_26_out;
  wire [0:0] direct_interc_27_out;
  wire [0:0] direct_interc_28_out;
  wire [0:0] direct_interc_29_out;
  wire [0:0] direct_interc_2_out;
  wire [0:0] direct_interc_30_out;
  wire [0:0] direct_interc_31_out;
  wire [0:0] direct_interc_32_out;
  wire [0:0] direct_interc_33_out;
  wire [0:0] direct_interc_34_out;
  wire [0:0] direct_interc_35_out;
  wire [0:0] direct_interc_36_out;
  wire [0:0] direct_interc_37_out;
  wire [0:0] direct_interc_38_out;
  wire [0:0] direct_interc_39_out;
  wire [0:0] direct_interc_3_out;
  wire [0:0] direct_interc_40_out;
  wire [0:0] direct_interc_41_out;
  wire [0:0] direct_interc_42_out;
  wire [0:0] direct_interc_43_out;
  wire [0:0] direct_interc_44_out;
  wire [0:0] direct_interc_45_out;
  wire [0:0] direct_interc_46_out;
  wire [0:0] direct_interc_47_out;
  wire [0:0] direct_interc_48_out;
  wire [0:0] direct_interc_49_out;
  wire [0:0] direct_interc_4_out;
  wire [0:0] direct_interc_50_out;
  wire [0:0] direct_interc_51_out;
  wire [0:0] direct_interc_52_out;
  wire [0:0] direct_interc_53_out;
  wire [0:0] direct_interc_54_out;
  wire [0:0] direct_interc_55_out;
  wire [0:0] direct_interc_56_out;
  wire [0:0] direct_interc_57_out;
  wire [0:0] direct_interc_58_out;
  wire [0:0] direct_interc_59_out;
  wire [0:0] direct_interc_5_out;
  wire [0:0] direct_interc_60_out;
  wire [0:0] direct_interc_61_out;
  wire [0:0] direct_interc_62_out;
  wire [0:0] direct_interc_63_out;
  wire [0:0] direct_interc_64_out;
  wire [0:0] direct_interc_65_out;
  wire [0:0] direct_interc_66_out;
  wire [0:0] direct_interc_67_out;
  wire [0:0] direct_interc_68_out;
  wire [0:0] direct_interc_69_out;
  wire [0:0] direct_interc_6_out;
  wire [0:0] direct_interc_70_out;
  wire [0:0] direct_interc_71_out;
  wire [0:0] direct_interc_72_out;
  wire [0:0] direct_interc_73_out;
  wire [0:0] direct_interc_74_out;
  wire [0:0] direct_interc_75_out;
  wire [0:0] direct_interc_76_out;
  wire [0:0] direct_interc_77_out;
  wire [0:0] direct_interc_78_out;
  wire [0:0] direct_interc_79_out;
  wire [0:0] direct_interc_7_out;
  wire [0:0] direct_interc_80_out;
  wire [0:0] direct_interc_81_out;
  wire [0:0] direct_interc_82_out;
  wire [0:0] direct_interc_83_out;
  wire [0:0] direct_interc_84_out;
  wire [0:0] direct_interc_85_out;
  wire [0:0] direct_interc_86_out;
  wire [0:0] direct_interc_87_out;
  wire [0:0] direct_interc_88_out;
  wire [0:0] direct_interc_89_out;
  wire [0:0] direct_interc_8_out;
  wire [0:0] direct_interc_90_out;
  wire [0:0] direct_interc_91_out;
  wire [0:0] direct_interc_92_out;
  wire [0:0] direct_interc_93_out;
  wire [0:0] direct_interc_94_out;
  wire [0:0] direct_interc_95_out;
  wire [0:0] direct_interc_96_out;
  wire [0:0] direct_interc_97_out;
  wire [0:0] direct_interc_98_out;
  wire [0:0] direct_interc_99_out;
  wire [0:0] direct_interc_9_out;
  wire [0:0] grid_clb_0_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_0_ccff_tail;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_0_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_0_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_10_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_10_ccff_tail;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_10_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_10_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_11_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_11_ccff_tail;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_11_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_11_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_12_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_12_ccff_tail;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_12_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_12_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_13_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_13_ccff_tail;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_13_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_13_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_14_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_14_ccff_tail;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_14_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_14_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_15_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_15_ccff_tail;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_15_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_15_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_16_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_16_ccff_tail;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_16_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_16_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_17_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_17_ccff_tail;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_17_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_17_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_18_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_18_ccff_tail;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_18_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_18_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_19_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_19_ccff_tail;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_19_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_19_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_1__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_1__8__undriven_top_width_0_height_0__pin_33_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_1_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_1_ccff_tail;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_1_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_1_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_20_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_20_ccff_tail;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_20_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_20_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_21_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_21_ccff_tail;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_21_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_21_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_22_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_22_ccff_tail;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_22_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_22_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_23_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_23_ccff_tail;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_23_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_23_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_24_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_24_ccff_tail;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_24_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_24_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_25_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_25_ccff_tail;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_25_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_25_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_26_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_26_ccff_tail;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_26_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_26_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_27_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_27_ccff_tail;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_27_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_27_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_28_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_28_ccff_tail;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_28_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_28_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_29_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_29_ccff_tail;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_29_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_29_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_2__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_2_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_2_ccff_tail;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_2_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_2_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_30_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_30_ccff_tail;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_30_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_30_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_31_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_31_ccff_tail;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_31_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_31_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_32_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_32_ccff_tail;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_32_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_32_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_33_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_33_ccff_tail;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_33_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_33_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_34_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_34_ccff_tail;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_34_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_34_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_35_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_35_ccff_tail;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_35_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_35_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_36_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_36_ccff_tail;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_36_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_36_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_37_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_37_ccff_tail;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_37_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_37_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_38_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_38_ccff_tail;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_38_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_38_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_39_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_39_ccff_tail;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_39_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_39_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_3__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_3_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_3_ccff_tail;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_3_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_3_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_40_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_40_ccff_tail;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_40_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_40_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_41_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_41_ccff_tail;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_41_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_41_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_42_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_42_ccff_tail;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_42_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_42_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_43_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_43_ccff_tail;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_43_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_43_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_44_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_44_ccff_tail;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_44_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_44_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_45_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_45_ccff_tail;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_45_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_45_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_46_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_46_ccff_tail;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_46_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_46_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_47_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_47_ccff_tail;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_47_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_47_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_48_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_48_ccff_tail;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_48_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_48_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_49_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_49_ccff_tail;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_49_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_49_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_4__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_4_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_4_ccff_tail;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_4_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_4_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_50_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_50_ccff_tail;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_50_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_50_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_51_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_51_ccff_tail;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_51_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_51_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_52_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_52_ccff_tail;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_52_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_52_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_53_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_53_ccff_tail;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_53_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_53_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_54_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_54_ccff_tail;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_54_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_54_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_55_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_55_ccff_tail;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_55_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_55_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_56_ccff_tail;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_56_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_56_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_57_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_57_ccff_tail;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_57_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_57_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_58_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_58_ccff_tail;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_58_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_58_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_59_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_59_ccff_tail;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_59_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_59_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_5__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_5__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_5_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_5_ccff_tail;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_5_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_5_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_60_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_60_ccff_tail;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_60_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_60_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_61_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_61_ccff_tail;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_61_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_61_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_62_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_62_ccff_tail;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_62_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_62_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_63_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_63_ccff_tail;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_63_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_63_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_6__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_6__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_6_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_6_ccff_tail;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_6_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_6_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_7__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_7__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_7_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_7_ccff_tail;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_7_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_7_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_8__1__undriven_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_8__8__undriven_top_width_0_height_0__pin_32_;
  wire [0:0] grid_clb_8_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_8_ccff_tail;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_8_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_8_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_50_;
  wire [0:0] grid_clb_9_bottom_width_0_height_0__pin_51_;
  wire [0:0] grid_clb_9_ccff_tail;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_42_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_42_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_43_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_43_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_44_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_45_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_46_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_47_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_48_upper;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_lower;
  wire [0:0] grid_clb_9_right_width_0_height_0__pin_49_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_34_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_34_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_35_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_35_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_36_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_37_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_38_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_39_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_40_upper;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_lower;
  wire [0:0] grid_clb_9_top_width_0_height_0__pin_41_upper;
  wire [0:0] grid_io_bottom_0_ccff_tail;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_0_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_1_ccff_tail;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_1_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_2_ccff_tail;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_2_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_3_ccff_tail;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_3_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_4_ccff_tail;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_4_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_5_ccff_tail;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_5_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_6_ccff_tail;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_6_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_bottom_7_ccff_tail;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_11_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_11_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_13_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_13_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_15_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_15_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_17_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_17_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_3_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_3_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_5_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_5_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_7_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_7_upper;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_9_lower;
  wire [0:0] grid_io_bottom_7_top_width_0_height_0__pin_9_upper;
  wire [0:0] grid_io_left_0_ccff_tail;
  wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_0_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_1_ccff_tail;
  wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_1_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_2_ccff_tail;
  wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_2_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_3_ccff_tail;
  wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_3_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_4_ccff_tail;
  wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_4_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_5_ccff_tail;
  wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_5_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_6_ccff_tail;
  wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_6_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_left_7_ccff_tail;
  wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_left_7_right_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_0_ccff_tail;
  wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_0_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_1_ccff_tail;
  wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_1_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_2_ccff_tail;
  wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_2_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_3_ccff_tail;
  wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_3_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_4_ccff_tail;
  wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_4_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_5_ccff_tail;
  wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_5_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_6_ccff_tail;
  wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_6_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_right_7_ccff_tail;
  wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_right_7_left_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_0_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_0_ccff_tail;
  wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_1_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_1_ccff_tail;
  wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_2_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_2_ccff_tail;
  wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_3_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_3_ccff_tail;
  wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_4_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_4_ccff_tail;
  wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_5_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_5_ccff_tail;
  wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_6_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_6_ccff_tail;
  wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_lower;
  wire [0:0] grid_io_top_7_bottom_width_0_height_0__pin_1_upper;
  wire [0:0] grid_io_top_7_ccff_tail;
  wire [0:19] sb_0__0__0_chanx_right_out;
  wire [0:19] sb_0__0__0_chany_top_out;
  wire [0:0] sb_0__1__0_ccff_tail;
  wire [0:19] sb_0__1__0_chanx_right_out;
  wire [0:19] sb_0__1__0_chany_bottom_out;
  wire [0:19] sb_0__1__0_chany_top_out;
  wire [0:0] sb_0__1__1_ccff_tail;
  wire [0:19] sb_0__1__1_chanx_right_out;
  wire [0:19] sb_0__1__1_chany_bottom_out;
  wire [0:19] sb_0__1__1_chany_top_out;
  wire [0:0] sb_0__1__2_ccff_tail;
  wire [0:19] sb_0__1__2_chanx_right_out;
  wire [0:19] sb_0__1__2_chany_bottom_out;
  wire [0:19] sb_0__1__2_chany_top_out;
  wire [0:0] sb_0__1__3_ccff_tail;
  wire [0:19] sb_0__1__3_chanx_right_out;
  wire [0:19] sb_0__1__3_chany_bottom_out;
  wire [0:19] sb_0__1__3_chany_top_out;
  wire [0:0] sb_0__1__4_ccff_tail;
  wire [0:19] sb_0__1__4_chanx_right_out;
  wire [0:19] sb_0__1__4_chany_bottom_out;
  wire [0:19] sb_0__1__4_chany_top_out;
  wire [0:0] sb_0__1__5_ccff_tail;
  wire [0:19] sb_0__1__5_chanx_right_out;
  wire [0:19] sb_0__1__5_chany_bottom_out;
  wire [0:19] sb_0__1__5_chany_top_out;
  wire [0:0] sb_0__1__6_ccff_tail;
  wire [0:19] sb_0__1__6_chanx_right_out;
  wire [0:19] sb_0__1__6_chany_bottom_out;
  wire [0:19] sb_0__1__6_chany_top_out;
  wire [0:0] sb_0__8__0_ccff_tail;
  wire [0:19] sb_0__8__0_chanx_right_out;
  wire [0:19] sb_0__8__0_chany_bottom_out;
  wire [0:0] sb_1__0__0_ccff_tail;
  wire [0:19] sb_1__0__0_chanx_left_out;
  wire [0:19] sb_1__0__0_chanx_right_out;
  wire [0:19] sb_1__0__0_chany_top_out;
  wire [0:0] sb_1__0__1_ccff_tail;
  wire [0:19] sb_1__0__1_chanx_left_out;
  wire [0:19] sb_1__0__1_chanx_right_out;
  wire [0:19] sb_1__0__1_chany_top_out;
  wire [0:0] sb_1__0__2_ccff_tail;
  wire [0:19] sb_1__0__2_chanx_left_out;
  wire [0:19] sb_1__0__2_chanx_right_out;
  wire [0:19] sb_1__0__2_chany_top_out;
  wire [0:0] sb_1__0__3_ccff_tail;
  wire [0:19] sb_1__0__3_chanx_left_out;
  wire [0:19] sb_1__0__3_chanx_right_out;
  wire [0:19] sb_1__0__3_chany_top_out;
  wire [0:0] sb_1__0__4_ccff_tail;
  wire [0:19] sb_1__0__4_chanx_left_out;
  wire [0:19] sb_1__0__4_chanx_right_out;
  wire [0:19] sb_1__0__4_chany_top_out;
  wire [0:0] sb_1__0__5_ccff_tail;
  wire [0:19] sb_1__0__5_chanx_left_out;
  wire [0:19] sb_1__0__5_chanx_right_out;
  wire [0:19] sb_1__0__5_chany_top_out;
  wire [0:0] sb_1__0__6_ccff_tail;
  wire [0:19] sb_1__0__6_chanx_left_out;
  wire [0:19] sb_1__0__6_chanx_right_out;
  wire [0:19] sb_1__0__6_chany_top_out;
  wire [0:0] sb_1__1__0_ccff_tail;
  wire [0:19] sb_1__1__0_chanx_left_out;
  wire [0:19] sb_1__1__0_chanx_right_out;
  wire [0:19] sb_1__1__0_chany_bottom_out;
  wire [0:19] sb_1__1__0_chany_top_out;
  wire [0:0] sb_1__1__10_ccff_tail;
  wire [0:19] sb_1__1__10_chanx_left_out;
  wire [0:19] sb_1__1__10_chanx_right_out;
  wire [0:19] sb_1__1__10_chany_bottom_out;
  wire [0:19] sb_1__1__10_chany_top_out;
  wire [0:0] sb_1__1__11_ccff_tail;
  wire [0:19] sb_1__1__11_chanx_left_out;
  wire [0:19] sb_1__1__11_chanx_right_out;
  wire [0:19] sb_1__1__11_chany_bottom_out;
  wire [0:19] sb_1__1__11_chany_top_out;
  wire [0:0] sb_1__1__12_ccff_tail;
  wire [0:19] sb_1__1__12_chanx_left_out;
  wire [0:19] sb_1__1__12_chanx_right_out;
  wire [0:19] sb_1__1__12_chany_bottom_out;
  wire [0:19] sb_1__1__12_chany_top_out;
  wire [0:0] sb_1__1__13_ccff_tail;
  wire [0:19] sb_1__1__13_chanx_left_out;
  wire [0:19] sb_1__1__13_chanx_right_out;
  wire [0:19] sb_1__1__13_chany_bottom_out;
  wire [0:19] sb_1__1__13_chany_top_out;
  wire [0:0] sb_1__1__14_ccff_tail;
  wire [0:19] sb_1__1__14_chanx_left_out;
  wire [0:19] sb_1__1__14_chanx_right_out;
  wire [0:19] sb_1__1__14_chany_bottom_out;
  wire [0:19] sb_1__1__14_chany_top_out;
  wire [0:0] sb_1__1__15_ccff_tail;
  wire [0:19] sb_1__1__15_chanx_left_out;
  wire [0:19] sb_1__1__15_chanx_right_out;
  wire [0:19] sb_1__1__15_chany_bottom_out;
  wire [0:19] sb_1__1__15_chany_top_out;
  wire [0:0] sb_1__1__16_ccff_tail;
  wire [0:19] sb_1__1__16_chanx_left_out;
  wire [0:19] sb_1__1__16_chanx_right_out;
  wire [0:19] sb_1__1__16_chany_bottom_out;
  wire [0:19] sb_1__1__16_chany_top_out;
  wire [0:0] sb_1__1__17_ccff_tail;
  wire [0:19] sb_1__1__17_chanx_left_out;
  wire [0:19] sb_1__1__17_chanx_right_out;
  wire [0:19] sb_1__1__17_chany_bottom_out;
  wire [0:19] sb_1__1__17_chany_top_out;
  wire [0:0] sb_1__1__18_ccff_tail;
  wire [0:19] sb_1__1__18_chanx_left_out;
  wire [0:19] sb_1__1__18_chanx_right_out;
  wire [0:19] sb_1__1__18_chany_bottom_out;
  wire [0:19] sb_1__1__18_chany_top_out;
  wire [0:0] sb_1__1__19_ccff_tail;
  wire [0:19] sb_1__1__19_chanx_left_out;
  wire [0:19] sb_1__1__19_chanx_right_out;
  wire [0:19] sb_1__1__19_chany_bottom_out;
  wire [0:19] sb_1__1__19_chany_top_out;
  wire [0:0] sb_1__1__1_ccff_tail;
  wire [0:19] sb_1__1__1_chanx_left_out;
  wire [0:19] sb_1__1__1_chanx_right_out;
  wire [0:19] sb_1__1__1_chany_bottom_out;
  wire [0:19] sb_1__1__1_chany_top_out;
  wire [0:0] sb_1__1__20_ccff_tail;
  wire [0:19] sb_1__1__20_chanx_left_out;
  wire [0:19] sb_1__1__20_chanx_right_out;
  wire [0:19] sb_1__1__20_chany_bottom_out;
  wire [0:19] sb_1__1__20_chany_top_out;
  wire [0:0] sb_1__1__21_ccff_tail;
  wire [0:19] sb_1__1__21_chanx_left_out;
  wire [0:19] sb_1__1__21_chanx_right_out;
  wire [0:19] sb_1__1__21_chany_bottom_out;
  wire [0:19] sb_1__1__21_chany_top_out;
  wire [0:0] sb_1__1__22_ccff_tail;
  wire [0:19] sb_1__1__22_chanx_left_out;
  wire [0:19] sb_1__1__22_chanx_right_out;
  wire [0:19] sb_1__1__22_chany_bottom_out;
  wire [0:19] sb_1__1__22_chany_top_out;
  wire [0:0] sb_1__1__23_ccff_tail;
  wire [0:19] sb_1__1__23_chanx_left_out;
  wire [0:19] sb_1__1__23_chanx_right_out;
  wire [0:19] sb_1__1__23_chany_bottom_out;
  wire [0:19] sb_1__1__23_chany_top_out;
  wire [0:0] sb_1__1__24_ccff_tail;
  wire [0:19] sb_1__1__24_chanx_left_out;
  wire [0:19] sb_1__1__24_chanx_right_out;
  wire [0:19] sb_1__1__24_chany_bottom_out;
  wire [0:19] sb_1__1__24_chany_top_out;
  wire [0:0] sb_1__1__25_ccff_tail;
  wire [0:19] sb_1__1__25_chanx_left_out;
  wire [0:19] sb_1__1__25_chanx_right_out;
  wire [0:19] sb_1__1__25_chany_bottom_out;
  wire [0:19] sb_1__1__25_chany_top_out;
  wire [0:0] sb_1__1__26_ccff_tail;
  wire [0:19] sb_1__1__26_chanx_left_out;
  wire [0:19] sb_1__1__26_chanx_right_out;
  wire [0:19] sb_1__1__26_chany_bottom_out;
  wire [0:19] sb_1__1__26_chany_top_out;
  wire [0:0] sb_1__1__27_ccff_tail;
  wire [0:19] sb_1__1__27_chanx_left_out;
  wire [0:19] sb_1__1__27_chanx_right_out;
  wire [0:19] sb_1__1__27_chany_bottom_out;
  wire [0:19] sb_1__1__27_chany_top_out;
  wire [0:0] sb_1__1__28_ccff_tail;
  wire [0:19] sb_1__1__28_chanx_left_out;
  wire [0:19] sb_1__1__28_chanx_right_out;
  wire [0:19] sb_1__1__28_chany_bottom_out;
  wire [0:19] sb_1__1__28_chany_top_out;
  wire [0:0] sb_1__1__29_ccff_tail;
  wire [0:19] sb_1__1__29_chanx_left_out;
  wire [0:19] sb_1__1__29_chanx_right_out;
  wire [0:19] sb_1__1__29_chany_bottom_out;
  wire [0:19] sb_1__1__29_chany_top_out;
  wire [0:0] sb_1__1__2_ccff_tail;
  wire [0:19] sb_1__1__2_chanx_left_out;
  wire [0:19] sb_1__1__2_chanx_right_out;
  wire [0:19] sb_1__1__2_chany_bottom_out;
  wire [0:19] sb_1__1__2_chany_top_out;
  wire [0:0] sb_1__1__30_ccff_tail;
  wire [0:19] sb_1__1__30_chanx_left_out;
  wire [0:19] sb_1__1__30_chanx_right_out;
  wire [0:19] sb_1__1__30_chany_bottom_out;
  wire [0:19] sb_1__1__30_chany_top_out;
  wire [0:0] sb_1__1__31_ccff_tail;
  wire [0:19] sb_1__1__31_chanx_left_out;
  wire [0:19] sb_1__1__31_chanx_right_out;
  wire [0:19] sb_1__1__31_chany_bottom_out;
  wire [0:19] sb_1__1__31_chany_top_out;
  wire [0:0] sb_1__1__32_ccff_tail;
  wire [0:19] sb_1__1__32_chanx_left_out;
  wire [0:19] sb_1__1__32_chanx_right_out;
  wire [0:19] sb_1__1__32_chany_bottom_out;
  wire [0:19] sb_1__1__32_chany_top_out;
  wire [0:0] sb_1__1__33_ccff_tail;
  wire [0:19] sb_1__1__33_chanx_left_out;
  wire [0:19] sb_1__1__33_chanx_right_out;
  wire [0:19] sb_1__1__33_chany_bottom_out;
  wire [0:19] sb_1__1__33_chany_top_out;
  wire [0:0] sb_1__1__34_ccff_tail;
  wire [0:19] sb_1__1__34_chanx_left_out;
  wire [0:19] sb_1__1__34_chanx_right_out;
  wire [0:19] sb_1__1__34_chany_bottom_out;
  wire [0:19] sb_1__1__34_chany_top_out;
  wire [0:0] sb_1__1__35_ccff_tail;
  wire [0:19] sb_1__1__35_chanx_left_out;
  wire [0:19] sb_1__1__35_chanx_right_out;
  wire [0:19] sb_1__1__35_chany_bottom_out;
  wire [0:19] sb_1__1__35_chany_top_out;
  wire [0:0] sb_1__1__36_ccff_tail;
  wire [0:19] sb_1__1__36_chanx_left_out;
  wire [0:19] sb_1__1__36_chanx_right_out;
  wire [0:19] sb_1__1__36_chany_bottom_out;
  wire [0:19] sb_1__1__36_chany_top_out;
  wire [0:0] sb_1__1__37_ccff_tail;
  wire [0:19] sb_1__1__37_chanx_left_out;
  wire [0:19] sb_1__1__37_chanx_right_out;
  wire [0:19] sb_1__1__37_chany_bottom_out;
  wire [0:19] sb_1__1__37_chany_top_out;
  wire [0:0] sb_1__1__38_ccff_tail;
  wire [0:19] sb_1__1__38_chanx_left_out;
  wire [0:19] sb_1__1__38_chanx_right_out;
  wire [0:19] sb_1__1__38_chany_bottom_out;
  wire [0:19] sb_1__1__38_chany_top_out;
  wire [0:0] sb_1__1__39_ccff_tail;
  wire [0:19] sb_1__1__39_chanx_left_out;
  wire [0:19] sb_1__1__39_chanx_right_out;
  wire [0:19] sb_1__1__39_chany_bottom_out;
  wire [0:19] sb_1__1__39_chany_top_out;
  wire [0:0] sb_1__1__3_ccff_tail;
  wire [0:19] sb_1__1__3_chanx_left_out;
  wire [0:19] sb_1__1__3_chanx_right_out;
  wire [0:19] sb_1__1__3_chany_bottom_out;
  wire [0:19] sb_1__1__3_chany_top_out;
  wire [0:0] sb_1__1__40_ccff_tail;
  wire [0:19] sb_1__1__40_chanx_left_out;
  wire [0:19] sb_1__1__40_chanx_right_out;
  wire [0:19] sb_1__1__40_chany_bottom_out;
  wire [0:19] sb_1__1__40_chany_top_out;
  wire [0:0] sb_1__1__41_ccff_tail;
  wire [0:19] sb_1__1__41_chanx_left_out;
  wire [0:19] sb_1__1__41_chanx_right_out;
  wire [0:19] sb_1__1__41_chany_bottom_out;
  wire [0:19] sb_1__1__41_chany_top_out;
  wire [0:0] sb_1__1__42_ccff_tail;
  wire [0:19] sb_1__1__42_chanx_left_out;
  wire [0:19] sb_1__1__42_chanx_right_out;
  wire [0:19] sb_1__1__42_chany_bottom_out;
  wire [0:19] sb_1__1__42_chany_top_out;
  wire [0:0] sb_1__1__43_ccff_tail;
  wire [0:19] sb_1__1__43_chanx_left_out;
  wire [0:19] sb_1__1__43_chanx_right_out;
  wire [0:19] sb_1__1__43_chany_bottom_out;
  wire [0:19] sb_1__1__43_chany_top_out;
  wire [0:0] sb_1__1__44_ccff_tail;
  wire [0:19] sb_1__1__44_chanx_left_out;
  wire [0:19] sb_1__1__44_chanx_right_out;
  wire [0:19] sb_1__1__44_chany_bottom_out;
  wire [0:19] sb_1__1__44_chany_top_out;
  wire [0:0] sb_1__1__45_ccff_tail;
  wire [0:19] sb_1__1__45_chanx_left_out;
  wire [0:19] sb_1__1__45_chanx_right_out;
  wire [0:19] sb_1__1__45_chany_bottom_out;
  wire [0:19] sb_1__1__45_chany_top_out;
  wire [0:0] sb_1__1__46_ccff_tail;
  wire [0:19] sb_1__1__46_chanx_left_out;
  wire [0:19] sb_1__1__46_chanx_right_out;
  wire [0:19] sb_1__1__46_chany_bottom_out;
  wire [0:19] sb_1__1__46_chany_top_out;
  wire [0:0] sb_1__1__47_ccff_tail;
  wire [0:19] sb_1__1__47_chanx_left_out;
  wire [0:19] sb_1__1__47_chanx_right_out;
  wire [0:19] sb_1__1__47_chany_bottom_out;
  wire [0:19] sb_1__1__47_chany_top_out;
  wire [0:0] sb_1__1__48_ccff_tail;
  wire [0:19] sb_1__1__48_chanx_left_out;
  wire [0:19] sb_1__1__48_chanx_right_out;
  wire [0:19] sb_1__1__48_chany_bottom_out;
  wire [0:19] sb_1__1__48_chany_top_out;
  wire [0:0] sb_1__1__4_ccff_tail;
  wire [0:19] sb_1__1__4_chanx_left_out;
  wire [0:19] sb_1__1__4_chanx_right_out;
  wire [0:19] sb_1__1__4_chany_bottom_out;
  wire [0:19] sb_1__1__4_chany_top_out;
  wire [0:0] sb_1__1__5_ccff_tail;
  wire [0:19] sb_1__1__5_chanx_left_out;
  wire [0:19] sb_1__1__5_chanx_right_out;
  wire [0:19] sb_1__1__5_chany_bottom_out;
  wire [0:19] sb_1__1__5_chany_top_out;
  wire [0:0] sb_1__1__6_ccff_tail;
  wire [0:19] sb_1__1__6_chanx_left_out;
  wire [0:19] sb_1__1__6_chanx_right_out;
  wire [0:19] sb_1__1__6_chany_bottom_out;
  wire [0:19] sb_1__1__6_chany_top_out;
  wire [0:0] sb_1__1__7_ccff_tail;
  wire [0:19] sb_1__1__7_chanx_left_out;
  wire [0:19] sb_1__1__7_chanx_right_out;
  wire [0:19] sb_1__1__7_chany_bottom_out;
  wire [0:19] sb_1__1__7_chany_top_out;
  wire [0:0] sb_1__1__8_ccff_tail;
  wire [0:19] sb_1__1__8_chanx_left_out;
  wire [0:19] sb_1__1__8_chanx_right_out;
  wire [0:19] sb_1__1__8_chany_bottom_out;
  wire [0:19] sb_1__1__8_chany_top_out;
  wire [0:0] sb_1__1__9_ccff_tail;
  wire [0:19] sb_1__1__9_chanx_left_out;
  wire [0:19] sb_1__1__9_chanx_right_out;
  wire [0:19] sb_1__1__9_chany_bottom_out;
  wire [0:19] sb_1__1__9_chany_top_out;
  wire [0:0] sb_1__8__0_ccff_tail;
  wire [0:19] sb_1__8__0_chanx_left_out;
  wire [0:19] sb_1__8__0_chanx_right_out;
  wire [0:19] sb_1__8__0_chany_bottom_out;
  wire [0:0] sb_1__8__1_ccff_tail;
  wire [0:19] sb_1__8__1_chanx_left_out;
  wire [0:19] sb_1__8__1_chanx_right_out;
  wire [0:19] sb_1__8__1_chany_bottom_out;
  wire [0:0] sb_1__8__2_ccff_tail;
  wire [0:19] sb_1__8__2_chanx_left_out;
  wire [0:19] sb_1__8__2_chanx_right_out;
  wire [0:19] sb_1__8__2_chany_bottom_out;
  wire [0:0] sb_1__8__3_ccff_tail;
  wire [0:19] sb_1__8__3_chanx_left_out;
  wire [0:19] sb_1__8__3_chanx_right_out;
  wire [0:19] sb_1__8__3_chany_bottom_out;
  wire [0:0] sb_1__8__4_ccff_tail;
  wire [0:19] sb_1__8__4_chanx_left_out;
  wire [0:19] sb_1__8__4_chanx_right_out;
  wire [0:19] sb_1__8__4_chany_bottom_out;
  wire [0:0] sb_1__8__5_ccff_tail;
  wire [0:19] sb_1__8__5_chanx_left_out;
  wire [0:19] sb_1__8__5_chanx_right_out;
  wire [0:19] sb_1__8__5_chany_bottom_out;
  wire [0:0] sb_1__8__6_ccff_tail;
  wire [0:19] sb_1__8__6_chanx_left_out;
  wire [0:19] sb_1__8__6_chanx_right_out;
  wire [0:19] sb_1__8__6_chany_bottom_out;
  wire [0:0] sb_8__0__0_ccff_tail;
  wire [0:19] sb_8__0__0_chanx_left_out;
  wire [0:19] sb_8__0__0_chany_top_out;
  wire [0:0] sb_8__1__0_ccff_tail;
  wire [0:19] sb_8__1__0_chanx_left_out;
  wire [0:19] sb_8__1__0_chany_bottom_out;
  wire [0:19] sb_8__1__0_chany_top_out;
  wire [0:0] sb_8__1__1_ccff_tail;
  wire [0:19] sb_8__1__1_chanx_left_out;
  wire [0:19] sb_8__1__1_chany_bottom_out;
  wire [0:19] sb_8__1__1_chany_top_out;
  wire [0:0] sb_8__1__2_ccff_tail;
  wire [0:19] sb_8__1__2_chanx_left_out;
  wire [0:19] sb_8__1__2_chany_bottom_out;
  wire [0:19] sb_8__1__2_chany_top_out;
  wire [0:0] sb_8__1__3_ccff_tail;
  wire [0:19] sb_8__1__3_chanx_left_out;
  wire [0:19] sb_8__1__3_chany_bottom_out;
  wire [0:19] sb_8__1__3_chany_top_out;
  wire [0:0] sb_8__1__4_ccff_tail;
  wire [0:19] sb_8__1__4_chanx_left_out;
  wire [0:19] sb_8__1__4_chany_bottom_out;
  wire [0:19] sb_8__1__4_chany_top_out;
  wire [0:0] sb_8__1__5_ccff_tail;
  wire [0:19] sb_8__1__5_chanx_left_out;
  wire [0:19] sb_8__1__5_chany_bottom_out;
  wire [0:19] sb_8__1__5_chany_top_out;
  wire [0:0] sb_8__1__6_ccff_tail;
  wire [0:19] sb_8__1__6_chanx_left_out;
  wire [0:19] sb_8__1__6_chany_bottom_out;
  wire [0:19] sb_8__1__6_chany_top_out;
  wire [0:0] sb_8__8__0_ccff_tail;
  wire [0:19] sb_8__8__0_chanx_left_out;
  wire [0:19] sb_8__8__0_chany_bottom_out;
  wire [1:0] UNCONN;
  wire [147:0] scff_Wires;
  wire [56:0] regin_feedthrough_wires;
  wire [56:0] regout_feedthrough_wires;
  wire [127:0] Test_enWires;
  wire [288:0] prog_clk_0_wires;
  wire [111:0] prog_clk_1_wires;
  wire [51:0] prog_clk_2_wires;
  wire [34:0] prog_clk_3_wires;
  wire [111:0] clk_1_wires;
  wire [51:0] clk_2_wires;
  wire [34:0] clk_3_wires;

  grid_clb
  grid_clb_1__1_
  (
    .clk_0_N_in(clk_1_wires[4]),
    .prog_clk_0_N_in(prog_clk_1_wires[4]),
    .prog_clk_0_W_out(prog_clk_0_wires[3]),
    .prog_clk_0_E_out(prog_clk_0_wires[1]),
    .prog_clk_0_S_out(prog_clk_0_wires[0]),
    .Test_en_E_in(Test_enWires[16]),
    .SC_OUT_BOT(scff_Wires[17]),
    .SC_IN_TOP(scff_Wires[15]),
    .top_width_0_height_0__pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_0_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_0_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_0_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_0_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_0_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_0_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_0_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_0_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_0_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_1__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_0_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__2_
  (
    .clk_0_S_in(clk_1_wires[3]),
    .prog_clk_0_S_in(prog_clk_1_wires[3]),
    .prog_clk_0_W_out(prog_clk_0_wires[9]),
    .prog_clk_0_E_out(prog_clk_0_wires[7]),
    .prog_clk_0_S_out(prog_clk_0_wires[6]),
    .Test_en_E_in(Test_enWires[30]),
    .SC_OUT_BOT(scff_Wires[14]),
    .SC_IN_TOP(scff_Wires[13]),
    .top_width_0_height_0__pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[1]),
    .right_width_0_height_0__pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_1_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_1_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_1_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_1_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_1_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_1_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_1_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_1_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_1_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[0]),
    .ccff_tail(grid_clb_1_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__3_
  (
    .clk_0_N_in(clk_1_wires[11]),
    .prog_clk_0_N_in(prog_clk_1_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[14]),
    .prog_clk_0_E_out(prog_clk_0_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[11]),
    .Test_en_E_in(Test_enWires[44]),
    .SC_OUT_BOT(scff_Wires[12]),
    .SC_IN_TOP(scff_Wires[11]),
    .top_width_0_height_0__pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[2]),
    .right_width_0_height_0__pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_2_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_2_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_2_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_2_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_2_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_2_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_2_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_2_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_2_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[1]),
    .ccff_tail(grid_clb_2_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__4_
  (
    .clk_0_S_in(clk_1_wires[10]),
    .prog_clk_0_S_in(prog_clk_1_wires[10]),
    .prog_clk_0_W_out(prog_clk_0_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[17]),
    .prog_clk_0_S_out(prog_clk_0_wires[16]),
    .Test_en_E_in(Test_enWires[58]),
    .SC_OUT_BOT(scff_Wires[10]),
    .SC_IN_TOP(scff_Wires[9]),
    .top_width_0_height_0__pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[3]),
    .right_width_0_height_0__pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_3_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_3_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_3_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_3_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_3_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_3_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_3_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_3_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_3_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[2]),
    .ccff_tail(grid_clb_3_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__5_
  (
    .clk_0_N_in(clk_1_wires[18]),
    .prog_clk_0_N_in(prog_clk_1_wires[18]),
    .prog_clk_0_W_out(prog_clk_0_wires[24]),
    .prog_clk_0_E_out(prog_clk_0_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[21]),
    .Test_en_E_in(Test_enWires[72]),
    .SC_OUT_BOT(scff_Wires[8]),
    .SC_IN_TOP(scff_Wires[7]),
    .top_width_0_height_0__pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[4]),
    .right_width_0_height_0__pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_4_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_4_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_4_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_4_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_4_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_4_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_4_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_4_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_4_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[3]),
    .ccff_tail(grid_clb_4_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__6_
  (
    .clk_0_S_in(clk_1_wires[17]),
    .prog_clk_0_S_in(prog_clk_1_wires[17]),
    .prog_clk_0_W_out(prog_clk_0_wires[29]),
    .prog_clk_0_E_out(prog_clk_0_wires[27]),
    .prog_clk_0_S_out(prog_clk_0_wires[26]),
    .Test_en_E_in(Test_enWires[86]),
    .SC_OUT_BOT(scff_Wires[6]),
    .SC_IN_TOP(scff_Wires[5]),
    .top_width_0_height_0__pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[5]),
    .right_width_0_height_0__pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_5_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_5_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_5_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_5_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_5_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_5_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_5_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_5_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_5_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[4]),
    .ccff_tail(grid_clb_5_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__7_
  (
    .clk_0_N_in(clk_1_wires[25]),
    .prog_clk_0_N_in(prog_clk_1_wires[25]),
    .prog_clk_0_W_out(prog_clk_0_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[32]),
    .prog_clk_0_S_out(prog_clk_0_wires[31]),
    .Test_en_E_in(Test_enWires[100]),
    .SC_OUT_BOT(scff_Wires[4]),
    .SC_IN_TOP(scff_Wires[3]),
    .top_width_0_height_0__pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[6]),
    .right_width_0_height_0__pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_6_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_6_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_6_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_6_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_6_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_6_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_6_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_6_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_6_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[5]),
    .ccff_tail(grid_clb_6_ccff_tail[0])
  );


  grid_clb
  grid_clb_1__8_
  (
    .clk_0_S_in(clk_1_wires[24]),
    .prog_clk_0_S_in(prog_clk_1_wires[24]),
    .prog_clk_0_W_out(prog_clk_0_wires[41]),
    .prog_clk_0_N_out(prog_clk_0_wires[39]),
    .prog_clk_0_E_out(prog_clk_0_wires[37]),
    .prog_clk_0_S_out(prog_clk_0_wires[36]),
    .Test_en_E_in(Test_enWires[114]),
    .SC_OUT_BOT(scff_Wires[2]),
    .SC_IN_TOP(scff_Wires[1]),
    .top_width_0_height_0__pin_0_(cbx_1__8__0_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__0_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__0_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__0_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__0_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__0_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__0_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__0_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__0_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_1__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
    .ccff_head(grid_io_left_7_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_7_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_7_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_7_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_7_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_7_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_7_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_7_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_7_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[6]),
    .ccff_tail(grid_clb_7_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__1_
  (
    .clk_0_N_in(clk_1_wires[6]),
    .prog_clk_0_N_in(prog_clk_1_wires[6]),
    .prog_clk_0_E_out(prog_clk_0_wires[44]),
    .prog_clk_0_S_out(prog_clk_0_wires[43]),
    .Test_en_W_out(Test_enWires[18]),
    .Test_en_E_in(Test_enWires[17]),
    .SC_OUT_TOP(scff_Wires[21]),
    .SC_IN_BOT(scff_Wires[20]),
    .top_width_0_height_0__pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[7]),
    .right_width_0_height_0__pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__0_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_8_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_8_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_8_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_8_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_8_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_8_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_8_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_8_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_2__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_8_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__2_
  (
    .clk_0_S_in(clk_1_wires[5]),
    .prog_clk_0_S_in(prog_clk_1_wires[5]),
    .prog_clk_0_E_out(prog_clk_0_wires[47]),
    .prog_clk_0_S_out(prog_clk_0_wires[46]),
    .Test_en_W_out(Test_enWires[32]),
    .Test_en_E_in(Test_enWires[31]),
    .SC_OUT_TOP(scff_Wires[23]),
    .SC_IN_BOT(scff_Wires[22]),
    .top_width_0_height_0__pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[8]),
    .right_width_0_height_0__pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__1_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_9_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_9_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_9_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_9_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_9_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_9_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_9_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_9_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[7]),
    .ccff_tail(grid_clb_9_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__3_
  (
    .clk_0_N_in(clk_1_wires[13]),
    .prog_clk_0_N_in(prog_clk_1_wires[13]),
    .prog_clk_0_E_out(prog_clk_0_wires[50]),
    .prog_clk_0_S_out(prog_clk_0_wires[49]),
    .Test_en_W_out(Test_enWires[46]),
    .Test_en_E_in(Test_enWires[45]),
    .SC_OUT_TOP(scff_Wires[25]),
    .SC_IN_BOT(scff_Wires[24]),
    .top_width_0_height_0__pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[9]),
    .right_width_0_height_0__pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__2_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_10_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_10_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_10_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_10_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_10_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_10_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_10_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_10_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[8]),
    .ccff_tail(grid_clb_10_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__4_
  (
    .clk_0_S_in(clk_1_wires[12]),
    .prog_clk_0_S_in(prog_clk_1_wires[12]),
    .prog_clk_0_E_out(prog_clk_0_wires[53]),
    .prog_clk_0_S_out(prog_clk_0_wires[52]),
    .Test_en_W_out(Test_enWires[60]),
    .Test_en_E_in(Test_enWires[59]),
    .SC_OUT_TOP(scff_Wires[27]),
    .SC_IN_BOT(scff_Wires[26]),
    .top_width_0_height_0__pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[10]),
    .right_width_0_height_0__pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__3_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_11_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_11_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_11_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_11_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_11_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_11_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_11_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_11_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[9]),
    .ccff_tail(grid_clb_11_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__5_
  (
    .clk_0_N_in(clk_1_wires[20]),
    .prog_clk_0_N_in(prog_clk_1_wires[20]),
    .prog_clk_0_E_out(prog_clk_0_wires[56]),
    .prog_clk_0_S_out(prog_clk_0_wires[55]),
    .Test_en_W_out(Test_enWires[74]),
    .Test_en_E_in(Test_enWires[73]),
    .SC_OUT_TOP(scff_Wires[29]),
    .SC_IN_BOT(scff_Wires[28]),
    .top_width_0_height_0__pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[11]),
    .right_width_0_height_0__pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__4_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_12_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_12_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_12_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_12_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_12_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_12_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_12_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_12_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[10]),
    .ccff_tail(grid_clb_12_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__6_
  (
    .clk_0_S_in(clk_1_wires[19]),
    .prog_clk_0_S_in(prog_clk_1_wires[19]),
    .prog_clk_0_E_out(prog_clk_0_wires[59]),
    .prog_clk_0_S_out(prog_clk_0_wires[58]),
    .Test_en_W_out(Test_enWires[88]),
    .Test_en_E_in(Test_enWires[87]),
    .SC_OUT_TOP(scff_Wires[31]),
    .SC_IN_BOT(scff_Wires[30]),
    .top_width_0_height_0__pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[12]),
    .right_width_0_height_0__pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__5_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_13_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_13_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_13_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_13_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_13_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_13_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_13_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_13_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[11]),
    .ccff_tail(grid_clb_13_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__7_
  (
    .clk_0_N_in(clk_1_wires[27]),
    .prog_clk_0_N_in(prog_clk_1_wires[27]),
    .prog_clk_0_E_out(prog_clk_0_wires[62]),
    .prog_clk_0_S_out(prog_clk_0_wires[61]),
    .Test_en_W_out(Test_enWires[102]),
    .Test_en_E_in(Test_enWires[101]),
    .SC_OUT_TOP(scff_Wires[33]),
    .SC_IN_BOT(scff_Wires[32]),
    .top_width_0_height_0__pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[13]),
    .right_width_0_height_0__pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__6_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_14_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_14_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_14_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_14_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_14_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_14_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_14_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_14_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[12]),
    .ccff_tail(grid_clb_14_ccff_tail[0])
  );


  grid_clb
  grid_clb_2__8_
  (
    .clk_0_S_in(clk_1_wires[26]),
    .prog_clk_0_S_in(prog_clk_1_wires[26]),
    .prog_clk_0_N_out(prog_clk_0_wires[67]),
    .prog_clk_0_E_out(prog_clk_0_wires[65]),
    .prog_clk_0_S_out(prog_clk_0_wires[64]),
    .Test_en_W_out(Test_enWires[116]),
    .Test_en_E_in(Test_enWires[115]),
    .SC_OUT_TOP(scff_Wires[35]),
    .SC_IN_BOT(scff_Wires[34]),
    .top_width_0_height_0__pin_0_(cbx_1__8__1_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__1_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__1_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__1_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__1_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__1_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__1_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__1_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__1_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_2__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__7_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_15_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_15_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_15_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_15_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_15_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_15_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_15_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_15_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[13]),
    .ccff_tail(grid_clb_15_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__1_
  (
    .clk_0_N_in(clk_1_wires[32]),
    .prog_clk_0_N_in(prog_clk_1_wires[32]),
    .prog_clk_0_E_out(prog_clk_0_wires[70]),
    .prog_clk_0_S_out(prog_clk_0_wires[69]),
    .Test_en_W_out(Test_enWires[20]),
    .Test_en_E_in(Test_enWires[19]),
    .SC_OUT_BOT(scff_Wires[54]),
    .SC_IN_TOP(scff_Wires[52]),
    .top_width_0_height_0__pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[14]),
    .right_width_0_height_0__pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__8_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_16_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_16_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_16_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_16_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_16_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_16_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_16_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_16_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_3__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_16_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__2_
  (
    .clk_0_S_in(clk_1_wires[31]),
    .prog_clk_0_S_in(prog_clk_1_wires[31]),
    .prog_clk_0_E_out(prog_clk_0_wires[73]),
    .prog_clk_0_S_out(prog_clk_0_wires[72]),
    .Test_en_W_out(Test_enWires[34]),
    .Test_en_E_in(Test_enWires[33]),
    .SC_OUT_BOT(scff_Wires[51]),
    .SC_IN_TOP(scff_Wires[50]),
    .top_width_0_height_0__pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[15]),
    .right_width_0_height_0__pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__9_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_17_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_17_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_17_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_17_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_17_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_17_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_17_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_17_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[14]),
    .ccff_tail(grid_clb_17_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__3_
  (
    .clk_0_N_in(clk_1_wires[39]),
    .prog_clk_0_N_in(prog_clk_1_wires[39]),
    .prog_clk_0_E_out(prog_clk_0_wires[76]),
    .prog_clk_0_S_out(prog_clk_0_wires[75]),
    .Test_en_W_out(Test_enWires[48]),
    .Test_en_E_in(Test_enWires[47]),
    .SC_OUT_BOT(scff_Wires[49]),
    .SC_IN_TOP(scff_Wires[48]),
    .top_width_0_height_0__pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[16]),
    .right_width_0_height_0__pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__10_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_18_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_18_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_18_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_18_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_18_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_18_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_18_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_18_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[15]),
    .ccff_tail(grid_clb_18_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__4_
  (
    .clk_0_S_in(clk_1_wires[38]),
    .prog_clk_0_S_in(prog_clk_1_wires[38]),
    .prog_clk_0_E_out(prog_clk_0_wires[79]),
    .prog_clk_0_S_out(prog_clk_0_wires[78]),
    .Test_en_W_out(Test_enWires[62]),
    .Test_en_E_in(Test_enWires[61]),
    .SC_OUT_BOT(scff_Wires[47]),
    .SC_IN_TOP(scff_Wires[46]),
    .top_width_0_height_0__pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[17]),
    .right_width_0_height_0__pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__11_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_19_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_19_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_19_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_19_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_19_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_19_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_19_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_19_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[16]),
    .ccff_tail(grid_clb_19_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__5_
  (
    .clk_0_N_in(clk_1_wires[46]),
    .prog_clk_0_N_in(prog_clk_1_wires[46]),
    .prog_clk_0_E_out(prog_clk_0_wires[82]),
    .prog_clk_0_S_out(prog_clk_0_wires[81]),
    .Test_en_W_out(Test_enWires[76]),
    .Test_en_E_in(Test_enWires[75]),
    .SC_OUT_BOT(scff_Wires[45]),
    .SC_IN_TOP(scff_Wires[44]),
    .top_width_0_height_0__pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[18]),
    .right_width_0_height_0__pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__12_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_20_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_20_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_20_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_20_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_20_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_20_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_20_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_20_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[17]),
    .ccff_tail(grid_clb_20_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__6_
  (
    .clk_0_S_in(clk_1_wires[45]),
    .prog_clk_0_S_in(prog_clk_1_wires[45]),
    .prog_clk_0_E_out(prog_clk_0_wires[85]),
    .prog_clk_0_S_out(prog_clk_0_wires[84]),
    .Test_en_W_out(Test_enWires[90]),
    .Test_en_E_in(Test_enWires[89]),
    .SC_OUT_BOT(scff_Wires[43]),
    .SC_IN_TOP(scff_Wires[42]),
    .top_width_0_height_0__pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[19]),
    .right_width_0_height_0__pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__13_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_21_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_21_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_21_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_21_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_21_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_21_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_21_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_21_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[18]),
    .ccff_tail(grid_clb_21_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__7_
  (
    .clk_0_N_in(clk_1_wires[53]),
    .prog_clk_0_N_in(prog_clk_1_wires[53]),
    .prog_clk_0_E_out(prog_clk_0_wires[88]),
    .prog_clk_0_S_out(prog_clk_0_wires[87]),
    .Test_en_W_out(Test_enWires[104]),
    .Test_en_E_in(Test_enWires[103]),
    .SC_OUT_BOT(scff_Wires[41]),
    .SC_IN_TOP(scff_Wires[40]),
    .top_width_0_height_0__pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[20]),
    .right_width_0_height_0__pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__14_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_22_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_22_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_22_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_22_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_22_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_22_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_22_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_22_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[19]),
    .ccff_tail(grid_clb_22_ccff_tail[0])
  );


  grid_clb
  grid_clb_3__8_
  (
    .clk_0_S_in(clk_1_wires[52]),
    .prog_clk_0_S_in(prog_clk_1_wires[52]),
    .prog_clk_0_N_out(prog_clk_0_wires[93]),
    .prog_clk_0_E_out(prog_clk_0_wires[91]),
    .prog_clk_0_S_out(prog_clk_0_wires[90]),
    .Test_en_W_out(Test_enWires[118]),
    .Test_en_E_in(Test_enWires[117]),
    .SC_OUT_BOT(scff_Wires[39]),
    .SC_IN_TOP(scff_Wires[38]),
    .top_width_0_height_0__pin_0_(cbx_1__8__2_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__2_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__2_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__2_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__2_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__2_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__2_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__2_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__2_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_3__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__15_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_23_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_23_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_23_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_23_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_23_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_23_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_23_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_23_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[20]),
    .ccff_tail(grid_clb_23_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__1_
  (
    .clk_0_N_in(clk_1_wires[34]),
    .prog_clk_0_N_in(prog_clk_1_wires[34]),
    .prog_clk_0_E_out(prog_clk_0_wires[96]),
    .prog_clk_0_S_out(prog_clk_0_wires[95]),
    .Test_en_W_out(Test_enWires[22]),
    .Test_en_E_in(Test_enWires[21]),
    .SC_OUT_TOP(scff_Wires[58]),
    .SC_IN_BOT(scff_Wires[57]),
    .top_width_0_height_0__pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[21]),
    .right_width_0_height_0__pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__16_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_24_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_24_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_24_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_24_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_24_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_24_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_24_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_24_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_4__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_24_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__2_
  (
    .clk_0_S_in(clk_1_wires[33]),
    .prog_clk_0_S_in(prog_clk_1_wires[33]),
    .prog_clk_0_E_out(prog_clk_0_wires[99]),
    .prog_clk_0_S_out(prog_clk_0_wires[98]),
    .Test_en_W_out(Test_enWires[36]),
    .Test_en_E_in(Test_enWires[35]),
    .SC_OUT_TOP(scff_Wires[60]),
    .SC_IN_BOT(scff_Wires[59]),
    .top_width_0_height_0__pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[22]),
    .right_width_0_height_0__pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__17_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_25_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_25_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_25_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_25_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_25_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_25_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_25_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_25_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[21]),
    .ccff_tail(grid_clb_25_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__3_
  (
    .clk_0_N_in(clk_1_wires[41]),
    .prog_clk_0_N_in(prog_clk_1_wires[41]),
    .prog_clk_0_E_out(prog_clk_0_wires[102]),
    .prog_clk_0_S_out(prog_clk_0_wires[101]),
    .Test_en_W_out(Test_enWires[50]),
    .Test_en_E_in(Test_enWires[49]),
    .SC_OUT_TOP(scff_Wires[62]),
    .SC_IN_BOT(scff_Wires[61]),
    .top_width_0_height_0__pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[23]),
    .right_width_0_height_0__pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__18_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_26_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_26_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_26_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_26_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_26_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_26_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_26_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_26_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[22]),
    .ccff_tail(grid_clb_26_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__4_
  (
    .clk_0_S_in(clk_1_wires[40]),
    .prog_clk_0_S_in(prog_clk_1_wires[40]),
    .prog_clk_0_E_out(prog_clk_0_wires[105]),
    .prog_clk_0_S_out(prog_clk_0_wires[104]),
    .Test_en_W_out(Test_enWires[64]),
    .Test_en_E_in(Test_enWires[63]),
    .SC_OUT_TOP(scff_Wires[64]),
    .SC_IN_BOT(scff_Wires[63]),
    .top_width_0_height_0__pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[24]),
    .right_width_0_height_0__pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__19_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_27_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_27_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_27_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_27_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_27_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_27_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_27_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_27_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[23]),
    .ccff_tail(grid_clb_27_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__5_
  (
    .clk_0_N_in(clk_1_wires[48]),
    .prog_clk_0_N_in(prog_clk_1_wires[48]),
    .prog_clk_0_E_out(prog_clk_0_wires[108]),
    .prog_clk_0_S_out(prog_clk_0_wires[107]),
    .Test_en_W_out(Test_enWires[78]),
    .Test_en_E_in(Test_enWires[77]),
    .SC_OUT_TOP(scff_Wires[66]),
    .SC_IN_BOT(scff_Wires[65]),
    .top_width_0_height_0__pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[25]),
    .right_width_0_height_0__pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__20_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_28_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_28_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_28_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_28_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_28_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_28_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_28_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_28_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[24]),
    .ccff_tail(grid_clb_28_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__6_
  (
    .clk_0_S_in(clk_1_wires[47]),
    .prog_clk_0_S_in(prog_clk_1_wires[47]),
    .prog_clk_0_E_out(prog_clk_0_wires[111]),
    .prog_clk_0_S_out(prog_clk_0_wires[110]),
    .Test_en_W_out(Test_enWires[92]),
    .Test_en_E_in(Test_enWires[91]),
    .SC_OUT_TOP(scff_Wires[68]),
    .SC_IN_BOT(scff_Wires[67]),
    .top_width_0_height_0__pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[26]),
    .right_width_0_height_0__pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__21_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_29_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_29_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_29_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_29_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_29_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_29_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_29_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_29_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[25]),
    .ccff_tail(grid_clb_29_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__7_
  (
    .clk_0_N_in(clk_1_wires[55]),
    .prog_clk_0_N_in(prog_clk_1_wires[55]),
    .prog_clk_0_E_out(prog_clk_0_wires[114]),
    .prog_clk_0_S_out(prog_clk_0_wires[113]),
    .Test_en_W_out(Test_enWires[106]),
    .Test_en_E_in(Test_enWires[105]),
    .SC_OUT_TOP(scff_Wires[70]),
    .SC_IN_BOT(scff_Wires[69]),
    .top_width_0_height_0__pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[27]),
    .right_width_0_height_0__pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__22_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_30_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_30_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_30_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_30_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_30_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_30_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_30_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_30_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[26]),
    .ccff_tail(grid_clb_30_ccff_tail[0])
  );


  grid_clb
  grid_clb_4__8_
  (
    .clk_0_S_in(clk_1_wires[54]),
    .prog_clk_0_S_in(prog_clk_1_wires[54]),
    .prog_clk_0_N_out(prog_clk_0_wires[119]),
    .prog_clk_0_E_out(prog_clk_0_wires[117]),
    .prog_clk_0_S_out(prog_clk_0_wires[116]),
    .Test_en_W_out(Test_enWires[120]),
    .Test_en_E_in(Test_enWires[119]),
    .SC_OUT_TOP(scff_Wires[72]),
    .SC_IN_BOT(scff_Wires[71]),
    .top_width_0_height_0__pin_0_(cbx_1__8__3_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__3_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__3_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__3_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__3_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__3_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__3_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__3_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__3_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_4__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__23_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_31_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_31_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_31_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_31_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_31_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_31_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_31_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_31_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[27]),
    .ccff_tail(grid_clb_31_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__1_
  (
    .clk_0_N_in(clk_1_wires[60]),
    .prog_clk_0_N_in(prog_clk_1_wires[60]),
    .prog_clk_0_E_out(prog_clk_0_wires[122]),
    .prog_clk_0_S_out(prog_clk_0_wires[121]),
    .Test_en_E_out(Test_enWires[24]),
    .Test_en_W_in(Test_enWires[23]),
    .SC_OUT_BOT(scff_Wires[91]),
    .SC_IN_TOP(scff_Wires[89]),
    .top_width_0_height_0__pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[28]),
    .right_width_0_height_0__pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__24_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_32_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_32_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_32_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_32_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_32_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_32_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_32_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_32_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_5__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_32_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__2_
  (
    .clk_0_S_in(clk_1_wires[59]),
    .prog_clk_0_S_in(prog_clk_1_wires[59]),
    .prog_clk_0_E_out(prog_clk_0_wires[125]),
    .prog_clk_0_S_out(prog_clk_0_wires[124]),
    .Test_en_E_out(Test_enWires[38]),
    .Test_en_W_in(Test_enWires[37]),
    .SC_OUT_BOT(scff_Wires[88]),
    .SC_IN_TOP(scff_Wires[87]),
    .top_width_0_height_0__pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[29]),
    .right_width_0_height_0__pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__25_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_33_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_33_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_33_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_33_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_33_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_33_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_33_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_33_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[28]),
    .ccff_tail(grid_clb_33_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__3_
  (
    .clk_0_N_in(clk_1_wires[67]),
    .prog_clk_0_N_in(prog_clk_1_wires[67]),
    .prog_clk_0_E_out(prog_clk_0_wires[128]),
    .prog_clk_0_S_out(prog_clk_0_wires[127]),
    .Test_en_E_out(Test_enWires[52]),
    .Test_en_W_in(Test_enWires[51]),
    .SC_OUT_BOT(scff_Wires[86]),
    .SC_IN_TOP(scff_Wires[85]),
    .top_width_0_height_0__pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[30]),
    .right_width_0_height_0__pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__26_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_34_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_34_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_34_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_34_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_34_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_34_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_34_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_34_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[29]),
    .ccff_tail(grid_clb_34_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__4_
  (
    .clk_0_S_in(clk_1_wires[66]),
    .prog_clk_0_S_in(prog_clk_1_wires[66]),
    .prog_clk_0_E_out(prog_clk_0_wires[131]),
    .prog_clk_0_S_out(prog_clk_0_wires[130]),
    .Test_en_E_out(Test_enWires[66]),
    .Test_en_W_in(Test_enWires[65]),
    .SC_OUT_BOT(scff_Wires[84]),
    .SC_IN_TOP(scff_Wires[83]),
    .top_width_0_height_0__pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[31]),
    .right_width_0_height_0__pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__27_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_35_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_35_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_35_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_35_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_35_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_35_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_35_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_35_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[30]),
    .ccff_tail(grid_clb_35_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__5_
  (
    .clk_0_N_in(clk_1_wires[74]),
    .prog_clk_0_N_in(prog_clk_1_wires[74]),
    .prog_clk_0_E_out(prog_clk_0_wires[134]),
    .prog_clk_0_S_out(prog_clk_0_wires[133]),
    .Test_en_E_out(Test_enWires[80]),
    .Test_en_W_in(Test_enWires[79]),
    .SC_OUT_BOT(scff_Wires[82]),
    .SC_IN_TOP(scff_Wires[81]),
    .top_width_0_height_0__pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[32]),
    .right_width_0_height_0__pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__28_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_36_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_36_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_36_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_36_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_36_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_36_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_36_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_36_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[31]),
    .ccff_tail(grid_clb_36_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__6_
  (
    .clk_0_S_in(clk_1_wires[73]),
    .prog_clk_0_S_in(prog_clk_1_wires[73]),
    .prog_clk_0_E_out(prog_clk_0_wires[137]),
    .prog_clk_0_S_out(prog_clk_0_wires[136]),
    .Test_en_E_out(Test_enWires[94]),
    .Test_en_W_in(Test_enWires[93]),
    .SC_OUT_BOT(scff_Wires[80]),
    .SC_IN_TOP(scff_Wires[79]),
    .top_width_0_height_0__pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[33]),
    .right_width_0_height_0__pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__29_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_37_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_37_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_37_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_37_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_37_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_37_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_37_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_37_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[32]),
    .ccff_tail(grid_clb_37_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__7_
  (
    .clk_0_N_in(clk_1_wires[81]),
    .prog_clk_0_N_in(prog_clk_1_wires[81]),
    .prog_clk_0_E_out(prog_clk_0_wires[140]),
    .prog_clk_0_S_out(prog_clk_0_wires[139]),
    .Test_en_E_out(Test_enWires[108]),
    .Test_en_W_in(Test_enWires[107]),
    .SC_OUT_BOT(scff_Wires[78]),
    .SC_IN_TOP(scff_Wires[77]),
    .top_width_0_height_0__pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[34]),
    .right_width_0_height_0__pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__30_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_38_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_38_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_38_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_38_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_38_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_38_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_38_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_38_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[33]),
    .ccff_tail(grid_clb_38_ccff_tail[0])
  );


  grid_clb
  grid_clb_5__8_
  (
    .clk_0_S_in(clk_1_wires[80]),
    .prog_clk_0_S_in(prog_clk_1_wires[80]),
    .prog_clk_0_N_out(prog_clk_0_wires[145]),
    .prog_clk_0_E_out(prog_clk_0_wires[143]),
    .prog_clk_0_S_out(prog_clk_0_wires[142]),
    .Test_en_E_out(Test_enWires[122]),
    .Test_en_W_in(Test_enWires[121]),
    .SC_OUT_BOT(scff_Wires[76]),
    .SC_IN_TOP(scff_Wires[75]),
    .top_width_0_height_0__pin_0_(cbx_1__8__4_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__4_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__4_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__4_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__4_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__4_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__4_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__4_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__4_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_5__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__31_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_39_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_39_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_39_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_39_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_39_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_39_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_39_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_39_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[34]),
    .ccff_tail(grid_clb_39_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__1_
  (
    .clk_0_N_in(clk_1_wires[62]),
    .prog_clk_0_N_in(prog_clk_1_wires[62]),
    .prog_clk_0_E_out(prog_clk_0_wires[148]),
    .prog_clk_0_S_out(prog_clk_0_wires[147]),
    .Test_en_E_out(Test_enWires[26]),
    .Test_en_W_in(Test_enWires[25]),
    .SC_OUT_TOP(scff_Wires[95]),
    .SC_IN_BOT(scff_Wires[94]),
    .top_width_0_height_0__pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[35]),
    .right_width_0_height_0__pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__32_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_40_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_40_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_40_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_40_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_40_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_40_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_40_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_40_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_6__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_40_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__2_
  (
    .clk_0_S_in(clk_1_wires[61]),
    .prog_clk_0_S_in(prog_clk_1_wires[61]),
    .prog_clk_0_E_out(prog_clk_0_wires[151]),
    .prog_clk_0_S_out(prog_clk_0_wires[150]),
    .Test_en_E_out(Test_enWires[40]),
    .Test_en_W_in(Test_enWires[39]),
    .SC_OUT_TOP(scff_Wires[97]),
    .SC_IN_BOT(scff_Wires[96]),
    .top_width_0_height_0__pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[36]),
    .right_width_0_height_0__pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__33_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_41_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_41_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_41_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_41_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_41_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_41_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_41_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_41_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[35]),
    .ccff_tail(grid_clb_41_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__3_
  (
    .clk_0_N_in(clk_1_wires[69]),
    .prog_clk_0_N_in(prog_clk_1_wires[69]),
    .prog_clk_0_E_out(prog_clk_0_wires[154]),
    .prog_clk_0_S_out(prog_clk_0_wires[153]),
    .Test_en_E_out(Test_enWires[54]),
    .Test_en_W_in(Test_enWires[53]),
    .SC_OUT_TOP(scff_Wires[99]),
    .SC_IN_BOT(scff_Wires[98]),
    .top_width_0_height_0__pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[37]),
    .right_width_0_height_0__pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__34_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_42_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_42_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_42_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_42_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_42_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_42_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_42_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_42_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[36]),
    .ccff_tail(grid_clb_42_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__4_
  (
    .clk_0_S_in(clk_1_wires[68]),
    .prog_clk_0_S_in(prog_clk_1_wires[68]),
    .prog_clk_0_E_out(prog_clk_0_wires[157]),
    .prog_clk_0_S_out(prog_clk_0_wires[156]),
    .Test_en_E_out(Test_enWires[68]),
    .Test_en_W_in(Test_enWires[67]),
    .SC_OUT_TOP(scff_Wires[101]),
    .SC_IN_BOT(scff_Wires[100]),
    .top_width_0_height_0__pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[38]),
    .right_width_0_height_0__pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__35_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_43_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_43_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_43_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_43_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_43_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_43_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_43_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_43_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[37]),
    .ccff_tail(grid_clb_43_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__5_
  (
    .clk_0_N_in(clk_1_wires[76]),
    .prog_clk_0_N_in(prog_clk_1_wires[76]),
    .prog_clk_0_E_out(prog_clk_0_wires[160]),
    .prog_clk_0_S_out(prog_clk_0_wires[159]),
    .Test_en_E_out(Test_enWires[82]),
    .Test_en_W_in(Test_enWires[81]),
    .SC_OUT_TOP(scff_Wires[103]),
    .SC_IN_BOT(scff_Wires[102]),
    .top_width_0_height_0__pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[39]),
    .right_width_0_height_0__pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__36_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_44_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_44_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_44_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_44_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_44_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_44_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_44_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_44_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[38]),
    .ccff_tail(grid_clb_44_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__6_
  (
    .clk_0_S_in(clk_1_wires[75]),
    .prog_clk_0_S_in(prog_clk_1_wires[75]),
    .prog_clk_0_E_out(prog_clk_0_wires[163]),
    .prog_clk_0_S_out(prog_clk_0_wires[162]),
    .Test_en_E_out(Test_enWires[96]),
    .Test_en_W_in(Test_enWires[95]),
    .SC_OUT_TOP(scff_Wires[105]),
    .SC_IN_BOT(scff_Wires[104]),
    .top_width_0_height_0__pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[40]),
    .right_width_0_height_0__pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__37_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_45_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_45_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_45_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_45_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_45_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_45_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_45_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_45_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[39]),
    .ccff_tail(grid_clb_45_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__7_
  (
    .clk_0_N_in(clk_1_wires[83]),
    .prog_clk_0_N_in(prog_clk_1_wires[83]),
    .prog_clk_0_E_out(prog_clk_0_wires[166]),
    .prog_clk_0_S_out(prog_clk_0_wires[165]),
    .Test_en_E_out(Test_enWires[110]),
    .Test_en_W_in(Test_enWires[109]),
    .SC_OUT_TOP(scff_Wires[107]),
    .SC_IN_BOT(scff_Wires[106]),
    .top_width_0_height_0__pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[41]),
    .right_width_0_height_0__pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__38_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_46_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_46_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_46_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_46_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_46_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_46_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_46_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_46_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[40]),
    .ccff_tail(grid_clb_46_ccff_tail[0])
  );


  grid_clb
  grid_clb_6__8_
  (
    .clk_0_S_in(clk_1_wires[82]),
    .prog_clk_0_S_in(prog_clk_1_wires[82]),
    .prog_clk_0_N_out(prog_clk_0_wires[171]),
    .prog_clk_0_E_out(prog_clk_0_wires[169]),
    .prog_clk_0_S_out(prog_clk_0_wires[168]),
    .Test_en_E_out(Test_enWires[124]),
    .Test_en_W_in(Test_enWires[123]),
    .SC_OUT_TOP(scff_Wires[109]),
    .SC_IN_BOT(scff_Wires[108]),
    .top_width_0_height_0__pin_0_(cbx_1__8__5_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__5_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__5_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__5_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__5_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__5_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__5_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__5_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__5_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_6__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__39_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_47_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_47_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_47_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_47_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_47_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_47_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_47_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_47_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[41]),
    .ccff_tail(grid_clb_47_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__1_
  (
    .clk_0_N_in(clk_1_wires[88]),
    .prog_clk_0_N_in(prog_clk_1_wires[88]),
    .prog_clk_0_E_out(prog_clk_0_wires[174]),
    .prog_clk_0_S_out(prog_clk_0_wires[173]),
    .Test_en_E_out(Test_enWires[28]),
    .Test_en_W_in(Test_enWires[27]),
    .SC_OUT_BOT(scff_Wires[128]),
    .SC_IN_TOP(scff_Wires[126]),
    .top_width_0_height_0__pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[42]),
    .right_width_0_height_0__pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__40_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_48_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_48_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_48_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_48_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_48_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_48_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_48_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_48_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_7__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_48_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__2_
  (
    .clk_0_S_in(clk_1_wires[87]),
    .prog_clk_0_S_in(prog_clk_1_wires[87]),
    .prog_clk_0_E_out(prog_clk_0_wires[177]),
    .prog_clk_0_S_out(prog_clk_0_wires[176]),
    .Test_en_E_out(Test_enWires[42]),
    .Test_en_W_in(Test_enWires[41]),
    .SC_OUT_BOT(scff_Wires[125]),
    .SC_IN_TOP(scff_Wires[124]),
    .top_width_0_height_0__pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[43]),
    .right_width_0_height_0__pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__41_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_49_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_49_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_49_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_49_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_49_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_49_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_49_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_49_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[42]),
    .ccff_tail(grid_clb_49_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__3_
  (
    .clk_0_N_in(clk_1_wires[95]),
    .prog_clk_0_N_in(prog_clk_1_wires[95]),
    .prog_clk_0_E_out(prog_clk_0_wires[180]),
    .prog_clk_0_S_out(prog_clk_0_wires[179]),
    .Test_en_E_out(Test_enWires[56]),
    .Test_en_W_in(Test_enWires[55]),
    .SC_OUT_BOT(scff_Wires[123]),
    .SC_IN_TOP(scff_Wires[122]),
    .top_width_0_height_0__pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[44]),
    .right_width_0_height_0__pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__42_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_50_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_50_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_50_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_50_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_50_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_50_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_50_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_50_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[43]),
    .ccff_tail(grid_clb_50_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__4_
  (
    .clk_0_S_in(clk_1_wires[94]),
    .prog_clk_0_S_in(prog_clk_1_wires[94]),
    .prog_clk_0_E_out(prog_clk_0_wires[183]),
    .prog_clk_0_S_out(prog_clk_0_wires[182]),
    .Test_en_E_out(Test_enWires[70]),
    .Test_en_W_in(Test_enWires[69]),
    .SC_OUT_BOT(scff_Wires[121]),
    .SC_IN_TOP(scff_Wires[120]),
    .top_width_0_height_0__pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[45]),
    .right_width_0_height_0__pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__43_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_51_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_51_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_51_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_51_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_51_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_51_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_51_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_51_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[44]),
    .ccff_tail(grid_clb_51_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__5_
  (
    .clk_0_N_in(clk_1_wires[102]),
    .prog_clk_0_N_in(prog_clk_1_wires[102]),
    .prog_clk_0_E_out(prog_clk_0_wires[186]),
    .prog_clk_0_S_out(prog_clk_0_wires[185]),
    .Test_en_E_out(Test_enWires[84]),
    .Test_en_W_in(Test_enWires[83]),
    .SC_OUT_BOT(scff_Wires[119]),
    .SC_IN_TOP(scff_Wires[118]),
    .top_width_0_height_0__pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[46]),
    .right_width_0_height_0__pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__44_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_52_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_52_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_52_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_52_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_52_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_52_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_52_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_52_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[45]),
    .ccff_tail(grid_clb_52_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__6_
  (
    .clk_0_S_in(clk_1_wires[101]),
    .prog_clk_0_S_in(prog_clk_1_wires[101]),
    .prog_clk_0_E_out(prog_clk_0_wires[189]),
    .prog_clk_0_S_out(prog_clk_0_wires[188]),
    .Test_en_E_out(Test_enWires[98]),
    .Test_en_W_in(Test_enWires[97]),
    .SC_OUT_BOT(scff_Wires[117]),
    .SC_IN_TOP(scff_Wires[116]),
    .top_width_0_height_0__pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[47]),
    .right_width_0_height_0__pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__45_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_53_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_53_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_53_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_53_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_53_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_53_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_53_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_53_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[46]),
    .ccff_tail(grid_clb_53_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__7_
  (
    .clk_0_N_in(clk_1_wires[109]),
    .prog_clk_0_N_in(prog_clk_1_wires[109]),
    .prog_clk_0_E_out(prog_clk_0_wires[192]),
    .prog_clk_0_S_out(prog_clk_0_wires[191]),
    .Test_en_E_out(Test_enWires[112]),
    .Test_en_W_in(Test_enWires[111]),
    .SC_OUT_BOT(scff_Wires[115]),
    .SC_IN_TOP(scff_Wires[114]),
    .top_width_0_height_0__pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[48]),
    .right_width_0_height_0__pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__46_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_54_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_54_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_54_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_54_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_54_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_54_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_54_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_54_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[47]),
    .ccff_tail(grid_clb_54_ccff_tail[0])
  );


  grid_clb
  grid_clb_7__8_
  (
    .clk_0_S_in(clk_1_wires[108]),
    .prog_clk_0_S_in(prog_clk_1_wires[108]),
    .prog_clk_0_N_out(prog_clk_0_wires[197]),
    .prog_clk_0_E_out(prog_clk_0_wires[195]),
    .prog_clk_0_S_out(prog_clk_0_wires[194]),
    .Test_en_E_out(Test_enWires[126]),
    .Test_en_W_in(Test_enWires[125]),
    .SC_OUT_BOT(scff_Wires[113]),
    .SC_IN_TOP(scff_Wires[112]),
    .top_width_0_height_0__pin_0_(cbx_1__8__6_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__6_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__6_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__6_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__6_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__6_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__6_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__6_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__6_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_7__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__47_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_55_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_55_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_55_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_55_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_55_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_55_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_55_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_55_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[48]),
    .ccff_tail(grid_clb_55_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__1_
  (
    .clk_0_N_in(clk_1_wires[90]),
    .prog_clk_0_N_in(prog_clk_1_wires[90]),
    .prog_clk_0_E_out(prog_clk_0_wires[200]),
    .prog_clk_0_S_out(prog_clk_0_wires[199]),
    .Test_en_W_in(Test_enWires[29]),
    .SC_OUT_TOP(scff_Wires[132]),
    .SC_IN_BOT(scff_Wires[131]),
    .top_width_0_height_0__pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[49]),
    .right_width_0_height_0__pin_16_(cby_8__1__0_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__0_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__0_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__0_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__0_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__0_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__0_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__0_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__0_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__0_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__0_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__0_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__0_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__0_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__0_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__0_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__48_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_56_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_56_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_56_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_56_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_56_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_56_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_56_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_56_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(grid_clb_8__1__undriven_bottom_width_0_height_0__pin_50_[0]),
    .ccff_tail(grid_clb_56_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__2_
  (
    .clk_0_S_in(clk_1_wires[89]),
    .prog_clk_0_S_in(prog_clk_1_wires[89]),
    .prog_clk_0_E_out(prog_clk_0_wires[203]),
    .prog_clk_0_S_out(prog_clk_0_wires[202]),
    .Test_en_W_in(Test_enWires[43]),
    .SC_OUT_TOP(scff_Wires[134]),
    .SC_IN_BOT(scff_Wires[133]),
    .top_width_0_height_0__pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[50]),
    .right_width_0_height_0__pin_16_(cby_8__1__1_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__1_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__1_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__1_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__1_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__1_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__1_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__1_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__1_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__1_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__1_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__1_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__1_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__1_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__1_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__1_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__49_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_57_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_57_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_57_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_57_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_57_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_57_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_57_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_57_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[49]),
    .ccff_tail(grid_clb_57_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__3_
  (
    .clk_0_N_in(clk_1_wires[97]),
    .prog_clk_0_N_in(prog_clk_1_wires[97]),
    .prog_clk_0_E_out(prog_clk_0_wires[206]),
    .prog_clk_0_S_out(prog_clk_0_wires[205]),
    .Test_en_W_in(Test_enWires[57]),
    .SC_OUT_TOP(scff_Wires[136]),
    .SC_IN_BOT(scff_Wires[135]),
    .top_width_0_height_0__pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[51]),
    .right_width_0_height_0__pin_16_(cby_8__1__2_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__2_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__2_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__2_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__2_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__2_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__2_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__2_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__2_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__2_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__2_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__2_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__2_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__2_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__2_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__2_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__50_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_58_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_58_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_58_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_58_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_58_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_58_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_58_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_58_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[50]),
    .ccff_tail(grid_clb_58_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__4_
  (
    .clk_0_S_in(clk_1_wires[96]),
    .prog_clk_0_S_in(prog_clk_1_wires[96]),
    .prog_clk_0_E_out(prog_clk_0_wires[209]),
    .prog_clk_0_S_out(prog_clk_0_wires[208]),
    .Test_en_W_in(Test_enWires[71]),
    .SC_OUT_TOP(scff_Wires[138]),
    .SC_IN_BOT(scff_Wires[137]),
    .top_width_0_height_0__pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[52]),
    .right_width_0_height_0__pin_16_(cby_8__1__3_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__3_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__3_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__3_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__3_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__3_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__3_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__3_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__3_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__3_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__3_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__3_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__3_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__3_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__3_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__3_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__51_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_59_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_59_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_59_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_59_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_59_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_59_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_59_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_59_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[51]),
    .ccff_tail(grid_clb_59_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__5_
  (
    .clk_0_N_in(clk_1_wires[104]),
    .prog_clk_0_N_in(prog_clk_1_wires[104]),
    .prog_clk_0_E_out(prog_clk_0_wires[212]),
    .prog_clk_0_S_out(prog_clk_0_wires[211]),
    .Test_en_W_in(Test_enWires[85]),
    .SC_OUT_TOP(scff_Wires[140]),
    .SC_IN_BOT(scff_Wires[139]),
    .top_width_0_height_0__pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[53]),
    .right_width_0_height_0__pin_16_(cby_8__1__4_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__4_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__4_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__4_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__4_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__4_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__4_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__4_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__4_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__4_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__4_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__4_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__4_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__4_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__4_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__4_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__52_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_60_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_60_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_60_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_60_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_60_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_60_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_60_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_60_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[52]),
    .ccff_tail(grid_clb_60_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__6_
  (
    .clk_0_S_in(clk_1_wires[103]),
    .prog_clk_0_S_in(prog_clk_1_wires[103]),
    .prog_clk_0_E_out(prog_clk_0_wires[215]),
    .prog_clk_0_S_out(prog_clk_0_wires[214]),
    .Test_en_W_in(Test_enWires[99]),
    .SC_OUT_TOP(scff_Wires[142]),
    .SC_IN_BOT(scff_Wires[141]),
    .top_width_0_height_0__pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[54]),
    .right_width_0_height_0__pin_16_(cby_8__1__5_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__5_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__5_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__5_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__5_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__5_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__5_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__5_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__5_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__5_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__5_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__5_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__5_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__5_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__5_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__5_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__53_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_61_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_61_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_61_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_61_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_61_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_61_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_61_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_61_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[53]),
    .ccff_tail(grid_clb_61_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__7_
  (
    .clk_0_N_in(clk_1_wires[111]),
    .prog_clk_0_N_in(prog_clk_1_wires[111]),
    .prog_clk_0_E_out(prog_clk_0_wires[218]),
    .prog_clk_0_S_out(prog_clk_0_wires[217]),
    .Test_en_W_in(Test_enWires[113]),
    .SC_OUT_TOP(scff_Wires[144]),
    .SC_IN_BOT(scff_Wires[143]),
    .top_width_0_height_0__pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(regout_feedthrough_wires[55]),
    .right_width_0_height_0__pin_16_(cby_8__1__6_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__6_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__6_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__6_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__6_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__6_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__6_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__6_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__6_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__6_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__6_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__6_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__6_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__6_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__6_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__6_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__54_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_62_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_62_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_62_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_62_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_62_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_62_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_62_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_62_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[54]),
    .ccff_tail(grid_clb_62_ccff_tail[0])
  );


  grid_clb
  grid_clb_8__8_
  (
    .clk_0_S_in(clk_1_wires[110]),
    .prog_clk_0_S_in(prog_clk_1_wires[110]),
    .prog_clk_0_N_out(prog_clk_0_wires[223]),
    .prog_clk_0_E_out(prog_clk_0_wires[221]),
    .prog_clk_0_S_out(prog_clk_0_wires[220]),
    .Test_en_W_in(Test_enWires[127]),
    .SC_OUT_TOP(scff_Wires[146]),
    .SC_IN_BOT(scff_Wires[145]),
    .top_width_0_height_0__pin_0_(cbx_1__8__7_bottom_grid_pin_0_[0]),
    .top_width_0_height_0__pin_1_(cbx_1__8__7_bottom_grid_pin_1_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__8__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_3_(cbx_1__8__7_bottom_grid_pin_3_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__8__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_5_(cbx_1__8__7_bottom_grid_pin_5_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__8__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_7_(cbx_1__8__7_bottom_grid_pin_7_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__8__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_9_(cbx_1__8__7_bottom_grid_pin_9_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__8__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_11_(cbx_1__8__7_bottom_grid_pin_11_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__8__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_13_(cbx_1__8__7_bottom_grid_pin_13_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__8__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_15_(cbx_1__8__7_bottom_grid_pin_15_[0]),
    .top_width_0_height_0__pin_32_(grid_clb_8__8__undriven_top_width_0_height_0__pin_32_[0]),
    .right_width_0_height_0__pin_16_(cby_8__1__7_left_grid_pin_16_[0]),
    .right_width_0_height_0__pin_17_(cby_8__1__7_left_grid_pin_17_[0]),
    .right_width_0_height_0__pin_18_(cby_8__1__7_left_grid_pin_18_[0]),
    .right_width_0_height_0__pin_19_(cby_8__1__7_left_grid_pin_19_[0]),
    .right_width_0_height_0__pin_20_(cby_8__1__7_left_grid_pin_20_[0]),
    .right_width_0_height_0__pin_21_(cby_8__1__7_left_grid_pin_21_[0]),
    .right_width_0_height_0__pin_22_(cby_8__1__7_left_grid_pin_22_[0]),
    .right_width_0_height_0__pin_23_(cby_8__1__7_left_grid_pin_23_[0]),
    .right_width_0_height_0__pin_24_(cby_8__1__7_left_grid_pin_24_[0]),
    .right_width_0_height_0__pin_25_(cby_8__1__7_left_grid_pin_25_[0]),
    .right_width_0_height_0__pin_26_(cby_8__1__7_left_grid_pin_26_[0]),
    .right_width_0_height_0__pin_27_(cby_8__1__7_left_grid_pin_27_[0]),
    .right_width_0_height_0__pin_28_(cby_8__1__7_left_grid_pin_28_[0]),
    .right_width_0_height_0__pin_29_(cby_8__1__7_left_grid_pin_29_[0]),
    .right_width_0_height_0__pin_30_(cby_8__1__7_left_grid_pin_30_[0]),
    .right_width_0_height_0__pin_31_(cby_8__1__7_left_grid_pin_31_[0]),
    .ccff_head(cby_1__1__55_ccff_tail[0]),
    .top_width_0_height_0__pin_34_upper(grid_clb_63_top_width_0_height_0__pin_34_upper[0]),
    .top_width_0_height_0__pin_34_lower(grid_clb_63_top_width_0_height_0__pin_34_lower[0]),
    .top_width_0_height_0__pin_35_upper(grid_clb_63_top_width_0_height_0__pin_35_upper[0]),
    .top_width_0_height_0__pin_35_lower(grid_clb_63_top_width_0_height_0__pin_35_lower[0]),
    .top_width_0_height_0__pin_36_upper(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
    .top_width_0_height_0__pin_36_lower(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
    .top_width_0_height_0__pin_37_upper(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
    .top_width_0_height_0__pin_37_lower(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
    .top_width_0_height_0__pin_38_upper(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
    .top_width_0_height_0__pin_38_lower(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
    .top_width_0_height_0__pin_39_upper(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
    .top_width_0_height_0__pin_39_lower(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
    .top_width_0_height_0__pin_40_upper(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
    .top_width_0_height_0__pin_40_lower(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
    .top_width_0_height_0__pin_41_upper(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
    .top_width_0_height_0__pin_41_lower(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
    .right_width_0_height_0__pin_42_upper(grid_clb_63_right_width_0_height_0__pin_42_upper[0]),
    .right_width_0_height_0__pin_42_lower(grid_clb_63_right_width_0_height_0__pin_42_lower[0]),
    .right_width_0_height_0__pin_43_upper(grid_clb_63_right_width_0_height_0__pin_43_upper[0]),
    .right_width_0_height_0__pin_43_lower(grid_clb_63_right_width_0_height_0__pin_43_lower[0]),
    .right_width_0_height_0__pin_44_upper(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
    .right_width_0_height_0__pin_44_lower(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
    .right_width_0_height_0__pin_45_upper(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
    .right_width_0_height_0__pin_45_lower(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
    .right_width_0_height_0__pin_46_upper(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
    .right_width_0_height_0__pin_46_lower(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
    .right_width_0_height_0__pin_47_upper(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
    .right_width_0_height_0__pin_47_lower(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
    .right_width_0_height_0__pin_48_upper(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
    .right_width_0_height_0__pin_48_lower(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
    .right_width_0_height_0__pin_49_upper(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
    .right_width_0_height_0__pin_49_lower(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
    .bottom_width_0_height_0__pin_50_(regin_feedthrough_wires[55]),
    .ccff_tail(grid_clb_63_ccff_tail[0])
  );


  sb_0__0_
  sb_0__0_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[5]),
    .chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_upper[0]),
    .ccff_head(grid_io_bottom_7_ccff_tail[0]),
    .chany_top_out(sb_0__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
    .ccff_tail(ccff_tail[0])
  );


  sb_0__1_
  sb_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[4]),
    .chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__0_ccff_tail[0]),
    .chany_top_out(sb_0__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__0_ccff_tail[0])
  );


  sb_0__1_
  sb_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[10]),
    .chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__1_ccff_tail[0]),
    .chany_top_out(sb_0__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__1_ccff_tail[0])
  );


  sb_0__1_
  sb_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[15]),
    .chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__2_ccff_tail[0]),
    .chany_top_out(sb_0__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__2_ccff_tail[0])
  );


  sb_0__1_
  sb_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[20]),
    .chany_top_in(cby_0__1__4_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__3_ccff_tail[0]),
    .chany_top_out(sb_0__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__3_ccff_tail[0])
  );


  sb_0__1_
  sb_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[25]),
    .chany_top_in(cby_0__1__5_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__4_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__4_ccff_tail[0]),
    .chany_top_out(sb_0__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__4_ccff_tail[0])
  );


  sb_0__1_
  sb_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[30]),
    .chany_top_in(cby_0__1__6_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__5_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__5_ccff_tail[0]),
    .chany_top_out(sb_0__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__5_ccff_tail[0])
  );


  sb_0__1_
  sb_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[35]),
    .chany_top_in(cby_0__1__7_chany_bottom_out[0:19]),
    .top_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
    .chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__6_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(cbx_1__1__6_ccff_tail[0]),
    .chany_top_out(sb_0__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_0__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__1__6_ccff_tail[0])
  );


  sb_0__2_
  sb_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[42]),
    .SC_OUT_BOT(scff_Wires[0]),
    .SC_IN_TOP(sc_head),
    .chanx_right_in(cbx_1__8__0_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_0__1__7_chany_top_out[0:19]),
    .bottom_left_grid_pin_1_(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
    .ccff_head(grid_io_top_0_ccff_tail[0]),
    .chanx_right_out(sb_0__8__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_0__8__0_chany_bottom_out[0:19]),
    .ccff_tail(sb_0__8__0_ccff_tail[0])
  );


  sb_1__0_
  sb_1__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[2]),
    .SC_OUT_TOP(scff_Wires[19]),
    .SC_IN_TOP(scff_Wires[18]),
    .chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_7_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_7_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_7_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_7_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_7_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_7_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_7_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_7_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_6_ccff_tail[0]),
    .chany_top_out(sb_1__0__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__0_ccff_tail[0])
  );


  sb_1__0_
  sb_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[45]),
    .chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_6_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_6_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_6_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_6_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_6_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_6_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_6_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_6_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_5_ccff_tail[0]),
    .chany_top_out(sb_1__0__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__1_ccff_tail[0])
  );


  sb_1__0_
  sb_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[71]),
    .SC_OUT_TOP(scff_Wires[56]),
    .SC_IN_TOP(scff_Wires[55]),
    .chany_top_in(cby_1__1__16_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_5_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_5_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_5_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_5_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_5_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_5_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_5_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_5_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_4_ccff_tail[0]),
    .chany_top_out(sb_1__0__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__2_ccff_tail[0])
  );


  sb_1__0_
  sb_4__0_
  (
    .clk_3_N_out(clk_3_wires[28]),
    .clk_3_S_in(clk),
    .prog_clk_3_N_out(prog_clk_3_wires[28]),
    .prog_clk_3_S_in(prog_clk),
    .prog_clk_0_N_in(prog_clk_0_wires[97]),
    .Test_en_N_out(Test_enWires[1]),
    .Test_en_S_in(Test_en),
    .chany_top_in(cby_1__1__24_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__4_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_4_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_4_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_4_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_4_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_4_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_4_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_4_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_4_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_3_ccff_tail[0]),
    .chany_top_out(sb_1__0__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__3_ccff_tail[0])
  );


  sb_1__0_
  sb_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[123]),
    .SC_OUT_TOP(scff_Wires[93]),
    .SC_IN_TOP(scff_Wires[92]),
    .chany_top_in(cby_1__1__32_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__5_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__4_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_3_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_3_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_3_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_3_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_3_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_3_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_3_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_3_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_2_ccff_tail[0]),
    .chany_top_out(sb_1__0__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__4_ccff_tail[0])
  );


  sb_1__0_
  sb_6__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[149]),
    .chany_top_in(cby_1__1__40_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__6_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__5_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_2_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_2_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_2_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_2_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_2_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_2_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_2_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_2_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_1_ccff_tail[0]),
    .chany_top_out(sb_1__0__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__5_ccff_tail[0])
  );


  sb_1__0_
  sb_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[175]),
    .SC_OUT_TOP(scff_Wires[130]),
    .SC_IN_TOP(scff_Wires[129]),
    .chany_top_in(cby_1__1__48_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__0__7_chanx_left_out[0:19]),
    .right_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_upper[0]),
    .right_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_upper[0]),
    .right_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_upper[0]),
    .right_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_upper[0]),
    .right_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_upper[0]),
    .right_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_upper[0]),
    .right_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_upper[0]),
    .right_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_upper[0]),
    .chanx_left_in(cbx_1__0__6_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_1_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_1_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_1_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_1_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_1_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_1_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_1_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_1_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_bottom_0_ccff_tail[0]),
    .chany_top_out(sb_1__0__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_left_out(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__0__6_ccff_tail[0])
  );


  sb_1__1_
  sb_1__1_
  (
    .clk_1_N_in(clk_2_wires[8]),
    .clk_1_W_out(clk_1_wires[2]),
    .clk_1_E_out(clk_1_wires[1]),
    .prog_clk_1_N_in(prog_clk_2_wires[8]),
    .prog_clk_1_W_out(prog_clk_1_wires[2]),
    .prog_clk_1_E_out(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[8]),
    .chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_0_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_0_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_0_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_0_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_0_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_0_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_0_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_0_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_0_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_0_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_0_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_0_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_0_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_0_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_0_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_0_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__7_ccff_tail[0]),
    .chany_top_out(sb_1__1__0_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__0_ccff_tail[0])
  );


  sb_1__1_
  sb_1__2_
  (
    .clk_2_S_out(clk_2_wires[7]),
    .clk_2_N_out(clk_2_wires[5]),
    .clk_2_E_in(clk_2_wires[4]),
    .prog_clk_2_S_out(prog_clk_2_wires[7]),
    .prog_clk_2_N_out(prog_clk_2_wires[5]),
    .prog_clk_2_E_in(prog_clk_2_wires[4]),
    .prog_clk_0_N_in(prog_clk_0_wires[13]),
    .chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_1_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_1_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_1_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_1_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_1_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_1_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_1_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_1_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_1_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_1_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_1_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_1_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_1_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_1_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_1_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_1_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__8_ccff_tail[0]),
    .chany_top_out(sb_1__1__1_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__1_ccff_tail[0])
  );


  sb_1__1_
  sb_1__3_
  (
    .clk_1_S_in(clk_2_wires[6]),
    .clk_1_W_out(clk_1_wires[9]),
    .clk_1_E_out(clk_1_wires[8]),
    .prog_clk_1_S_in(prog_clk_2_wires[6]),
    .prog_clk_1_W_out(prog_clk_1_wires[9]),
    .prog_clk_1_E_out(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[18]),
    .chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_2_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_2_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_2_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_2_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_2_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_2_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_2_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_2_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_2_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_2_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_2_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_2_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_2_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_2_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_2_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_2_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__9_ccff_tail[0]),
    .chany_top_out(sb_1__1__2_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__2_ccff_tail[0])
  );


  sb_1__1_
  sb_1__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[23]),
    .chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_3_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_3_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_3_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_3_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_3_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_3_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_3_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_3_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_3_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_3_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_3_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_3_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_3_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_3_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_3_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_3_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__10_ccff_tail[0]),
    .chany_top_out(sb_1__1__3_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__3_ccff_tail[0])
  );


  sb_1__1_
  sb_1__5_
  (
    .clk_1_N_in(clk_2_wires[21]),
    .clk_1_W_out(clk_1_wires[16]),
    .clk_1_E_out(clk_1_wires[15]),
    .prog_clk_1_N_in(prog_clk_2_wires[21]),
    .prog_clk_1_W_out(prog_clk_1_wires[16]),
    .prog_clk_1_E_out(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[28]),
    .chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_4_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_4_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_4_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_4_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_4_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_4_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_4_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_4_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_4_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_4_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_4_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_4_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_4_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_4_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_4_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_4_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__11_ccff_tail[0]),
    .chany_top_out(sb_1__1__4_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__4_ccff_tail[0])
  );


  sb_1__1_
  sb_1__6_
  (
    .clk_2_S_out(clk_2_wires[20]),
    .clk_2_N_out(clk_2_wires[18]),
    .clk_2_E_in(clk_2_wires[17]),
    .prog_clk_2_S_out(prog_clk_2_wires[20]),
    .prog_clk_2_N_out(prog_clk_2_wires[18]),
    .prog_clk_2_E_in(prog_clk_2_wires[17]),
    .prog_clk_0_N_in(prog_clk_0_wires[33]),
    .chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__12_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_5_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_5_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_5_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_5_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_5_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_5_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_5_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_5_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_5_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_5_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_5_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_5_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_5_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_5_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_5_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_5_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__12_ccff_tail[0]),
    .chany_top_out(sb_1__1__5_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__5_ccff_tail[0])
  );


  sb_1__1_
  sb_1__7_
  (
    .clk_1_S_in(clk_2_wires[19]),
    .clk_1_W_out(clk_1_wires[23]),
    .clk_1_E_out(clk_1_wires[22]),
    .prog_clk_1_S_in(prog_clk_2_wires[19]),
    .prog_clk_1_W_out(prog_clk_1_wires[23]),
    .prog_clk_1_E_out(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[38]),
    .chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__13_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_6_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_6_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_6_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_6_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_6_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_6_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_6_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_6_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_6_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_6_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_6_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_6_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_6_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_6_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_6_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_6_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__13_ccff_tail[0]),
    .chany_top_out(sb_1__1__6_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__6_ccff_tail[0])
  );


  sb_1__1_
  sb_2__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[48]),
    .chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__14_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_8_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_8_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_8_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_8_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_8_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_8_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_8_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_8_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_8_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_8_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_8_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_8_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_8_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_8_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_8_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_8_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__14_ccff_tail[0]),
    .chany_top_out(sb_1__1__7_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__7_ccff_tail[0])
  );


  sb_1__1_
  sb_2__2_
  (
    .clk_2_N_in(clk_3_wires[17]),
    .clk_2_W_out(clk_2_wires[3]),
    .clk_2_E_out(clk_2_wires[1]),
    .prog_clk_2_N_in(prog_clk_3_wires[17]),
    .prog_clk_2_W_out(prog_clk_2_wires[3]),
    .prog_clk_2_E_out(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[51]),
    .chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__15_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_9_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_9_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_9_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_9_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_9_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_9_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_9_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_9_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_9_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_9_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_9_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_9_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_9_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_9_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_9_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_9_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__15_ccff_tail[0]),
    .chany_top_out(sb_1__1__8_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__8_ccff_tail[0])
  );


  sb_1__1_
  sb_2__3_
  (
    .clk_3_S_out(clk_3_wires[16]),
    .clk_3_N_in(clk_3_wires[13]),
    .prog_clk_3_S_out(prog_clk_3_wires[16]),
    .prog_clk_3_N_in(prog_clk_3_wires[13]),
    .prog_clk_0_N_in(prog_clk_0_wires[54]),
    .chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__16_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_10_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_10_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_10_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_10_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_10_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_10_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_10_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_10_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_10_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_10_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_10_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_10_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_10_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_10_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_10_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_10_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__16_ccff_tail[0]),
    .chany_top_out(sb_1__1__9_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__9_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__9_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__9_ccff_tail[0])
  );


  sb_1__1_
  sb_2__4_
  (
    .clk_3_S_out(clk_3_wires[12]),
    .clk_3_N_out(clk_3_wires[10]),
    .clk_3_E_in(clk_3_wires[9]),
    .prog_clk_3_S_out(prog_clk_3_wires[12]),
    .prog_clk_3_N_out(prog_clk_3_wires[10]),
    .prog_clk_3_E_in(prog_clk_3_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[57]),
    .chany_top_in(cby_1__1__12_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__17_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_11_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_11_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_11_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_11_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_11_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_11_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_11_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_11_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_11_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_11_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_11_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_11_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_11_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_11_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_11_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_11_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__17_ccff_tail[0]),
    .chany_top_out(sb_1__1__10_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__10_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__10_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__10_ccff_tail[0])
  );


  sb_1__1_
  sb_2__5_
  (
    .clk_3_N_out(clk_3_wires[14]),
    .clk_3_S_in(clk_3_wires[11]),
    .prog_clk_3_N_out(prog_clk_3_wires[14]),
    .prog_clk_3_S_in(prog_clk_3_wires[11]),
    .prog_clk_0_N_in(prog_clk_0_wires[60]),
    .chany_top_in(cby_1__1__13_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__18_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__12_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_12_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_12_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_12_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_12_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_12_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_12_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_12_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_12_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_12_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_12_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_12_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_12_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_12_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_12_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_12_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_12_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__18_ccff_tail[0]),
    .chany_top_out(sb_1__1__11_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__11_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__11_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__11_ccff_tail[0])
  );


  sb_1__1_
  sb_2__6_
  (
    .clk_2_S_in(clk_3_wires[15]),
    .clk_2_W_out(clk_2_wires[16]),
    .clk_2_E_out(clk_2_wires[14]),
    .prog_clk_2_S_in(prog_clk_3_wires[15]),
    .prog_clk_2_W_out(prog_clk_2_wires[16]),
    .prog_clk_2_E_out(prog_clk_2_wires[14]),
    .prog_clk_0_N_in(prog_clk_0_wires[63]),
    .chany_top_in(cby_1__1__14_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__19_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__13_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_13_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_13_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_13_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_13_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_13_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_13_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_13_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_13_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__12_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_13_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_13_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_13_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_13_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_13_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_13_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_13_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_13_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__19_ccff_tail[0]),
    .chany_top_out(sb_1__1__12_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__12_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__12_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__12_ccff_tail[0])
  );


  sb_1__1_
  sb_2__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[66]),
    .chany_top_in(cby_1__1__15_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__20_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__14_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_14_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_14_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_14_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_14_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_14_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_14_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_14_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_14_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__13_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_14_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_14_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_14_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_14_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_14_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_14_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_14_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_14_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__20_ccff_tail[0]),
    .chany_top_out(sb_1__1__13_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__13_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__13_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__13_ccff_tail[0])
  );


  sb_1__1_
  sb_3__1_
  (
    .clk_1_N_in(clk_2_wires[12]),
    .clk_1_W_out(clk_1_wires[30]),
    .clk_1_E_out(clk_1_wires[29]),
    .prog_clk_1_N_in(prog_clk_2_wires[12]),
    .prog_clk_1_W_out(prog_clk_1_wires[30]),
    .prog_clk_1_E_out(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[74]),
    .chany_top_in(cby_1__1__17_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__21_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__16_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_16_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_16_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_16_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_16_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_16_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_16_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_16_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_16_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__14_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_16_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_16_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_16_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_16_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_16_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_16_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_16_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_16_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__21_ccff_tail[0]),
    .chany_top_out(sb_1__1__14_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__14_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__14_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__14_ccff_tail[0])
  );


  sb_1__1_
  sb_3__2_
  (
    .clk_2_S_out(clk_2_wires[11]),
    .clk_2_N_out(clk_2_wires[9]),
    .clk_2_W_in(clk_2_wires[2]),
    .prog_clk_2_S_out(prog_clk_2_wires[11]),
    .prog_clk_2_N_out(prog_clk_2_wires[9]),
    .prog_clk_2_W_in(prog_clk_2_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[77]),
    .chany_top_in(cby_1__1__18_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__22_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__17_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_17_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_17_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_17_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_17_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_17_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_17_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_17_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_17_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__15_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_17_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_17_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_17_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_17_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_17_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_17_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_17_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_17_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__22_ccff_tail[0]),
    .chany_top_out(sb_1__1__15_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__15_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__15_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__15_ccff_tail[0])
  );


  sb_1__1_
  sb_3__3_
  (
    .clk_1_S_in(clk_2_wires[10]),
    .clk_1_W_out(clk_1_wires[37]),
    .clk_1_E_out(clk_1_wires[36]),
    .prog_clk_1_S_in(prog_clk_2_wires[10]),
    .prog_clk_1_W_out(prog_clk_1_wires[37]),
    .prog_clk_1_E_out(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[80]),
    .chany_top_in(cby_1__1__19_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__23_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__18_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_18_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_18_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_18_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_18_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_18_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_18_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_18_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_18_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__16_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_18_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_18_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_18_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_18_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_18_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_18_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_18_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_18_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__23_ccff_tail[0]),
    .chany_top_out(sb_1__1__16_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__16_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__16_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__16_ccff_tail[0])
  );


  sb_1__1_
  sb_3__4_
  (
    .clk_3_W_out(clk_3_wires[8]),
    .clk_3_E_in(clk_3_wires[4]),
    .prog_clk_3_W_out(prog_clk_3_wires[8]),
    .prog_clk_3_E_in(prog_clk_3_wires[4]),
    .prog_clk_0_N_in(prog_clk_0_wires[83]),
    .chany_top_in(cby_1__1__20_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__24_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__19_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_19_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_19_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_19_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_19_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_19_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_19_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_19_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_19_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__17_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_19_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_19_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_19_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_19_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_19_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_19_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_19_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_19_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__24_ccff_tail[0]),
    .chany_top_out(sb_1__1__17_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__17_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__17_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__17_ccff_tail[0])
  );


  sb_1__1_
  sb_3__5_
  (
    .clk_1_N_in(clk_2_wires[25]),
    .clk_1_W_out(clk_1_wires[44]),
    .clk_1_E_out(clk_1_wires[43]),
    .prog_clk_1_N_in(prog_clk_2_wires[25]),
    .prog_clk_1_W_out(prog_clk_1_wires[44]),
    .prog_clk_1_E_out(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[86]),
    .chany_top_in(cby_1__1__21_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__25_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__20_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_20_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_20_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_20_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_20_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_20_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_20_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_20_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_20_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__18_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_20_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_20_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_20_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_20_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_20_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_20_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_20_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_20_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__25_ccff_tail[0]),
    .chany_top_out(sb_1__1__18_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__18_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__18_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__18_ccff_tail[0])
  );


  sb_1__1_
  sb_3__6_
  (
    .clk_2_S_out(clk_2_wires[24]),
    .clk_2_N_out(clk_2_wires[22]),
    .clk_2_W_in(clk_2_wires[15]),
    .prog_clk_2_S_out(prog_clk_2_wires[24]),
    .prog_clk_2_N_out(prog_clk_2_wires[22]),
    .prog_clk_2_W_in(prog_clk_2_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[89]),
    .chany_top_in(cby_1__1__22_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__26_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__21_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_21_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_21_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_21_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_21_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_21_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_21_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_21_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_21_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__19_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_21_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_21_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_21_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_21_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_21_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_21_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_21_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_21_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__26_ccff_tail[0]),
    .chany_top_out(sb_1__1__19_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__19_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__19_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__19_ccff_tail[0])
  );


  sb_1__1_
  sb_3__7_
  (
    .clk_1_S_in(clk_2_wires[23]),
    .clk_1_W_out(clk_1_wires[51]),
    .clk_1_E_out(clk_1_wires[50]),
    .prog_clk_1_S_in(prog_clk_2_wires[23]),
    .prog_clk_1_W_out(prog_clk_1_wires[51]),
    .prog_clk_1_E_out(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[92]),
    .chany_top_in(cby_1__1__23_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__27_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__22_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_22_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_22_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_22_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_22_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_22_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_22_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_22_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_22_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__20_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_22_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_22_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_22_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_22_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_22_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_22_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_22_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_22_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__27_ccff_tail[0]),
    .chany_top_out(sb_1__1__20_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__20_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__20_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__20_ccff_tail[0])
  );


  sb_1__1_
  sb_4__1_
  (
    .clk_3_N_out(clk_3_wires[30]),
    .clk_3_S_in(clk_3_wires[27]),
    .prog_clk_3_N_out(prog_clk_3_wires[30]),
    .prog_clk_3_S_in(prog_clk_3_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[100]),
    .Test_en_N_out(Test_enWires[3]),
    .Test_en_S_in(Test_enWires[2]),
    .chany_top_in(cby_1__1__25_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__28_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__24_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_24_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_24_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_24_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_24_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_24_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_24_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_24_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_24_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__21_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_24_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_24_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_24_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_24_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_24_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_24_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_24_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_24_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__28_ccff_tail[0]),
    .chany_top_out(sb_1__1__21_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__21_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__21_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__21_ccff_tail[0])
  );


  sb_1__1_
  sb_4__2_
  (
    .clk_3_N_out(clk_3_wires[32]),
    .clk_3_S_in(clk_3_wires[29]),
    .prog_clk_3_N_out(prog_clk_3_wires[32]),
    .prog_clk_3_S_in(prog_clk_3_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[103]),
    .Test_en_N_out(Test_enWires[5]),
    .Test_en_S_in(Test_enWires[4]),
    .chany_top_in(cby_1__1__26_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__29_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__25_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_25_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_25_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_25_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_25_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_25_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_25_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_25_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_25_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__22_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_25_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_25_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_25_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_25_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_25_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_25_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_25_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_25_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__29_ccff_tail[0]),
    .chany_top_out(sb_1__1__22_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__22_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__22_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__22_ccff_tail[0])
  );


  sb_1__1_
  sb_4__3_
  (
    .clk_3_N_out(clk_3_wires[34]),
    .clk_3_S_in(clk_3_wires[31]),
    .prog_clk_3_N_out(prog_clk_3_wires[34]),
    .prog_clk_3_S_in(prog_clk_3_wires[31]),
    .prog_clk_0_N_in(prog_clk_0_wires[106]),
    .Test_en_N_out(Test_enWires[7]),
    .Test_en_S_in(Test_enWires[6]),
    .chany_top_in(cby_1__1__27_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__30_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__26_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_26_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_26_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_26_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_26_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_26_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_26_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_26_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_26_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__23_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_26_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_26_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_26_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_26_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_26_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_26_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_26_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_26_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__30_ccff_tail[0]),
    .chany_top_out(sb_1__1__23_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__23_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__23_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__23_ccff_tail[0])
  );


  sb_1__1_
  sb_4__4_
  (
    .clk_3_S_in(clk_3_wires[33]),
    .clk_3_W_out(clk_3_wires[3]),
    .clk_3_E_out(clk_3_wires[1]),
    .prog_clk_3_S_in(prog_clk_3_wires[33]),
    .prog_clk_3_W_out(prog_clk_3_wires[3]),
    .prog_clk_3_E_out(prog_clk_3_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[109]),
    .Test_en_N_out(Test_enWires[9]),
    .Test_en_S_in(Test_enWires[8]),
    .chany_top_in(cby_1__1__28_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__31_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__27_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_27_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_27_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_27_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_27_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_27_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_27_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_27_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_27_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__24_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_27_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_27_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_27_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_27_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_27_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_27_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_27_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_27_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__31_ccff_tail[0]),
    .chany_top_out(sb_1__1__24_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__24_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__24_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__24_ccff_tail[0])
  );


  sb_1__1_
  sb_4__5_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[112]),
    .Test_en_N_out(Test_enWires[11]),
    .Test_en_S_in(Test_enWires[10]),
    .chany_top_in(cby_1__1__29_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__32_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__28_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_28_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_28_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_28_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_28_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_28_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_28_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_28_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_28_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__25_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_28_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_28_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_28_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_28_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_28_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_28_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_28_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_28_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__32_ccff_tail[0]),
    .chany_top_out(sb_1__1__25_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__25_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__25_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__25_ccff_tail[0])
  );


  sb_1__1_
  sb_4__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[115]),
    .Test_en_N_out(Test_enWires[13]),
    .Test_en_S_in(Test_enWires[12]),
    .chany_top_in(cby_1__1__30_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__33_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__29_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_29_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_29_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_29_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_29_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_29_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_29_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_29_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_29_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__26_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_29_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_29_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_29_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_29_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_29_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_29_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_29_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_29_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__33_ccff_tail[0]),
    .chany_top_out(sb_1__1__26_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__26_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__26_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__26_ccff_tail[0])
  );


  sb_1__1_
  sb_4__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[118]),
    .Test_en_N_out(Test_enWires[15]),
    .Test_en_S_in(Test_enWires[14]),
    .chany_top_in(cby_1__1__31_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__34_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__30_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_30_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_30_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_30_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_30_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_30_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_30_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_30_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_30_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__27_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_30_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_30_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_30_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_30_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_30_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_30_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_30_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_30_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__34_ccff_tail[0]),
    .chany_top_out(sb_1__1__27_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__27_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__27_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__27_ccff_tail[0])
  );


  sb_1__1_
  sb_5__1_
  (
    .clk_1_N_in(clk_2_wires[34]),
    .clk_1_W_out(clk_1_wires[58]),
    .clk_1_E_out(clk_1_wires[57]),
    .prog_clk_1_N_in(prog_clk_2_wires[34]),
    .prog_clk_1_W_out(prog_clk_1_wires[58]),
    .prog_clk_1_E_out(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[126]),
    .chany_top_in(cby_1__1__33_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__35_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__32_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_32_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_32_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_32_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_32_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_32_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_32_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_32_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_32_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__28_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_32_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_32_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_32_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_32_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_32_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_32_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_32_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_32_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__35_ccff_tail[0]),
    .chany_top_out(sb_1__1__28_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__28_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__28_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__28_ccff_tail[0])
  );


  sb_1__1_
  sb_5__2_
  (
    .clk_2_S_out(clk_2_wires[33]),
    .clk_2_N_out(clk_2_wires[31]),
    .clk_2_E_in(clk_2_wires[30]),
    .prog_clk_2_S_out(prog_clk_2_wires[33]),
    .prog_clk_2_N_out(prog_clk_2_wires[31]),
    .prog_clk_2_E_in(prog_clk_2_wires[30]),
    .prog_clk_0_N_in(prog_clk_0_wires[129]),
    .chany_top_in(cby_1__1__34_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__36_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__33_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_33_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_33_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_33_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_33_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_33_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_33_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_33_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_33_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__29_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_33_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_33_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_33_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_33_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_33_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_33_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_33_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_33_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__36_ccff_tail[0]),
    .chany_top_out(sb_1__1__29_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__29_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__29_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__29_ccff_tail[0])
  );


  sb_1__1_
  sb_5__3_
  (
    .clk_1_S_in(clk_2_wires[32]),
    .clk_1_W_out(clk_1_wires[65]),
    .clk_1_E_out(clk_1_wires[64]),
    .prog_clk_1_S_in(prog_clk_2_wires[32]),
    .prog_clk_1_W_out(prog_clk_1_wires[65]),
    .prog_clk_1_E_out(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[132]),
    .chany_top_in(cby_1__1__35_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__37_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__34_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_34_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_34_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_34_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_34_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_34_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_34_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_34_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_34_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__30_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_34_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_34_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_34_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_34_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_34_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_34_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_34_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_34_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__37_ccff_tail[0]),
    .chany_top_out(sb_1__1__30_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__30_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__30_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__30_ccff_tail[0])
  );


  sb_1__1_
  sb_5__4_
  (
    .clk_3_E_out(clk_3_wires[6]),
    .clk_3_W_in(clk_3_wires[2]),
    .prog_clk_3_E_out(prog_clk_3_wires[6]),
    .prog_clk_3_W_in(prog_clk_3_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[135]),
    .chany_top_in(cby_1__1__36_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__38_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__35_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_35_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_35_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_35_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_35_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_35_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_35_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_35_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_35_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__31_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_35_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_35_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_35_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_35_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_35_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_35_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_35_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_35_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__38_ccff_tail[0]),
    .chany_top_out(sb_1__1__31_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__31_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__31_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__31_ccff_tail[0])
  );


  sb_1__1_
  sb_5__5_
  (
    .clk_1_N_in(clk_2_wires[47]),
    .clk_1_W_out(clk_1_wires[72]),
    .clk_1_E_out(clk_1_wires[71]),
    .prog_clk_1_N_in(prog_clk_2_wires[47]),
    .prog_clk_1_W_out(prog_clk_1_wires[72]),
    .prog_clk_1_E_out(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[138]),
    .chany_top_in(cby_1__1__37_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__39_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__36_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_36_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_36_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_36_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_36_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_36_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_36_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_36_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_36_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__32_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_36_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_36_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_36_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_36_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_36_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_36_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_36_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_36_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__39_ccff_tail[0]),
    .chany_top_out(sb_1__1__32_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__32_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__32_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__32_ccff_tail[0])
  );


  sb_1__1_
  sb_5__6_
  (
    .clk_2_S_out(clk_2_wires[46]),
    .clk_2_N_out(clk_2_wires[44]),
    .clk_2_E_in(clk_2_wires[43]),
    .prog_clk_2_S_out(prog_clk_2_wires[46]),
    .prog_clk_2_N_out(prog_clk_2_wires[44]),
    .prog_clk_2_E_in(prog_clk_2_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[141]),
    .chany_top_in(cby_1__1__38_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__40_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__37_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_37_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_37_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_37_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_37_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_37_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_37_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_37_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_37_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__33_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_37_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_37_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_37_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_37_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_37_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_37_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_37_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_37_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__40_ccff_tail[0]),
    .chany_top_out(sb_1__1__33_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__33_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__33_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__33_ccff_tail[0])
  );


  sb_1__1_
  sb_5__7_
  (
    .clk_1_S_in(clk_2_wires[45]),
    .clk_1_W_out(clk_1_wires[79]),
    .clk_1_E_out(clk_1_wires[78]),
    .prog_clk_1_S_in(prog_clk_2_wires[45]),
    .prog_clk_1_W_out(prog_clk_1_wires[79]),
    .prog_clk_1_E_out(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[144]),
    .chany_top_in(cby_1__1__39_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__41_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__38_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_38_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_38_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_38_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_38_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_38_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_38_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_38_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_38_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__34_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_38_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_38_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_38_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_38_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_38_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_38_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_38_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_38_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__41_ccff_tail[0]),
    .chany_top_out(sb_1__1__34_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__34_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__34_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__34_ccff_tail[0])
  );


  sb_1__1_
  sb_6__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[152]),
    .chany_top_in(cby_1__1__41_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__42_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__40_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_40_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_40_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_40_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_40_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_40_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_40_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_40_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_40_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__35_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_40_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_40_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_40_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_40_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_40_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_40_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_40_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_40_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__42_ccff_tail[0]),
    .chany_top_out(sb_1__1__35_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__35_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__35_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__35_ccff_tail[0])
  );


  sb_1__1_
  sb_6__2_
  (
    .clk_2_N_in(clk_3_wires[25]),
    .clk_2_W_out(clk_2_wires[29]),
    .clk_2_E_out(clk_2_wires[27]),
    .prog_clk_2_N_in(prog_clk_3_wires[25]),
    .prog_clk_2_W_out(prog_clk_2_wires[29]),
    .prog_clk_2_E_out(prog_clk_2_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[155]),
    .chany_top_in(cby_1__1__42_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__43_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__41_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_41_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_41_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_41_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_41_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_41_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_41_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_41_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_41_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__36_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_41_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_41_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_41_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_41_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_41_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_41_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_41_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_41_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__43_ccff_tail[0]),
    .chany_top_out(sb_1__1__36_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__36_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__36_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__36_ccff_tail[0])
  );


  sb_1__1_
  sb_6__3_
  (
    .clk_3_S_out(clk_3_wires[24]),
    .clk_3_N_in(clk_3_wires[21]),
    .prog_clk_3_S_out(prog_clk_3_wires[24]),
    .prog_clk_3_N_in(prog_clk_3_wires[21]),
    .prog_clk_0_N_in(prog_clk_0_wires[158]),
    .chany_top_in(cby_1__1__43_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__44_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__42_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_42_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_42_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_42_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_42_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_42_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_42_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_42_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_42_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__37_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_42_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_42_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_42_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_42_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_42_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_42_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_42_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_42_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__44_ccff_tail[0]),
    .chany_top_out(sb_1__1__37_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__37_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__37_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__37_ccff_tail[0])
  );


  sb_1__1_
  sb_6__4_
  (
    .clk_3_S_out(clk_3_wires[20]),
    .clk_3_N_out(clk_3_wires[18]),
    .clk_3_W_in(clk_3_wires[7]),
    .prog_clk_3_S_out(prog_clk_3_wires[20]),
    .prog_clk_3_N_out(prog_clk_3_wires[18]),
    .prog_clk_3_W_in(prog_clk_3_wires[7]),
    .prog_clk_0_N_in(prog_clk_0_wires[161]),
    .chany_top_in(cby_1__1__44_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__45_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__43_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_43_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_43_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_43_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_43_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_43_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_43_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_43_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_43_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__38_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_43_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_43_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_43_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_43_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_43_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_43_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_43_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_43_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__45_ccff_tail[0]),
    .chany_top_out(sb_1__1__38_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__38_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__38_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__38_ccff_tail[0])
  );


  sb_1__1_
  sb_6__5_
  (
    .clk_3_N_out(clk_3_wires[22]),
    .clk_3_S_in(clk_3_wires[19]),
    .prog_clk_3_N_out(prog_clk_3_wires[22]),
    .prog_clk_3_S_in(prog_clk_3_wires[19]),
    .prog_clk_0_N_in(prog_clk_0_wires[164]),
    .chany_top_in(cby_1__1__45_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__46_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__44_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_44_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_44_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_44_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_44_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_44_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_44_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_44_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_44_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__39_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_44_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_44_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_44_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_44_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_44_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_44_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_44_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_44_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__46_ccff_tail[0]),
    .chany_top_out(sb_1__1__39_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__39_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__39_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__39_ccff_tail[0])
  );


  sb_1__1_
  sb_6__6_
  (
    .clk_2_S_in(clk_3_wires[23]),
    .clk_2_W_out(clk_2_wires[42]),
    .clk_2_E_out(clk_2_wires[40]),
    .prog_clk_2_S_in(prog_clk_3_wires[23]),
    .prog_clk_2_W_out(prog_clk_2_wires[42]),
    .prog_clk_2_E_out(prog_clk_2_wires[40]),
    .prog_clk_0_N_in(prog_clk_0_wires[167]),
    .chany_top_in(cby_1__1__46_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__47_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__45_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_45_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_45_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_45_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_45_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_45_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_45_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_45_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_45_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__40_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_45_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_45_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_45_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_45_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_45_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_45_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_45_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_45_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__47_ccff_tail[0]),
    .chany_top_out(sb_1__1__40_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__40_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__40_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__40_ccff_tail[0])
  );


  sb_1__1_
  sb_6__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[170]),
    .chany_top_in(cby_1__1__47_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__48_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__46_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_46_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_46_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_46_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_46_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_46_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_46_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_46_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_46_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__41_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_46_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_46_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_46_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_46_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_46_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_46_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_46_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_46_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__48_ccff_tail[0]),
    .chany_top_out(sb_1__1__41_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__41_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__41_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__41_ccff_tail[0])
  );


  sb_1__1_
  sb_7__1_
  (
    .clk_1_N_in(clk_2_wires[38]),
    .clk_1_W_out(clk_1_wires[86]),
    .clk_1_E_out(clk_1_wires[85]),
    .prog_clk_1_N_in(prog_clk_2_wires[38]),
    .prog_clk_1_W_out(prog_clk_1_wires[86]),
    .prog_clk_1_E_out(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[178]),
    .chany_top_in(cby_1__1__49_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__49_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__48_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_48_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_48_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_48_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_48_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_48_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_48_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_48_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_48_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__42_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_48_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_48_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_48_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_48_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_48_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_48_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_48_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_48_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__49_ccff_tail[0]),
    .chany_top_out(sb_1__1__42_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__42_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__42_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__42_ccff_tail[0])
  );


  sb_1__1_
  sb_7__2_
  (
    .clk_2_S_out(clk_2_wires[37]),
    .clk_2_N_out(clk_2_wires[35]),
    .clk_2_W_in(clk_2_wires[28]),
    .prog_clk_2_S_out(prog_clk_2_wires[37]),
    .prog_clk_2_N_out(prog_clk_2_wires[35]),
    .prog_clk_2_W_in(prog_clk_2_wires[28]),
    .prog_clk_0_N_in(prog_clk_0_wires[181]),
    .chany_top_in(cby_1__1__50_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__50_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__49_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_49_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_49_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_49_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_49_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_49_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_49_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_49_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_49_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__43_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_49_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_49_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_49_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_49_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_49_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_49_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_49_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_49_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__50_ccff_tail[0]),
    .chany_top_out(sb_1__1__43_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__43_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__43_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__43_ccff_tail[0])
  );


  sb_1__1_
  sb_7__3_
  (
    .clk_1_S_in(clk_2_wires[36]),
    .clk_1_W_out(clk_1_wires[93]),
    .clk_1_E_out(clk_1_wires[92]),
    .prog_clk_1_S_in(prog_clk_2_wires[36]),
    .prog_clk_1_W_out(prog_clk_1_wires[93]),
    .prog_clk_1_E_out(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[184]),
    .chany_top_in(cby_1__1__51_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__51_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__50_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_50_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_50_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_50_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_50_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_50_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_50_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_50_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_50_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__44_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_50_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_50_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_50_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_50_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_50_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_50_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_50_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_50_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__51_ccff_tail[0]),
    .chany_top_out(sb_1__1__44_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__44_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__44_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__44_ccff_tail[0])
  );


  sb_1__1_
  sb_7__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[187]),
    .chany_top_in(cby_1__1__52_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__52_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__51_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_51_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_51_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_51_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_51_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_51_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_51_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_51_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_51_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__45_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_51_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_51_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_51_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_51_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_51_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_51_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_51_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_51_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__52_ccff_tail[0]),
    .chany_top_out(sb_1__1__45_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__45_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__45_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__45_ccff_tail[0])
  );


  sb_1__1_
  sb_7__5_
  (
    .clk_1_N_in(clk_2_wires[51]),
    .clk_1_W_out(clk_1_wires[100]),
    .clk_1_E_out(clk_1_wires[99]),
    .prog_clk_1_N_in(prog_clk_2_wires[51]),
    .prog_clk_1_W_out(prog_clk_1_wires[100]),
    .prog_clk_1_E_out(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[190]),
    .chany_top_in(cby_1__1__53_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__53_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__52_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_52_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_52_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_52_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_52_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_52_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_52_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_52_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_52_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__46_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_52_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_52_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_52_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_52_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_52_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_52_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_52_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_52_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__53_ccff_tail[0]),
    .chany_top_out(sb_1__1__46_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__46_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__46_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__46_ccff_tail[0])
  );


  sb_1__1_
  sb_7__6_
  (
    .clk_2_S_out(clk_2_wires[50]),
    .clk_2_N_out(clk_2_wires[48]),
    .clk_2_W_in(clk_2_wires[41]),
    .prog_clk_2_S_out(prog_clk_2_wires[50]),
    .prog_clk_2_N_out(prog_clk_2_wires[48]),
    .prog_clk_2_W_in(prog_clk_2_wires[41]),
    .prog_clk_0_N_in(prog_clk_0_wires[193]),
    .chany_top_in(cby_1__1__54_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__54_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__53_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_53_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_53_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_53_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_53_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_53_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_53_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_53_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_53_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__47_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_53_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_53_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_53_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_53_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_53_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_53_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_53_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_53_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__54_ccff_tail[0]),
    .chany_top_out(sb_1__1__47_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__47_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__47_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__47_ccff_tail[0])
  );


  sb_1__1_
  sb_7__7_
  (
    .clk_1_S_in(clk_2_wires[49]),
    .clk_1_W_out(clk_1_wires[107]),
    .clk_1_E_out(clk_1_wires[106]),
    .prog_clk_1_S_in(prog_clk_2_wires[49]),
    .prog_clk_1_W_out(prog_clk_1_wires[107]),
    .prog_clk_1_E_out(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[196]),
    .chany_top_in(cby_1__1__55_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_lower[0]),
    .chanx_right_in(cbx_1__1__55_chanx_left_out[0:19]),
    .right_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__54_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_54_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_54_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_54_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_54_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_54_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_54_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_54_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_54_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__48_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_54_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_54_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_54_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_54_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_54_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_54_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_54_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_54_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(cbx_1__1__55_ccff_tail[0]),
    .chany_top_out(sb_1__1__48_chany_top_out[0:19]),
    .chanx_right_out(sb_1__1__48_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__1__48_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_tail(sb_1__1__48_ccff_tail[0])
  );


  sb_1__2_
  sb_1__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[40]),
    .chanx_right_in(cbx_1__8__1_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_7_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_7_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_7_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_7_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_7_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_7_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_7_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_7_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__0_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_7_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_7_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_7_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_7_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_7_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_7_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_7_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_7_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_1_ccff_tail[0]),
    .chanx_right_out(sb_1__8__0_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__0_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__0_ccff_tail[0])
  );


  sb_1__2_
  sb_2__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[68]),
    .SC_OUT_BOT(scff_Wires[37]),
    .SC_IN_BOT(scff_Wires[36]),
    .chanx_right_in(cbx_1__8__2_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__15_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_15_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_15_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_15_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_15_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_15_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_15_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_15_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_15_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__1_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_15_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_15_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_15_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_15_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_15_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_15_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_15_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_15_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_2_ccff_tail[0]),
    .chanx_right_out(sb_1__8__1_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__1_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__1_ccff_tail[0])
  );


  sb_1__2_
  sb_3__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[94]),
    .chanx_right_in(cbx_1__8__3_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__23_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_23_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_23_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_23_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_23_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_23_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_23_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_23_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_23_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__2_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_23_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_23_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_23_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_23_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_23_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_23_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_23_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_23_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_3_ccff_tail[0]),
    .chanx_right_out(sb_1__8__2_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__2_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__2_ccff_tail[0])
  );


  sb_1__2_
  sb_4__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[120]),
    .SC_OUT_BOT(scff_Wires[74]),
    .SC_IN_BOT(scff_Wires[73]),
    .chanx_right_in(cbx_1__8__4_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__31_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_31_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_31_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_31_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_31_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_31_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_31_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_31_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_31_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__3_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_31_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_31_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_31_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_31_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_31_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_31_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_31_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_31_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_4_ccff_tail[0]),
    .chanx_right_out(sb_1__8__3_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__3_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__3_ccff_tail[0])
  );


  sb_1__2_
  sb_5__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[146]),
    .chanx_right_in(cbx_1__8__5_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__39_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_39_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_39_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_39_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_39_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_39_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_39_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_39_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_39_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__4_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_39_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_39_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_39_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_39_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_39_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_39_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_39_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_39_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_5_ccff_tail[0]),
    .chanx_right_out(sb_1__8__4_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__4_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__4_ccff_tail[0])
  );


  sb_1__2_
  sb_6__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[172]),
    .SC_OUT_BOT(scff_Wires[111]),
    .SC_IN_BOT(scff_Wires[110]),
    .chanx_right_in(cbx_1__8__6_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__47_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_47_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_47_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_47_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_47_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_47_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_47_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_47_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_47_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__5_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_47_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_47_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_47_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_47_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_47_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_47_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_47_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_47_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_6_ccff_tail[0]),
    .chanx_right_out(sb_1__8__5_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__5_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__5_ccff_tail[0])
  );


  sb_1__2_
  sb_7__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[198]),
    .chanx_right_in(cbx_1__8__7_chanx_left_out[0:19]),
    .right_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
    .right_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_upper[0]),
    .right_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_upper[0]),
    .right_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_upper[0]),
    .right_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_upper[0]),
    .right_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_upper[0]),
    .right_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_upper[0]),
    .right_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_upper[0]),
    .right_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_upper[0]),
    .chany_bottom_in(cby_1__1__55_chany_top_out[0:19]),
    .bottom_left_grid_pin_42_(grid_clb_55_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_55_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_55_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_55_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_55_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_55_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_55_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_55_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__6_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_55_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_55_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_55_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_55_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_55_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_55_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_55_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_55_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_top_7_ccff_tail[0]),
    .chanx_right_out(sb_1__8__6_chanx_right_out[0:19]),
    .chany_bottom_out(sb_1__8__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_1__8__6_chanx_left_out[0:19]),
    .ccff_tail(sb_1__8__6_ccff_tail[0])
  );


  sb_2__0_
  sb_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[201]),
    .chany_top_in(cby_8__1__0_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
    .chanx_left_in(cbx_1__0__7_chanx_right_out[0:19]),
    .left_bottom_grid_pin_1_(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_3_(grid_io_bottom_0_top_width_0_height_0__pin_3_lower[0]),
    .left_bottom_grid_pin_5_(grid_io_bottom_0_top_width_0_height_0__pin_5_lower[0]),
    .left_bottom_grid_pin_7_(grid_io_bottom_0_top_width_0_height_0__pin_7_lower[0]),
    .left_bottom_grid_pin_9_(grid_io_bottom_0_top_width_0_height_0__pin_9_lower[0]),
    .left_bottom_grid_pin_11_(grid_io_bottom_0_top_width_0_height_0__pin_11_lower[0]),
    .left_bottom_grid_pin_13_(grid_io_bottom_0_top_width_0_height_0__pin_13_lower[0]),
    .left_bottom_grid_pin_15_(grid_io_bottom_0_top_width_0_height_0__pin_15_lower[0]),
    .left_bottom_grid_pin_17_(grid_io_bottom_0_top_width_0_height_0__pin_17_lower[0]),
    .ccff_head(grid_io_right_7_ccff_tail[0]),
    .chany_top_out(sb_8__0__0_chany_top_out[0:19]),
    .chanx_left_out(sb_8__0__0_chanx_left_out[0:19]),
    .ccff_tail(sb_8__0__0_ccff_tail[0])
  );


  sb_2__1_
  sb_8__1_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[204]),
    .chany_top_in(cby_8__1__1_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__0_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_56_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_56_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_56_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_56_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_56_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_56_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_56_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_56_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__49_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_56_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_56_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_56_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_56_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_56_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_56_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_56_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_56_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_6_ccff_tail[0]),
    .chany_top_out(sb_8__1__0_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__0_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__0_ccff_tail[0])
  );


  sb_2__1_
  sb_8__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[207]),
    .chany_top_in(cby_8__1__2_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__1_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_57_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_57_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_57_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_57_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_57_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_57_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_57_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_57_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__50_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_57_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_57_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_57_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_57_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_57_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_57_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_57_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_57_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_5_ccff_tail[0]),
    .chany_top_out(sb_8__1__1_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__1_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__1_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__1_ccff_tail[0])
  );


  sb_2__1_
  sb_8__3_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[210]),
    .chany_top_in(cby_8__1__3_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__2_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_58_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_58_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_58_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_58_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_58_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_58_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_58_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_58_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__51_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_58_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_58_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_58_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_58_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_58_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_58_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_58_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_58_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_4_ccff_tail[0]),
    .chany_top_out(sb_8__1__2_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__2_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__2_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__2_ccff_tail[0])
  );


  sb_2__1_
  sb_8__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[213]),
    .chany_top_in(cby_8__1__4_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__3_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_59_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_59_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_59_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_59_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_59_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_59_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_59_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_59_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__52_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_59_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_59_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_59_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_59_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_59_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_59_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_59_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_59_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_3_ccff_tail[0]),
    .chany_top_out(sb_8__1__3_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__3_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__3_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__3_ccff_tail[0])
  );


  sb_2__1_
  sb_8__5_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[216]),
    .chany_top_in(cby_8__1__5_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__4_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_60_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_60_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_60_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_60_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_60_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_60_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_60_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_60_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__53_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_60_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_60_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_60_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_60_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_60_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_60_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_60_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_60_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_2_ccff_tail[0]),
    .chany_top_out(sb_8__1__4_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__4_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__4_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__4_ccff_tail[0])
  );


  sb_2__1_
  sb_8__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[219]),
    .chany_top_in(cby_8__1__6_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__5_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_61_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_61_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_61_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_61_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_61_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_61_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_61_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_61_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__54_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_61_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_61_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_61_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_61_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_61_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_61_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_61_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_61_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_1_ccff_tail[0]),
    .chany_top_out(sb_8__1__5_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__5_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__5_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__5_ccff_tail[0])
  );


  sb_2__1_
  sb_8__7_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[222]),
    .chany_top_in(cby_8__1__7_chany_bottom_out[0:19]),
    .top_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_lower[0]),
    .top_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_lower[0]),
    .top_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_lower[0]),
    .top_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_lower[0]),
    .top_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_lower[0]),
    .top_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_lower[0]),
    .top_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_lower[0]),
    .top_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_lower[0]),
    .top_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
    .chany_bottom_in(cby_8__1__6_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_62_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_62_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_62_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_62_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_62_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_62_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_62_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_62_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__1__55_chanx_right_out[0:19]),
    .left_bottom_grid_pin_34_(grid_clb_62_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_62_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_62_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_62_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_62_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_62_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_62_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_62_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(grid_io_right_0_ccff_tail[0]),
    .chany_top_out(sb_8__1__6_chany_top_out[0:19]),
    .chany_bottom_out(sb_8__1__6_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__1__6_chanx_left_out[0:19]),
    .ccff_tail(sb_8__1__6_ccff_tail[0])
  );


  sb_2__2_
  sb_8__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[224]),
    .SC_OUT_BOT(sc_tail),
    .SC_IN_BOT(scff_Wires[147]),
    .chany_bottom_in(cby_8__1__7_chany_top_out[0:19]),
    .bottom_right_grid_pin_1_(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
    .bottom_left_grid_pin_42_(grid_clb_63_right_width_0_height_0__pin_42_upper[0]),
    .bottom_left_grid_pin_43_(grid_clb_63_right_width_0_height_0__pin_43_upper[0]),
    .bottom_left_grid_pin_44_(grid_clb_63_right_width_0_height_0__pin_44_upper[0]),
    .bottom_left_grid_pin_45_(grid_clb_63_right_width_0_height_0__pin_45_upper[0]),
    .bottom_left_grid_pin_46_(grid_clb_63_right_width_0_height_0__pin_46_upper[0]),
    .bottom_left_grid_pin_47_(grid_clb_63_right_width_0_height_0__pin_47_upper[0]),
    .bottom_left_grid_pin_48_(grid_clb_63_right_width_0_height_0__pin_48_upper[0]),
    .bottom_left_grid_pin_49_(grid_clb_63_right_width_0_height_0__pin_49_upper[0]),
    .chanx_left_in(cbx_1__8__7_chanx_right_out[0:19]),
    .left_top_grid_pin_1_(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
    .left_bottom_grid_pin_34_(grid_clb_63_top_width_0_height_0__pin_34_lower[0]),
    .left_bottom_grid_pin_35_(grid_clb_63_top_width_0_height_0__pin_35_lower[0]),
    .left_bottom_grid_pin_36_(grid_clb_63_top_width_0_height_0__pin_36_lower[0]),
    .left_bottom_grid_pin_37_(grid_clb_63_top_width_0_height_0__pin_37_lower[0]),
    .left_bottom_grid_pin_38_(grid_clb_63_top_width_0_height_0__pin_38_lower[0]),
    .left_bottom_grid_pin_39_(grid_clb_63_top_width_0_height_0__pin_39_lower[0]),
    .left_bottom_grid_pin_40_(grid_clb_63_top_width_0_height_0__pin_40_lower[0]),
    .left_bottom_grid_pin_41_(grid_clb_63_top_width_0_height_0__pin_41_lower[0]),
    .ccff_head(ccff_head[0]),
    .chany_bottom_out(sb_8__8__0_chany_bottom_out[0:19]),
    .chanx_left_out(sb_8__8__0_chanx_left_out[0:19]),
    .ccff_tail(sb_8__8__0_ccff_tail[0])
  );


  cbx_1__0_
  cbx_1__0_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[5]),
    .prog_clk_0_N_in(prog_clk_0_wires[0]),
    .SC_OUT_BOT(scff_Wires[18]),
    .SC_IN_TOP(scff_Wires[17]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_7_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_7_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_7_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_7_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_7_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_7_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_7_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_7_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_7_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_7_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_7_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_7_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_7_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_7_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_7_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_7_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_7_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_7_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79:87]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79:87]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79:87]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__0_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_7_ccff_tail[0])
  );


  cbx_1__0_
  cbx_2__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[43]),
    .SC_OUT_TOP(scff_Wires[20]),
    .SC_IN_BOT(scff_Wires[19]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_6_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_6_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_6_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_6_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_6_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_6_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_6_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_6_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_6_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_6_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_6_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_6_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_6_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_6_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_6_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_6_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_6_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_6_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70:78]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70:78]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70:78]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__1_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_6_ccff_tail[0])
  );


  cbx_1__0_
  cbx_3__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[69]),
    .SC_OUT_BOT(scff_Wires[55]),
    .SC_IN_TOP(scff_Wires[54]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_5_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_5_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_5_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_5_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_5_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_5_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_5_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_5_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_5_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_5_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_5_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_5_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_5_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_5_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_5_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_5_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_5_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_5_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61:69]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61:69]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61:69]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__2_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_5_ccff_tail[0])
  );


  cbx_1__0_
  cbx_4__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[95]),
    .SC_OUT_TOP(scff_Wires[57]),
    .SC_IN_BOT(scff_Wires[56]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_4_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_4_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_4_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_4_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_4_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_4_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_4_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_4_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_4_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_4_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_4_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_4_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_4_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_4_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_4_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_4_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_4_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_4_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52:60]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52:60]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52:60]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__3_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_4_ccff_tail[0])
  );


  cbx_1__0_
  cbx_5__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[121]),
    .SC_OUT_BOT(scff_Wires[92]),
    .SC_IN_TOP(scff_Wires[91]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_3_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_3_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_3_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_3_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_3_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_3_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_3_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_3_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_3_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_3_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_3_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_3_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_3_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_3_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_3_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_3_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_3_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_3_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43:51]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43:51]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43:51]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__4_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__4_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_3_ccff_tail[0])
  );


  cbx_1__0_
  cbx_6__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[147]),
    .SC_OUT_TOP(scff_Wires[94]),
    .SC_IN_BOT(scff_Wires[93]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_2_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_2_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_2_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_2_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_2_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_2_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_2_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_2_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_2_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_2_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_2_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_2_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_2_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_2_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_2_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_2_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_2_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_2_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34:42]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34:42]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34:42]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__5_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__5_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_2_ccff_tail[0])
  );


  cbx_1__0_
  cbx_7__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[173]),
    .SC_OUT_BOT(scff_Wires[129]),
    .SC_IN_TOP(scff_Wires[128]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_1_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_1_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_1_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_1_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_1_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_1_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_1_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_1_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_1_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_1_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_1_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_1_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_1_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_1_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_1_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_1_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_1_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_1_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25:33]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25:33]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25:33]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__0__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__0__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__6_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__6_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_1_ccff_tail[0])
  );


  cbx_1__0_
  cbx_8__0_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[199]),
    .SC_OUT_TOP(scff_Wires[131]),
    .SC_IN_BOT(scff_Wires[130]),
    .top_width_0_height_0__pin_17_lower(grid_io_bottom_0_top_width_0_height_0__pin_17_lower[0]),
    .top_width_0_height_0__pin_17_upper(grid_io_bottom_0_top_width_0_height_0__pin_17_upper[0]),
    .top_width_0_height_0__pin_15_lower(grid_io_bottom_0_top_width_0_height_0__pin_15_lower[0]),
    .top_width_0_height_0__pin_15_upper(grid_io_bottom_0_top_width_0_height_0__pin_15_upper[0]),
    .top_width_0_height_0__pin_13_lower(grid_io_bottom_0_top_width_0_height_0__pin_13_lower[0]),
    .top_width_0_height_0__pin_13_upper(grid_io_bottom_0_top_width_0_height_0__pin_13_upper[0]),
    .top_width_0_height_0__pin_11_lower(grid_io_bottom_0_top_width_0_height_0__pin_11_lower[0]),
    .top_width_0_height_0__pin_11_upper(grid_io_bottom_0_top_width_0_height_0__pin_11_upper[0]),
    .top_width_0_height_0__pin_9_lower(grid_io_bottom_0_top_width_0_height_0__pin_9_lower[0]),
    .top_width_0_height_0__pin_9_upper(grid_io_bottom_0_top_width_0_height_0__pin_9_upper[0]),
    .top_width_0_height_0__pin_7_lower(grid_io_bottom_0_top_width_0_height_0__pin_7_lower[0]),
    .top_width_0_height_0__pin_7_upper(grid_io_bottom_0_top_width_0_height_0__pin_7_upper[0]),
    .top_width_0_height_0__pin_5_lower(grid_io_bottom_0_top_width_0_height_0__pin_5_lower[0]),
    .top_width_0_height_0__pin_5_upper(grid_io_bottom_0_top_width_0_height_0__pin_5_upper[0]),
    .top_width_0_height_0__pin_3_lower(grid_io_bottom_0_top_width_0_height_0__pin_3_lower[0]),
    .top_width_0_height_0__pin_3_upper(grid_io_bottom_0_top_width_0_height_0__pin_3_upper[0]),
    .top_width_0_height_0__pin_1_lower(grid_io_bottom_0_top_width_0_height_0__pin_1_lower[0]),
    .top_width_0_height_0__pin_1_upper(grid_io_bottom_0_top_width_0_height_0__pin_1_upper[0]),
    .top_width_0_height_0__pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
    .top_width_0_height_0__pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
    .top_width_0_height_0__pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
    .top_width_0_height_0__pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
    .top_width_0_height_0__pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
    .top_width_0_height_0__pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
    .top_width_0_height_0__pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
    .top_width_0_height_0__pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
    .top_width_0_height_0__pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16:24]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16:24]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16:24]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__0__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__0__0_chanx_left_out[0:19]),
    .ccff_head(sb_8__0__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__0__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__0__7_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__0__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_2_(cbx_1__0__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_4_(cbx_1__0__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_6_(cbx_1__0__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_8_(cbx_1__0__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_10_(cbx_1__0__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_12_(cbx_1__0__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_14_(cbx_1__0__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_16_(cbx_1__0__7_bottom_grid_pin_16_[0]),
    .ccff_tail(grid_io_bottom_0_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__1_
  (
    .clk_1_S_out(clk_1_wires[4]),
    .clk_1_N_out(clk_1_wires[3]),
    .clk_1_E_in(clk_1_wires[2]),
    .prog_clk_1_S_out(prog_clk_1_wires[4]),
    .prog_clk_1_N_out(prog_clk_1_wires[3]),
    .prog_clk_1_E_in(prog_clk_1_wires[2]),
    .prog_clk_0_N_in(prog_clk_0_wires[6]),
    .prog_clk_0_W_out(prog_clk_0_wires[4]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[0]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[0]),
    .SC_OUT_BOT(scff_Wires[15]),
    .SC_IN_TOP(scff_Wires[14]),
    .chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__0_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__0_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__0_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__0_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__0_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__0_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__0_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__0_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__0_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[11]),
    .prog_clk_0_W_out(prog_clk_0_wires[10]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[1]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[1]),
    .SC_OUT_BOT(scff_Wires[13]),
    .SC_IN_TOP(scff_Wires[12]),
    .chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__1_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__1_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__1_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__1_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__1_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__1_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__1_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__1_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__1_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__3_
  (
    .clk_1_S_out(clk_1_wires[11]),
    .clk_1_N_out(clk_1_wires[10]),
    .clk_1_E_in(clk_1_wires[9]),
    .prog_clk_1_S_out(prog_clk_1_wires[11]),
    .prog_clk_1_N_out(prog_clk_1_wires[10]),
    .prog_clk_1_E_in(prog_clk_1_wires[9]),
    .prog_clk_0_N_in(prog_clk_0_wires[16]),
    .prog_clk_0_W_out(prog_clk_0_wires[15]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[2]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[2]),
    .SC_OUT_BOT(scff_Wires[11]),
    .SC_IN_TOP(scff_Wires[10]),
    .chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__2_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__2_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__2_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__2_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__2_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__2_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__2_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__2_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__2_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[21]),
    .prog_clk_0_W_out(prog_clk_0_wires[20]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[3]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[3]),
    .SC_OUT_BOT(scff_Wires[9]),
    .SC_IN_TOP(scff_Wires[8]),
    .chanx_left_in(sb_0__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__3_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__3_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__3_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__3_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__3_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__3_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__3_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__3_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__3_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__5_
  (
    .clk_1_S_out(clk_1_wires[18]),
    .clk_1_N_out(clk_1_wires[17]),
    .clk_1_E_in(clk_1_wires[16]),
    .prog_clk_1_S_out(prog_clk_1_wires[18]),
    .prog_clk_1_N_out(prog_clk_1_wires[17]),
    .prog_clk_1_E_in(prog_clk_1_wires[16]),
    .prog_clk_0_N_in(prog_clk_0_wires[26]),
    .prog_clk_0_W_out(prog_clk_0_wires[25]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[4]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[4]),
    .SC_OUT_BOT(scff_Wires[7]),
    .SC_IN_TOP(scff_Wires[6]),
    .chanx_left_in(sb_0__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__4_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__4_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__4_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__4_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__4_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__4_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__4_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__4_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__4_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[31]),
    .prog_clk_0_W_out(prog_clk_0_wires[30]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[5]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[5]),
    .SC_OUT_BOT(scff_Wires[5]),
    .SC_IN_TOP(scff_Wires[4]),
    .chanx_left_in(sb_0__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__5_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__5_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__5_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__5_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__5_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__5_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__5_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__5_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__5_ccff_tail[0])
  );


  cbx_1__1_
  cbx_1__7_
  (
    .clk_1_S_out(clk_1_wires[25]),
    .clk_1_N_out(clk_1_wires[24]),
    .clk_1_E_in(clk_1_wires[23]),
    .prog_clk_1_S_out(prog_clk_1_wires[25]),
    .prog_clk_1_N_out(prog_clk_1_wires[24]),
    .prog_clk_1_E_in(prog_clk_1_wires[23]),
    .prog_clk_0_N_in(prog_clk_0_wires[36]),
    .prog_clk_0_W_out(prog_clk_0_wires[35]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[6]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[6]),
    .SC_OUT_BOT(scff_Wires[3]),
    .SC_IN_TOP(scff_Wires[2]),
    .chanx_left_in(sb_0__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__6_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__6_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__6_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__6_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__6_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__6_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__6_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__6_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__6_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__1_
  (
    .clk_1_S_out(clk_1_wires[6]),
    .clk_1_N_out(clk_1_wires[5]),
    .clk_1_W_in(clk_1_wires[1]),
    .prog_clk_1_S_out(prog_clk_1_wires[6]),
    .prog_clk_1_N_out(prog_clk_1_wires[5]),
    .prog_clk_1_W_in(prog_clk_1_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[46]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[7]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[7]),
    .SC_OUT_TOP(scff_Wires[22]),
    .SC_IN_BOT(scff_Wires[21]),
    .chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__7_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__7_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__7_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__7_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__7_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__7_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__7_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__7_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__7_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__7_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__2_
  (
    .clk_2_W_out(clk_2_wires[4]),
    .clk_2_E_in(clk_2_wires[3]),
    .prog_clk_2_W_out(prog_clk_2_wires[4]),
    .prog_clk_2_E_in(prog_clk_2_wires[3]),
    .prog_clk_0_N_in(prog_clk_0_wires[49]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[8]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[8]),
    .SC_OUT_TOP(scff_Wires[24]),
    .SC_IN_BOT(scff_Wires[23]),
    .chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__8_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__8_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__8_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__8_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__8_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__8_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__8_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__8_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__8_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__8_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__8_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__8_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__8_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__8_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__8_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__8_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__8_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__8_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__3_
  (
    .clk_1_S_out(clk_1_wires[13]),
    .clk_1_N_out(clk_1_wires[12]),
    .clk_1_W_in(clk_1_wires[8]),
    .prog_clk_1_S_out(prog_clk_1_wires[13]),
    .prog_clk_1_N_out(prog_clk_1_wires[12]),
    .prog_clk_1_W_in(prog_clk_1_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[52]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[9]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[9]),
    .SC_OUT_TOP(scff_Wires[26]),
    .SC_IN_BOT(scff_Wires[25]),
    .chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__9_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__9_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__9_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__9_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__9_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__9_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__9_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__9_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__9_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__9_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__9_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__9_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__9_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__9_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__9_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__9_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__9_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__9_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__9_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[55]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[10]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[10]),
    .SC_OUT_TOP(scff_Wires[28]),
    .SC_IN_BOT(scff_Wires[27]),
    .chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__10_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__10_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__10_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__10_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__10_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__10_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__10_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__10_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__10_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__10_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__10_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__10_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__10_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__10_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__10_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__10_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__10_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__10_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__10_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__5_
  (
    .clk_1_S_out(clk_1_wires[20]),
    .clk_1_N_out(clk_1_wires[19]),
    .clk_1_W_in(clk_1_wires[15]),
    .prog_clk_1_S_out(prog_clk_1_wires[20]),
    .prog_clk_1_N_out(prog_clk_1_wires[19]),
    .prog_clk_1_W_in(prog_clk_1_wires[15]),
    .prog_clk_0_N_in(prog_clk_0_wires[58]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[11]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[11]),
    .SC_OUT_TOP(scff_Wires[30]),
    .SC_IN_BOT(scff_Wires[29]),
    .chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__11_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__11_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__11_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__11_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__11_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__11_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__11_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__11_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__11_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__11_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__11_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__11_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__11_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__11_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__11_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__11_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__11_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__11_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__11_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__6_
  (
    .clk_2_W_out(clk_2_wires[17]),
    .clk_2_E_in(clk_2_wires[16]),
    .prog_clk_2_W_out(prog_clk_2_wires[17]),
    .prog_clk_2_E_in(prog_clk_2_wires[16]),
    .prog_clk_0_N_in(prog_clk_0_wires[61]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[12]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[12]),
    .SC_OUT_TOP(scff_Wires[32]),
    .SC_IN_BOT(scff_Wires[31]),
    .chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__12_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__12_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__12_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__12_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__12_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__12_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__12_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__12_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__12_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__12_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__12_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__12_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__12_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__12_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__12_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__12_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__12_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__12_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__12_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__12_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__12_ccff_tail[0])
  );


  cbx_1__1_
  cbx_2__7_
  (
    .clk_1_S_out(clk_1_wires[27]),
    .clk_1_N_out(clk_1_wires[26]),
    .clk_1_W_in(clk_1_wires[22]),
    .prog_clk_1_S_out(prog_clk_1_wires[27]),
    .prog_clk_1_N_out(prog_clk_1_wires[26]),
    .prog_clk_1_W_in(prog_clk_1_wires[22]),
    .prog_clk_0_N_in(prog_clk_0_wires[64]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[13]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[13]),
    .SC_OUT_TOP(scff_Wires[34]),
    .SC_IN_BOT(scff_Wires[33]),
    .chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__13_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__13_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__13_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__13_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__13_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__13_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__13_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__13_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__13_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__13_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__13_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__13_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__13_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__13_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__13_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__13_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__13_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__13_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__13_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__13_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__13_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__1_
  (
    .clk_1_S_out(clk_1_wires[32]),
    .clk_1_N_out(clk_1_wires[31]),
    .clk_1_E_in(clk_1_wires[30]),
    .prog_clk_1_S_out(prog_clk_1_wires[32]),
    .prog_clk_1_N_out(prog_clk_1_wires[31]),
    .prog_clk_1_E_in(prog_clk_1_wires[30]),
    .prog_clk_0_N_in(prog_clk_0_wires[72]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[14]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[14]),
    .SC_OUT_BOT(scff_Wires[52]),
    .SC_IN_TOP(scff_Wires[51]),
    .chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__14_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__14_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__14_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__14_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__14_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__14_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__14_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__14_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__14_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__14_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__14_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__14_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__14_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__14_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__14_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__14_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__14_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__14_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__14_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__14_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__14_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__2_
  (
    .clk_2_E_out(clk_2_wires[2]),
    .clk_2_W_in(clk_2_wires[1]),
    .prog_clk_2_E_out(prog_clk_2_wires[2]),
    .prog_clk_2_W_in(prog_clk_2_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[75]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[15]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[15]),
    .SC_OUT_BOT(scff_Wires[50]),
    .SC_IN_TOP(scff_Wires[49]),
    .chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__15_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__15_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__15_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__15_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__15_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__15_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__15_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__15_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__15_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__15_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__15_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__15_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__15_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__15_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__15_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__15_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__15_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__15_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__15_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__15_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__15_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__3_
  (
    .clk_1_S_out(clk_1_wires[39]),
    .clk_1_N_out(clk_1_wires[38]),
    .clk_1_E_in(clk_1_wires[37]),
    .prog_clk_1_S_out(prog_clk_1_wires[39]),
    .prog_clk_1_N_out(prog_clk_1_wires[38]),
    .prog_clk_1_E_in(prog_clk_1_wires[37]),
    .prog_clk_0_N_in(prog_clk_0_wires[78]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[16]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[16]),
    .SC_OUT_BOT(scff_Wires[48]),
    .SC_IN_TOP(scff_Wires[47]),
    .chanx_left_in(sb_1__1__9_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__16_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__16_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__16_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__16_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__16_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__16_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__16_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__16_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__16_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__16_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__16_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__16_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__16_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__16_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__16_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__16_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__16_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__16_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__16_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__16_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__16_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__4_
  (
    .clk_3_W_out(clk_3_wires[9]),
    .clk_3_E_in(clk_3_wires[8]),
    .prog_clk_3_W_out(prog_clk_3_wires[9]),
    .prog_clk_3_E_in(prog_clk_3_wires[8]),
    .prog_clk_0_N_in(prog_clk_0_wires[81]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[17]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[17]),
    .SC_OUT_BOT(scff_Wires[46]),
    .SC_IN_TOP(scff_Wires[45]),
    .chanx_left_in(sb_1__1__10_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__17_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__17_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__17_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__17_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__17_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__17_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__17_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__17_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__17_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__17_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__17_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__17_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__17_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__17_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__17_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__17_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__17_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__17_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__17_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__17_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__17_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__5_
  (
    .clk_1_S_out(clk_1_wires[46]),
    .clk_1_N_out(clk_1_wires[45]),
    .clk_1_E_in(clk_1_wires[44]),
    .prog_clk_1_S_out(prog_clk_1_wires[46]),
    .prog_clk_1_N_out(prog_clk_1_wires[45]),
    .prog_clk_1_E_in(prog_clk_1_wires[44]),
    .prog_clk_0_N_in(prog_clk_0_wires[84]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[18]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[18]),
    .SC_OUT_BOT(scff_Wires[44]),
    .SC_IN_TOP(scff_Wires[43]),
    .chanx_left_in(sb_1__1__11_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__18_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__18_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__18_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__18_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__18_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__18_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__18_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__18_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__18_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__18_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__18_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__18_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__18_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__18_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__18_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__18_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__18_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__18_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__18_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__18_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__18_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__6_
  (
    .clk_2_E_out(clk_2_wires[15]),
    .clk_2_W_in(clk_2_wires[14]),
    .prog_clk_2_E_out(prog_clk_2_wires[15]),
    .prog_clk_2_W_in(prog_clk_2_wires[14]),
    .prog_clk_0_N_in(prog_clk_0_wires[87]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[19]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[19]),
    .SC_OUT_BOT(scff_Wires[42]),
    .SC_IN_TOP(scff_Wires[41]),
    .chanx_left_in(sb_1__1__12_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__19_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__19_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__19_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__19_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__19_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__19_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__19_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__19_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__19_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__19_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__19_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__19_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__19_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__19_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__19_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__19_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__19_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__19_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__19_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__19_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__19_ccff_tail[0])
  );


  cbx_1__1_
  cbx_3__7_
  (
    .clk_1_S_out(clk_1_wires[53]),
    .clk_1_N_out(clk_1_wires[52]),
    .clk_1_E_in(clk_1_wires[51]),
    .prog_clk_1_S_out(prog_clk_1_wires[53]),
    .prog_clk_1_N_out(prog_clk_1_wires[52]),
    .prog_clk_1_E_in(prog_clk_1_wires[51]),
    .prog_clk_0_N_in(prog_clk_0_wires[90]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[20]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[20]),
    .SC_OUT_BOT(scff_Wires[40]),
    .SC_IN_TOP(scff_Wires[39]),
    .chanx_left_in(sb_1__1__13_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__20_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__20_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__20_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__20_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__20_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__20_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__20_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__20_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__20_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__20_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__20_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__20_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__20_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__20_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__20_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__20_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__20_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__20_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__20_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__20_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__20_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__1_
  (
    .clk_1_S_out(clk_1_wires[34]),
    .clk_1_N_out(clk_1_wires[33]),
    .clk_1_W_in(clk_1_wires[29]),
    .prog_clk_1_S_out(prog_clk_1_wires[34]),
    .prog_clk_1_N_out(prog_clk_1_wires[33]),
    .prog_clk_1_W_in(prog_clk_1_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[98]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[21]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[21]),
    .SC_OUT_TOP(scff_Wires[59]),
    .SC_IN_BOT(scff_Wires[58]),
    .chanx_left_in(sb_1__1__14_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__21_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__21_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__21_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__21_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__21_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__21_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__21_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__21_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__21_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__21_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__21_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__21_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__21_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__21_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__21_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__21_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__21_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__21_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__21_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__21_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__21_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[101]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[22]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[22]),
    .SC_OUT_TOP(scff_Wires[61]),
    .SC_IN_BOT(scff_Wires[60]),
    .chanx_left_in(sb_1__1__15_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__22_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__22_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__22_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__22_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__22_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__22_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__22_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__22_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__22_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__22_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__22_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__22_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__22_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__22_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__22_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__22_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__22_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__22_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__22_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__22_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__22_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__3_
  (
    .clk_1_S_out(clk_1_wires[41]),
    .clk_1_N_out(clk_1_wires[40]),
    .clk_1_W_in(clk_1_wires[36]),
    .prog_clk_1_S_out(prog_clk_1_wires[41]),
    .prog_clk_1_N_out(prog_clk_1_wires[40]),
    .prog_clk_1_W_in(prog_clk_1_wires[36]),
    .prog_clk_0_N_in(prog_clk_0_wires[104]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[23]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[23]),
    .SC_OUT_TOP(scff_Wires[63]),
    .SC_IN_BOT(scff_Wires[62]),
    .chanx_left_in(sb_1__1__16_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__23_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__23_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__23_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__23_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__23_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__23_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__23_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__23_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__23_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__23_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__23_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__23_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__23_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__23_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__23_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__23_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__23_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__23_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__23_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__23_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__23_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__4_
  (
    .clk_3_W_out(clk_3_wires[4]),
    .clk_3_E_in(clk_3_wires[3]),
    .prog_clk_3_W_out(prog_clk_3_wires[4]),
    .prog_clk_3_E_in(prog_clk_3_wires[3]),
    .prog_clk_0_N_in(prog_clk_0_wires[107]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[24]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[24]),
    .SC_OUT_TOP(scff_Wires[65]),
    .SC_IN_BOT(scff_Wires[64]),
    .chanx_left_in(sb_1__1__17_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__24_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__24_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__24_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__24_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__24_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__24_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__24_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__24_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__24_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__24_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__24_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__24_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__24_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__24_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__24_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__24_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__24_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__24_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__24_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__24_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__24_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__5_
  (
    .clk_1_S_out(clk_1_wires[48]),
    .clk_1_N_out(clk_1_wires[47]),
    .clk_1_W_in(clk_1_wires[43]),
    .prog_clk_1_S_out(prog_clk_1_wires[48]),
    .prog_clk_1_N_out(prog_clk_1_wires[47]),
    .prog_clk_1_W_in(prog_clk_1_wires[43]),
    .prog_clk_0_N_in(prog_clk_0_wires[110]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[25]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[25]),
    .SC_OUT_TOP(scff_Wires[67]),
    .SC_IN_BOT(scff_Wires[66]),
    .chanx_left_in(sb_1__1__18_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__25_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__25_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__25_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__25_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__25_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__25_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__25_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__25_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__25_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__25_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__25_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__25_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__25_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__25_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__25_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__25_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__25_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__25_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__25_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__25_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__25_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[113]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[26]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[26]),
    .SC_OUT_TOP(scff_Wires[69]),
    .SC_IN_BOT(scff_Wires[68]),
    .chanx_left_in(sb_1__1__19_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__26_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__26_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__26_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__26_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__26_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__26_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__26_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__26_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__26_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__26_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__26_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__26_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__26_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__26_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__26_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__26_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__26_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__26_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__26_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__26_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__26_ccff_tail[0])
  );


  cbx_1__1_
  cbx_4__7_
  (
    .clk_1_S_out(clk_1_wires[55]),
    .clk_1_N_out(clk_1_wires[54]),
    .clk_1_W_in(clk_1_wires[50]),
    .prog_clk_1_S_out(prog_clk_1_wires[55]),
    .prog_clk_1_N_out(prog_clk_1_wires[54]),
    .prog_clk_1_W_in(prog_clk_1_wires[50]),
    .prog_clk_0_N_in(prog_clk_0_wires[116]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[27]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[27]),
    .SC_OUT_TOP(scff_Wires[71]),
    .SC_IN_BOT(scff_Wires[70]),
    .chanx_left_in(sb_1__1__20_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__27_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__27_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__27_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__27_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__27_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__27_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__27_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__27_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__27_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__27_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__27_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__27_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__27_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__27_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__27_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__27_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__27_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__27_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__27_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__27_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__27_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__1_
  (
    .clk_1_S_out(clk_1_wires[60]),
    .clk_1_N_out(clk_1_wires[59]),
    .clk_1_E_in(clk_1_wires[58]),
    .prog_clk_1_S_out(prog_clk_1_wires[60]),
    .prog_clk_1_N_out(prog_clk_1_wires[59]),
    .prog_clk_1_E_in(prog_clk_1_wires[58]),
    .prog_clk_0_N_in(prog_clk_0_wires[124]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[28]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[28]),
    .SC_OUT_BOT(scff_Wires[89]),
    .SC_IN_TOP(scff_Wires[88]),
    .chanx_left_in(sb_1__1__21_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__28_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__28_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__28_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__28_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__28_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__28_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__28_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__28_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__28_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__28_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__28_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__28_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__28_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__28_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__28_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__28_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__28_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__28_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__28_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__28_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__28_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[127]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[29]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[29]),
    .SC_OUT_BOT(scff_Wires[87]),
    .SC_IN_TOP(scff_Wires[86]),
    .chanx_left_in(sb_1__1__22_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__29_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__29_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__29_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__29_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__29_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__29_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__29_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__29_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__29_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__29_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__29_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__29_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__29_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__29_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__29_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__29_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__29_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__29_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__29_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__29_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__29_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__3_
  (
    .clk_1_S_out(clk_1_wires[67]),
    .clk_1_N_out(clk_1_wires[66]),
    .clk_1_E_in(clk_1_wires[65]),
    .prog_clk_1_S_out(prog_clk_1_wires[67]),
    .prog_clk_1_N_out(prog_clk_1_wires[66]),
    .prog_clk_1_E_in(prog_clk_1_wires[65]),
    .prog_clk_0_N_in(prog_clk_0_wires[130]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[30]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[30]),
    .SC_OUT_BOT(scff_Wires[85]),
    .SC_IN_TOP(scff_Wires[84]),
    .chanx_left_in(sb_1__1__23_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__30_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__30_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__30_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__30_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__30_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__30_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__30_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__30_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__30_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__30_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__30_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__30_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__30_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__30_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__30_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__30_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__30_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__30_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__30_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__30_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__30_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__4_
  (
    .clk_3_E_out(clk_3_wires[2]),
    .clk_3_W_in(clk_3_wires[1]),
    .prog_clk_3_E_out(prog_clk_3_wires[2]),
    .prog_clk_3_W_in(prog_clk_3_wires[1]),
    .prog_clk_0_N_in(prog_clk_0_wires[133]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[31]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[31]),
    .SC_OUT_BOT(scff_Wires[83]),
    .SC_IN_TOP(scff_Wires[82]),
    .chanx_left_in(sb_1__1__24_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__31_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__31_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__31_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__31_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__31_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__31_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__31_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__31_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__31_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__31_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__31_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__31_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__31_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__31_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__31_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__31_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__31_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__31_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__31_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__31_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__31_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__5_
  (
    .clk_1_S_out(clk_1_wires[74]),
    .clk_1_N_out(clk_1_wires[73]),
    .clk_1_E_in(clk_1_wires[72]),
    .prog_clk_1_S_out(prog_clk_1_wires[74]),
    .prog_clk_1_N_out(prog_clk_1_wires[73]),
    .prog_clk_1_E_in(prog_clk_1_wires[72]),
    .prog_clk_0_N_in(prog_clk_0_wires[136]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[32]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[32]),
    .SC_OUT_BOT(scff_Wires[81]),
    .SC_IN_TOP(scff_Wires[80]),
    .chanx_left_in(sb_1__1__25_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__32_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__32_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__32_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__32_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__32_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__32_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__32_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__32_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__32_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__32_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__32_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__32_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__32_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__32_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__32_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__32_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__32_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__32_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__32_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__32_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__32_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[139]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[33]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[33]),
    .SC_OUT_BOT(scff_Wires[79]),
    .SC_IN_TOP(scff_Wires[78]),
    .chanx_left_in(sb_1__1__26_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__33_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__33_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__33_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__33_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__33_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__33_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__33_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__33_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__33_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__33_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__33_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__33_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__33_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__33_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__33_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__33_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__33_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__33_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__33_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__33_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__33_ccff_tail[0])
  );


  cbx_1__1_
  cbx_5__7_
  (
    .clk_1_S_out(clk_1_wires[81]),
    .clk_1_N_out(clk_1_wires[80]),
    .clk_1_E_in(clk_1_wires[79]),
    .prog_clk_1_S_out(prog_clk_1_wires[81]),
    .prog_clk_1_N_out(prog_clk_1_wires[80]),
    .prog_clk_1_E_in(prog_clk_1_wires[79]),
    .prog_clk_0_N_in(prog_clk_0_wires[142]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[34]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[34]),
    .SC_OUT_BOT(scff_Wires[77]),
    .SC_IN_TOP(scff_Wires[76]),
    .chanx_left_in(sb_1__1__27_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__34_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__34_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__34_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__34_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__34_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__34_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__34_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__34_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__34_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__34_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__34_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__34_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__34_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__34_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__34_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__34_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__34_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__34_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__34_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__34_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__34_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__1_
  (
    .clk_1_S_out(clk_1_wires[62]),
    .clk_1_N_out(clk_1_wires[61]),
    .clk_1_W_in(clk_1_wires[57]),
    .prog_clk_1_S_out(prog_clk_1_wires[62]),
    .prog_clk_1_N_out(prog_clk_1_wires[61]),
    .prog_clk_1_W_in(prog_clk_1_wires[57]),
    .prog_clk_0_N_in(prog_clk_0_wires[150]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[35]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[35]),
    .SC_OUT_TOP(scff_Wires[96]),
    .SC_IN_BOT(scff_Wires[95]),
    .chanx_left_in(sb_1__1__28_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__35_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__35_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__35_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__35_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__35_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__35_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__35_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__35_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__35_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__35_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__35_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__35_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__35_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__35_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__35_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__35_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__35_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__35_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__35_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__35_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__35_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__2_
  (
    .clk_2_W_out(clk_2_wires[30]),
    .clk_2_E_in(clk_2_wires[29]),
    .prog_clk_2_W_out(prog_clk_2_wires[30]),
    .prog_clk_2_E_in(prog_clk_2_wires[29]),
    .prog_clk_0_N_in(prog_clk_0_wires[153]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[36]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[36]),
    .SC_OUT_TOP(scff_Wires[98]),
    .SC_IN_BOT(scff_Wires[97]),
    .chanx_left_in(sb_1__1__29_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__36_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__36_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__36_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__36_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__36_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__36_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__36_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__36_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__36_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__36_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__36_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__36_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__36_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__36_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__36_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__36_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__36_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__36_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__36_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__36_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__36_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__3_
  (
    .clk_1_S_out(clk_1_wires[69]),
    .clk_1_N_out(clk_1_wires[68]),
    .clk_1_W_in(clk_1_wires[64]),
    .prog_clk_1_S_out(prog_clk_1_wires[69]),
    .prog_clk_1_N_out(prog_clk_1_wires[68]),
    .prog_clk_1_W_in(prog_clk_1_wires[64]),
    .prog_clk_0_N_in(prog_clk_0_wires[156]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[37]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[37]),
    .SC_OUT_TOP(scff_Wires[100]),
    .SC_IN_BOT(scff_Wires[99]),
    .chanx_left_in(sb_1__1__30_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__37_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__37_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__37_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__37_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__37_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__37_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__37_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__37_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__37_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__37_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__37_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__37_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__37_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__37_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__37_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__37_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__37_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__37_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__37_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__37_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__37_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__4_
  (
    .clk_3_E_out(clk_3_wires[7]),
    .clk_3_W_in(clk_3_wires[6]),
    .prog_clk_3_E_out(prog_clk_3_wires[7]),
    .prog_clk_3_W_in(prog_clk_3_wires[6]),
    .prog_clk_0_N_in(prog_clk_0_wires[159]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[38]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[38]),
    .SC_OUT_TOP(scff_Wires[102]),
    .SC_IN_BOT(scff_Wires[101]),
    .chanx_left_in(sb_1__1__31_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__38_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__38_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__38_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__38_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__38_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__38_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__38_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__38_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__38_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__38_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__38_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__38_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__38_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__38_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__38_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__38_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__38_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__38_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__38_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__38_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__38_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__5_
  (
    .clk_1_S_out(clk_1_wires[76]),
    .clk_1_N_out(clk_1_wires[75]),
    .clk_1_W_in(clk_1_wires[71]),
    .prog_clk_1_S_out(prog_clk_1_wires[76]),
    .prog_clk_1_N_out(prog_clk_1_wires[75]),
    .prog_clk_1_W_in(prog_clk_1_wires[71]),
    .prog_clk_0_N_in(prog_clk_0_wires[162]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[39]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[39]),
    .SC_OUT_TOP(scff_Wires[104]),
    .SC_IN_BOT(scff_Wires[103]),
    .chanx_left_in(sb_1__1__32_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__39_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__39_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__39_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__39_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__39_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__39_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__39_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__39_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__39_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__39_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__39_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__39_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__39_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__39_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__39_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__39_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__39_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__39_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__39_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__39_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__39_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__6_
  (
    .clk_2_W_out(clk_2_wires[43]),
    .clk_2_E_in(clk_2_wires[42]),
    .prog_clk_2_W_out(prog_clk_2_wires[43]),
    .prog_clk_2_E_in(prog_clk_2_wires[42]),
    .prog_clk_0_N_in(prog_clk_0_wires[165]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[40]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[40]),
    .SC_OUT_TOP(scff_Wires[106]),
    .SC_IN_BOT(scff_Wires[105]),
    .chanx_left_in(sb_1__1__33_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__40_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__40_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__40_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__40_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__40_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__40_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__40_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__40_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__40_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__40_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__40_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__40_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__40_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__40_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__40_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__40_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__40_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__40_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__40_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__40_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__40_ccff_tail[0])
  );


  cbx_1__1_
  cbx_6__7_
  (
    .clk_1_S_out(clk_1_wires[83]),
    .clk_1_N_out(clk_1_wires[82]),
    .clk_1_W_in(clk_1_wires[78]),
    .prog_clk_1_S_out(prog_clk_1_wires[83]),
    .prog_clk_1_N_out(prog_clk_1_wires[82]),
    .prog_clk_1_W_in(prog_clk_1_wires[78]),
    .prog_clk_0_N_in(prog_clk_0_wires[168]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[41]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[41]),
    .SC_OUT_TOP(scff_Wires[108]),
    .SC_IN_BOT(scff_Wires[107]),
    .chanx_left_in(sb_1__1__34_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__41_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__41_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__41_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__41_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__41_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__41_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__41_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__41_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__41_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__41_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__41_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__41_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__41_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__41_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__41_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__41_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__41_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__41_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__41_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__41_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__41_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__1_
  (
    .clk_1_S_out(clk_1_wires[88]),
    .clk_1_N_out(clk_1_wires[87]),
    .clk_1_E_in(clk_1_wires[86]),
    .prog_clk_1_S_out(prog_clk_1_wires[88]),
    .prog_clk_1_N_out(prog_clk_1_wires[87]),
    .prog_clk_1_E_in(prog_clk_1_wires[86]),
    .prog_clk_0_N_in(prog_clk_0_wires[176]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[42]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[42]),
    .SC_OUT_BOT(scff_Wires[126]),
    .SC_IN_TOP(scff_Wires[125]),
    .chanx_left_in(sb_1__1__35_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__42_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__42_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__42_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__42_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__42_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__42_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__42_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__42_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__42_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__42_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__42_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__42_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__42_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__42_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__42_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__42_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__42_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__42_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__42_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__42_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__42_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__2_
  (
    .clk_2_E_out(clk_2_wires[28]),
    .clk_2_W_in(clk_2_wires[27]),
    .prog_clk_2_E_out(prog_clk_2_wires[28]),
    .prog_clk_2_W_in(prog_clk_2_wires[27]),
    .prog_clk_0_N_in(prog_clk_0_wires[179]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[43]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[43]),
    .SC_OUT_BOT(scff_Wires[124]),
    .SC_IN_TOP(scff_Wires[123]),
    .chanx_left_in(sb_1__1__36_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__43_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__43_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__43_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__43_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__43_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__43_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__43_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__43_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__43_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__43_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__43_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__43_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__43_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__43_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__43_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__43_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__43_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__43_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__43_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__43_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__43_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__3_
  (
    .clk_1_S_out(clk_1_wires[95]),
    .clk_1_N_out(clk_1_wires[94]),
    .clk_1_E_in(clk_1_wires[93]),
    .prog_clk_1_S_out(prog_clk_1_wires[95]),
    .prog_clk_1_N_out(prog_clk_1_wires[94]),
    .prog_clk_1_E_in(prog_clk_1_wires[93]),
    .prog_clk_0_N_in(prog_clk_0_wires[182]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[44]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[44]),
    .SC_OUT_BOT(scff_Wires[122]),
    .SC_IN_TOP(scff_Wires[121]),
    .chanx_left_in(sb_1__1__37_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__44_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__44_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__44_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__44_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__44_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__44_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__44_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__44_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__44_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__44_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__44_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__44_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__44_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__44_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__44_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__44_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__44_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__44_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__44_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__44_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__44_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[185]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[45]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[45]),
    .SC_OUT_BOT(scff_Wires[120]),
    .SC_IN_TOP(scff_Wires[119]),
    .chanx_left_in(sb_1__1__38_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__45_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__45_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__45_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__45_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__45_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__45_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__45_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__45_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__45_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__45_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__45_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__45_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__45_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__45_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__45_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__45_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__45_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__45_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__45_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__45_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__45_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__5_
  (
    .clk_1_S_out(clk_1_wires[102]),
    .clk_1_N_out(clk_1_wires[101]),
    .clk_1_E_in(clk_1_wires[100]),
    .prog_clk_1_S_out(prog_clk_1_wires[102]),
    .prog_clk_1_N_out(prog_clk_1_wires[101]),
    .prog_clk_1_E_in(prog_clk_1_wires[100]),
    .prog_clk_0_N_in(prog_clk_0_wires[188]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[46]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[46]),
    .SC_OUT_BOT(scff_Wires[118]),
    .SC_IN_TOP(scff_Wires[117]),
    .chanx_left_in(sb_1__1__39_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__46_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__46_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__46_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__46_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__46_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__46_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__46_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__46_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__46_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__46_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__46_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__46_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__46_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__46_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__46_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__46_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__46_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__46_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__46_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__46_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__46_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__6_
  (
    .clk_2_E_out(clk_2_wires[41]),
    .clk_2_W_in(clk_2_wires[40]),
    .prog_clk_2_E_out(prog_clk_2_wires[41]),
    .prog_clk_2_W_in(prog_clk_2_wires[40]),
    .prog_clk_0_N_in(prog_clk_0_wires[191]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[47]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[47]),
    .SC_OUT_BOT(scff_Wires[116]),
    .SC_IN_TOP(scff_Wires[115]),
    .chanx_left_in(sb_1__1__40_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__47_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__47_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__47_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__47_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__47_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__47_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__47_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__47_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__47_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__47_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__47_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__47_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__47_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__47_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__47_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__47_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__47_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__47_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__47_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__47_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__47_ccff_tail[0])
  );


  cbx_1__1_
  cbx_7__7_
  (
    .clk_1_S_out(clk_1_wires[109]),
    .clk_1_N_out(clk_1_wires[108]),
    .clk_1_E_in(clk_1_wires[107]),
    .prog_clk_1_S_out(prog_clk_1_wires[109]),
    .prog_clk_1_N_out(prog_clk_1_wires[108]),
    .prog_clk_1_E_in(prog_clk_1_wires[107]),
    .prog_clk_0_N_in(prog_clk_0_wires[194]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[48]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[48]),
    .SC_OUT_BOT(scff_Wires[114]),
    .SC_IN_TOP(scff_Wires[113]),
    .chanx_left_in(sb_1__1__41_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__1__48_chanx_left_out[0:19]),
    .ccff_head(sb_1__1__48_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__48_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__48_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__48_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__48_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__48_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__48_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__48_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__48_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__48_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__48_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__48_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__48_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__48_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__48_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__48_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__48_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__48_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__48_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__48_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__1_
  (
    .clk_1_S_out(clk_1_wires[90]),
    .clk_1_N_out(clk_1_wires[89]),
    .clk_1_W_in(clk_1_wires[85]),
    .prog_clk_1_S_out(prog_clk_1_wires[90]),
    .prog_clk_1_N_out(prog_clk_1_wires[89]),
    .prog_clk_1_W_in(prog_clk_1_wires[85]),
    .prog_clk_0_N_in(prog_clk_0_wires[202]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[49]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[49]),
    .SC_OUT_TOP(scff_Wires[133]),
    .SC_IN_BOT(scff_Wires[132]),
    .chanx_left_in(sb_1__1__42_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__0_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__49_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__49_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__49_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__49_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__49_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__49_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__49_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__49_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__49_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__49_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__49_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__49_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__49_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__49_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__49_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__49_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__49_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__49_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__49_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__2_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[205]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[50]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[50]),
    .SC_OUT_TOP(scff_Wires[135]),
    .SC_IN_BOT(scff_Wires[134]),
    .chanx_left_in(sb_1__1__43_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__1_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__50_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__50_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__50_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__50_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__50_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__50_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__50_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__50_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__50_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__50_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__50_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__50_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__50_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__50_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__50_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__50_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__50_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__50_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__50_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__3_
  (
    .clk_1_S_out(clk_1_wires[97]),
    .clk_1_N_out(clk_1_wires[96]),
    .clk_1_W_in(clk_1_wires[92]),
    .prog_clk_1_S_out(prog_clk_1_wires[97]),
    .prog_clk_1_N_out(prog_clk_1_wires[96]),
    .prog_clk_1_W_in(prog_clk_1_wires[92]),
    .prog_clk_0_N_in(prog_clk_0_wires[208]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[51]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[51]),
    .SC_OUT_TOP(scff_Wires[137]),
    .SC_IN_BOT(scff_Wires[136]),
    .chanx_left_in(sb_1__1__44_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__2_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__51_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__51_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__51_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__51_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__51_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__51_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__51_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__51_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__51_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__51_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__51_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__51_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__51_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__51_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__51_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__51_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__51_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__51_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__51_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__4_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[211]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[52]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[52]),
    .SC_OUT_TOP(scff_Wires[139]),
    .SC_IN_BOT(scff_Wires[138]),
    .chanx_left_in(sb_1__1__45_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__3_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__52_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__52_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__52_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__52_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__52_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__52_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__52_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__52_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__52_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__52_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__52_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__52_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__52_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__52_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__52_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__52_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__52_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__52_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__52_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__5_
  (
    .clk_1_S_out(clk_1_wires[104]),
    .clk_1_N_out(clk_1_wires[103]),
    .clk_1_W_in(clk_1_wires[99]),
    .prog_clk_1_S_out(prog_clk_1_wires[104]),
    .prog_clk_1_N_out(prog_clk_1_wires[103]),
    .prog_clk_1_W_in(prog_clk_1_wires[99]),
    .prog_clk_0_N_in(prog_clk_0_wires[214]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[53]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[53]),
    .SC_OUT_TOP(scff_Wires[141]),
    .SC_IN_BOT(scff_Wires[140]),
    .chanx_left_in(sb_1__1__46_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__4_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__53_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__53_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__53_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__53_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__53_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__53_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__53_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__53_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__53_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__53_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__53_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__53_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__53_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__53_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__53_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__53_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__53_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__53_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__53_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__6_
  (
    .prog_clk_0_N_in(prog_clk_0_wires[217]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[54]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[54]),
    .SC_OUT_TOP(scff_Wires[143]),
    .SC_IN_BOT(scff_Wires[142]),
    .chanx_left_in(sb_1__1__47_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__5_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__54_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__54_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__54_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__54_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__54_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__54_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__54_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__54_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__54_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__54_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__54_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__54_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__54_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__54_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__54_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__54_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__54_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__54_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__54_ccff_tail[0])
  );


  cbx_1__1_
  cbx_8__7_
  (
    .clk_1_S_out(clk_1_wires[111]),
    .clk_1_N_out(clk_1_wires[110]),
    .clk_1_W_in(clk_1_wires[106]),
    .prog_clk_1_S_out(prog_clk_1_wires[111]),
    .prog_clk_1_N_out(prog_clk_1_wires[110]),
    .prog_clk_1_W_in(prog_clk_1_wires[106]),
    .prog_clk_0_N_in(prog_clk_0_wires[220]),
    .REGOUT_FEEDTHROUGH(regout_feedthrough_wires[55]),
    .REGIN_FEEDTHROUGH(regin_feedthrough_wires[55]),
    .SC_OUT_TOP(scff_Wires[145]),
    .SC_IN_BOT(scff_Wires[144]),
    .chanx_left_in(sb_1__1__48_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__1__6_chanx_left_out[0:19]),
    .ccff_head(sb_8__1__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__1__55_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__1__55_chanx_right_out[0:19]),
    .bottom_grid_pin_0_(cbx_1__1__55_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__1__55_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__1__55_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__1__55_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__1__55_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__1__55_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__1__55_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__1__55_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__1__55_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__1__55_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__1__55_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__1__55_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__1__55_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__1__55_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__1__55_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__1__55_bottom_grid_pin_15_[0]),
    .ccff_tail(cbx_1__1__55_ccff_tail[0])
  );


  cbx_1__2_
  cbx_1__8_
  (
    .prog_clk_0_W_out(prog_clk_0_wires[42]),
    .prog_clk_0_S_in(prog_clk_0_wires[39]),
    .SC_OUT_BOT(scff_Wires[1]),
    .SC_IN_TOP(scff_Wires[0]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_0_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_0_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__0_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_0__8__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__0_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__0_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__0_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__0_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__0_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__0_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__0_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__0_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__0_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__0_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__0_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__0_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__0_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__0_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__0_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__0_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__0_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__0_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__0_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__0_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_0_ccff_tail[0])
  );


  cbx_1__2_
  cbx_2__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[67]),
    .SC_OUT_TOP(scff_Wires[36]),
    .SC_IN_BOT(scff_Wires[35]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_1_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_1_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__1_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__0_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__1_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__1_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__1_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__1_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__1_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__1_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__1_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__1_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__1_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__1_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__1_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__1_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__1_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__1_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__1_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__1_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__1_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__1_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__1_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__1_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__1_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_1_ccff_tail[0])
  );


  cbx_1__2_
  cbx_3__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[93]),
    .SC_OUT_BOT(scff_Wires[38]),
    .SC_IN_TOP(scff_Wires[37]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_2_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_2_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__2_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__1_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__2_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__2_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__2_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__2_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__2_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__2_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__2_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__2_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__2_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__2_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__2_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__2_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__2_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__2_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__2_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__2_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__2_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__2_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__2_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__2_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__2_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_2_ccff_tail[0])
  );


  cbx_1__2_
  cbx_4__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[119]),
    .SC_OUT_TOP(scff_Wires[73]),
    .SC_IN_BOT(scff_Wires[72]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_3_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_3_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__3_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__2_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__3_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__3_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__3_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__3_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__3_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__3_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__3_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__3_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__3_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__3_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__3_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__3_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__3_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__3_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__3_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__3_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__3_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__3_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__3_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__3_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__3_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_3_ccff_tail[0])
  );


  cbx_1__2_
  cbx_5__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[145]),
    .SC_OUT_BOT(scff_Wires[75]),
    .SC_IN_TOP(scff_Wires[74]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_4_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_4_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__4_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__3_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__4_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__4_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__4_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__4_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__4_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__4_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__4_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__4_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__4_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__4_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__4_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__4_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__4_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__4_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__4_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__4_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__4_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__4_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__4_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__4_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__4_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_4_ccff_tail[0])
  );


  cbx_1__2_
  cbx_6__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[171]),
    .SC_OUT_TOP(scff_Wires[110]),
    .SC_IN_BOT(scff_Wires[109]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_5_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_5_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__5_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__4_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__5_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__5_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__5_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__5_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__5_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__5_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__5_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__5_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__5_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__5_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__5_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__5_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__5_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__5_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__5_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__5_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__5_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__5_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__5_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__5_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__5_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_5_ccff_tail[0])
  );


  cbx_1__2_
  cbx_7__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[197]),
    .SC_OUT_BOT(scff_Wires[112]),
    .SC_IN_TOP(scff_Wires[111]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_6_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_6_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__6_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__5_chanx_right_out[0:19]),
    .chanx_right_in(sb_1__8__6_chanx_left_out[0:19]),
    .ccff_head(sb_1__8__6_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__6_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__6_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__6_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__6_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__6_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__6_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__6_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__6_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__6_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__6_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__6_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__6_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__6_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__6_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__6_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__6_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__6_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__6_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__6_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_6_ccff_tail[0])
  );


  cbx_1__2_
  cbx_8__8_
  (
    .prog_clk_0_S_in(prog_clk_0_wires[223]),
    .SC_OUT_TOP(scff_Wires[147]),
    .SC_IN_BOT(scff_Wires[146]),
    .bottom_width_0_height_0__pin_1_lower(grid_io_top_7_bottom_width_0_height_0__pin_1_lower[0]),
    .bottom_width_0_height_0__pin_1_upper(grid_io_top_7_bottom_width_0_height_0__pin_1_upper[0]),
    .bottom_width_0_height_0__pin_0_(cbx_1__8__7_top_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chanx_left_in(sb_1__8__6_chanx_right_out[0:19]),
    .chanx_right_in(sb_8__8__0_chanx_left_out[0:19]),
    .ccff_head(sb_8__8__0_ccff_tail[0]),
    .chanx_left_out(cbx_1__8__7_chanx_left_out[0:19]),
    .chanx_right_out(cbx_1__8__7_chanx_right_out[0:19]),
    .top_grid_pin_0_(cbx_1__8__7_top_grid_pin_0_[0]),
    .bottom_grid_pin_0_(cbx_1__8__7_bottom_grid_pin_0_[0]),
    .bottom_grid_pin_1_(cbx_1__8__7_bottom_grid_pin_1_[0]),
    .bottom_grid_pin_2_(cbx_1__8__7_bottom_grid_pin_2_[0]),
    .bottom_grid_pin_3_(cbx_1__8__7_bottom_grid_pin_3_[0]),
    .bottom_grid_pin_4_(cbx_1__8__7_bottom_grid_pin_4_[0]),
    .bottom_grid_pin_5_(cbx_1__8__7_bottom_grid_pin_5_[0]),
    .bottom_grid_pin_6_(cbx_1__8__7_bottom_grid_pin_6_[0]),
    .bottom_grid_pin_7_(cbx_1__8__7_bottom_grid_pin_7_[0]),
    .bottom_grid_pin_8_(cbx_1__8__7_bottom_grid_pin_8_[0]),
    .bottom_grid_pin_9_(cbx_1__8__7_bottom_grid_pin_9_[0]),
    .bottom_grid_pin_10_(cbx_1__8__7_bottom_grid_pin_10_[0]),
    .bottom_grid_pin_11_(cbx_1__8__7_bottom_grid_pin_11_[0]),
    .bottom_grid_pin_12_(cbx_1__8__7_bottom_grid_pin_12_[0]),
    .bottom_grid_pin_13_(cbx_1__8__7_bottom_grid_pin_13_[0]),
    .bottom_grid_pin_14_(cbx_1__8__7_bottom_grid_pin_14_[0]),
    .bottom_grid_pin_15_(cbx_1__8__7_bottom_grid_pin_15_[0]),
    .ccff_tail(grid_io_top_7_ccff_tail[0])
  );


  cby_0__1_
  cby_0__1_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[3]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_0_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_0_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__0_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__0_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__0_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_0_ccff_tail[0])
  );


  cby_0__1_
  cby_0__2_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[9]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_1_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_1_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__1_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__1_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__1_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_1_ccff_tail[0])
  );


  cby_0__1_
  cby_0__3_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[14]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_2_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_2_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__2_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__2_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__2_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_2_ccff_tail[0])
  );


  cby_0__1_
  cby_0__4_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[19]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_3_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_3_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__3_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__3_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__3_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__3_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_3_ccff_tail[0])
  );


  cby_0__1_
  cby_0__5_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[24]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_4_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_4_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__4_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__4_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__4_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__4_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_4_ccff_tail[0])
  );


  cby_0__1_
  cby_0__6_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[29]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_5_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_5_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__5_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__5_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__5_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__5_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_5_ccff_tail[0])
  );


  cby_0__1_
  cby_0__7_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[34]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_6_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_6_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_0__1__6_chany_bottom_out[0:19]),
    .ccff_head(sb_0__1__6_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__6_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__6_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_6_ccff_tail[0])
  );


  cby_0__1_
  cby_0__8_
  (
    .prog_clk_0_E_in(prog_clk_0_wires[41]),
    .right_width_0_height_0__pin_1_lower(grid_io_left_7_right_width_0_height_0__pin_1_lower[0]),
    .right_width_0_height_0__pin_1_upper(grid_io_left_7_right_width_0_height_0__pin_1_upper[0]),
    .right_width_0_height_0__pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_0__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_0__8__0_chany_bottom_out[0:19]),
    .ccff_head(sb_0__8__0_ccff_tail[0]),
    .chany_bottom_out(cby_0__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_0__1__7_chany_top_out[0:19]),
    .left_grid_pin_0_(cby_0__1__7_left_grid_pin_0_[0]),
    .ccff_tail(grid_io_left_7_ccff_tail[0])
  );


  cby_1__1_
  cby_1__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[2]),
    .prog_clk_0_W_in(prog_clk_0_wires[1]),
    .Test_en_E_in(Test_enWires[18]),
    .Test_en_W_out(Test_enWires[16]),
    .chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_0_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__0_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__0_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__0_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__0_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__0_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__0_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__0_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__0_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__0_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__0_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__0_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__0_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__0_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__0_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__0_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__0_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__0_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__0_ccff_tail[0])
  );


  cby_1__1_
  cby_1__2_
  (
    .clk_2_S_out(clk_2_wires[8]),
    .clk_2_N_in(clk_2_wires[7]),
    .prog_clk_2_S_out(prog_clk_2_wires[8]),
    .prog_clk_2_N_in(prog_clk_2_wires[7]),
    .prog_clk_0_S_out(prog_clk_0_wires[8]),
    .prog_clk_0_W_in(prog_clk_0_wires[7]),
    .Test_en_E_in(Test_enWires[32]),
    .Test_en_W_out(Test_enWires[30]),
    .chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_1_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__1_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__1_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__1_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__1_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__1_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__1_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__1_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__1_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__1_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__1_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__1_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__1_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__1_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__1_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__1_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__1_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__1_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__1_ccff_tail[0])
  );


  cby_1__1_
  cby_1__3_
  (
    .clk_2_N_out(clk_2_wires[6]),
    .clk_2_S_in(clk_2_wires[5]),
    .prog_clk_2_N_out(prog_clk_2_wires[6]),
    .prog_clk_2_S_in(prog_clk_2_wires[5]),
    .prog_clk_0_S_out(prog_clk_0_wires[13]),
    .prog_clk_0_W_in(prog_clk_0_wires[12]),
    .Test_en_E_in(Test_enWires[46]),
    .Test_en_W_out(Test_enWires[44]),
    .chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_2_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__2_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__2_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__2_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__2_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__2_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__2_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__2_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__2_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__2_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__2_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__2_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__2_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__2_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__2_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__2_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__2_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__2_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__2_ccff_tail[0])
  );


  cby_1__1_
  cby_1__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[18]),
    .prog_clk_0_W_in(prog_clk_0_wires[17]),
    .Test_en_E_in(Test_enWires[60]),
    .Test_en_W_out(Test_enWires[58]),
    .chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_3_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__3_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__3_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__3_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__3_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__3_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__3_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__3_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__3_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__3_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__3_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__3_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__3_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__3_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__3_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__3_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__3_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__3_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__3_ccff_tail[0])
  );


  cby_1__1_
  cby_1__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[23]),
    .prog_clk_0_W_in(prog_clk_0_wires[22]),
    .Test_en_E_in(Test_enWires[74]),
    .Test_en_W_out(Test_enWires[72]),
    .chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_4_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__4_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__4_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__4_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__4_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__4_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__4_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__4_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__4_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__4_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__4_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__4_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__4_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__4_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__4_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__4_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__4_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__4_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__4_ccff_tail[0])
  );


  cby_1__1_
  cby_1__6_
  (
    .clk_2_S_out(clk_2_wires[21]),
    .clk_2_N_in(clk_2_wires[20]),
    .prog_clk_2_S_out(prog_clk_2_wires[21]),
    .prog_clk_2_N_in(prog_clk_2_wires[20]),
    .prog_clk_0_S_out(prog_clk_0_wires[28]),
    .prog_clk_0_W_in(prog_clk_0_wires[27]),
    .Test_en_E_in(Test_enWires[88]),
    .Test_en_W_out(Test_enWires[86]),
    .chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_5_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__5_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__5_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__5_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__5_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__5_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__5_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__5_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__5_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__5_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__5_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__5_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__5_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__5_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__5_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__5_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__5_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__5_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__5_ccff_tail[0])
  );


  cby_1__1_
  cby_1__7_
  (
    .clk_2_N_out(clk_2_wires[19]),
    .clk_2_S_in(clk_2_wires[18]),
    .prog_clk_2_N_out(prog_clk_2_wires[19]),
    .prog_clk_2_S_in(prog_clk_2_wires[18]),
    .prog_clk_0_S_out(prog_clk_0_wires[33]),
    .prog_clk_0_W_in(prog_clk_0_wires[32]),
    .Test_en_E_in(Test_enWires[102]),
    .Test_en_W_out(Test_enWires[100]),
    .chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_6_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__6_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__6_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__6_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__6_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__6_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__6_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__6_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__6_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__6_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__6_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__6_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__6_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__6_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__6_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__6_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__6_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__6_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__6_ccff_tail[0])
  );


  cby_1__1_
  cby_1__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[40]),
    .prog_clk_0_S_out(prog_clk_0_wires[38]),
    .prog_clk_0_W_in(prog_clk_0_wires[37]),
    .Test_en_E_in(Test_enWires[116]),
    .Test_en_W_out(Test_enWires[114]),
    .chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_7_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__7_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__7_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__7_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__7_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__7_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__7_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__7_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__7_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__7_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__7_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__7_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__7_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__7_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__7_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__7_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__7_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__7_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__7_ccff_tail[0])
  );


  cby_1__1_
  cby_2__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[45]),
    .prog_clk_0_W_in(prog_clk_0_wires[44]),
    .Test_en_E_in(Test_enWires[20]),
    .Test_en_W_out(Test_enWires[17]),
    .chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_8_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__8_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__8_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__8_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__8_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__8_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__8_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__8_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__8_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__8_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__8_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__8_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__8_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__8_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__8_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__8_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__8_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__8_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__8_ccff_tail[0])
  );


  cby_1__1_
  cby_2__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[48]),
    .prog_clk_0_W_in(prog_clk_0_wires[47]),
    .Test_en_E_in(Test_enWires[34]),
    .Test_en_W_out(Test_enWires[31]),
    .chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_9_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__9_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__9_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__9_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__9_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__9_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__9_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__9_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__9_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__9_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__9_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__9_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__9_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__9_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__9_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__9_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__9_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__9_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__9_ccff_tail[0])
  );


  cby_1__1_
  cby_2__3_
  (
    .clk_3_S_out(clk_3_wires[17]),
    .clk_3_N_in(clk_3_wires[16]),
    .prog_clk_3_S_out(prog_clk_3_wires[17]),
    .prog_clk_3_N_in(prog_clk_3_wires[16]),
    .prog_clk_0_S_out(prog_clk_0_wires[51]),
    .prog_clk_0_W_in(prog_clk_0_wires[50]),
    .Test_en_E_in(Test_enWires[48]),
    .Test_en_W_out(Test_enWires[45]),
    .chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__9_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_10_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__10_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__10_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__10_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__10_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__10_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__10_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__10_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__10_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__10_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__10_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__10_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__10_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__10_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__10_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__10_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__10_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__10_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__10_ccff_tail[0])
  );


  cby_1__1_
  cby_2__4_
  (
    .clk_3_S_out(clk_3_wires[13]),
    .clk_3_N_in(clk_3_wires[12]),
    .prog_clk_3_S_out(prog_clk_3_wires[13]),
    .prog_clk_3_N_in(prog_clk_3_wires[12]),
    .prog_clk_0_S_out(prog_clk_0_wires[54]),
    .prog_clk_0_W_in(prog_clk_0_wires[53]),
    .Test_en_E_in(Test_enWires[62]),
    .Test_en_W_out(Test_enWires[59]),
    .chany_bottom_in(sb_1__1__9_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__10_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_11_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__11_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__11_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__11_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__11_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__11_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__11_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__11_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__11_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__11_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__11_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__11_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__11_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__11_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__11_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__11_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__11_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__11_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__11_ccff_tail[0])
  );


  cby_1__1_
  cby_2__5_
  (
    .clk_3_N_out(clk_3_wires[11]),
    .clk_3_S_in(clk_3_wires[10]),
    .prog_clk_3_N_out(prog_clk_3_wires[11]),
    .prog_clk_3_S_in(prog_clk_3_wires[10]),
    .prog_clk_0_S_out(prog_clk_0_wires[57]),
    .prog_clk_0_W_in(prog_clk_0_wires[56]),
    .Test_en_E_in(Test_enWires[76]),
    .Test_en_W_out(Test_enWires[73]),
    .chany_bottom_in(sb_1__1__10_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__11_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_12_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__12_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__12_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__12_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__12_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__12_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__12_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__12_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__12_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__12_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__12_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__12_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__12_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__12_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__12_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__12_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__12_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__12_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__12_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__12_ccff_tail[0])
  );


  cby_1__1_
  cby_2__6_
  (
    .clk_3_N_out(clk_3_wires[15]),
    .clk_3_S_in(clk_3_wires[14]),
    .prog_clk_3_N_out(prog_clk_3_wires[15]),
    .prog_clk_3_S_in(prog_clk_3_wires[14]),
    .prog_clk_0_S_out(prog_clk_0_wires[60]),
    .prog_clk_0_W_in(prog_clk_0_wires[59]),
    .Test_en_E_in(Test_enWires[90]),
    .Test_en_W_out(Test_enWires[87]),
    .chany_bottom_in(sb_1__1__11_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__12_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_13_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__13_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__13_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__13_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__13_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__13_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__13_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__13_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__13_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__13_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__13_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__13_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__13_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__13_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__13_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__13_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__13_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__13_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__13_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__13_ccff_tail[0])
  );


  cby_1__1_
  cby_2__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[63]),
    .prog_clk_0_W_in(prog_clk_0_wires[62]),
    .Test_en_E_in(Test_enWires[104]),
    .Test_en_W_out(Test_enWires[101]),
    .chany_bottom_in(sb_1__1__12_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__13_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_14_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__14_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__14_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__14_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__14_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__14_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__14_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__14_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__14_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__14_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__14_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__14_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__14_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__14_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__14_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__14_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__14_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__14_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__14_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__14_ccff_tail[0])
  );


  cby_1__1_
  cby_2__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[68]),
    .prog_clk_0_S_out(prog_clk_0_wires[66]),
    .prog_clk_0_W_in(prog_clk_0_wires[65]),
    .Test_en_E_in(Test_enWires[118]),
    .Test_en_W_out(Test_enWires[115]),
    .chany_bottom_in(sb_1__1__13_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_15_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__15_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__15_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__15_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__15_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__15_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__15_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__15_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__15_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__15_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__15_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__15_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__15_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__15_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__15_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__15_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__15_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__15_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__15_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__15_ccff_tail[0])
  );


  cby_1__1_
  cby_3__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[71]),
    .prog_clk_0_W_in(prog_clk_0_wires[70]),
    .Test_en_E_in(Test_enWires[22]),
    .Test_en_W_out(Test_enWires[19]),
    .chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__14_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_16_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__16_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__16_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__16_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__16_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__16_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__16_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__16_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__16_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__16_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__16_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__16_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__16_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__16_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__16_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__16_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__16_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__16_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__16_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__16_ccff_tail[0])
  );


  cby_1__1_
  cby_3__2_
  (
    .clk_2_S_out(clk_2_wires[12]),
    .clk_2_N_in(clk_2_wires[11]),
    .prog_clk_2_S_out(prog_clk_2_wires[12]),
    .prog_clk_2_N_in(prog_clk_2_wires[11]),
    .prog_clk_0_S_out(prog_clk_0_wires[74]),
    .prog_clk_0_W_in(prog_clk_0_wires[73]),
    .Test_en_E_in(Test_enWires[36]),
    .Test_en_W_out(Test_enWires[33]),
    .chany_bottom_in(sb_1__1__14_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__15_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_17_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__17_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__17_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__17_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__17_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__17_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__17_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__17_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__17_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__17_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__17_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__17_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__17_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__17_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__17_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__17_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__17_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__17_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__17_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__17_ccff_tail[0])
  );


  cby_1__1_
  cby_3__3_
  (
    .clk_2_N_out(clk_2_wires[10]),
    .clk_2_S_in(clk_2_wires[9]),
    .prog_clk_2_N_out(prog_clk_2_wires[10]),
    .prog_clk_2_S_in(prog_clk_2_wires[9]),
    .prog_clk_0_S_out(prog_clk_0_wires[77]),
    .prog_clk_0_W_in(prog_clk_0_wires[76]),
    .Test_en_E_in(Test_enWires[50]),
    .Test_en_W_out(Test_enWires[47]),
    .chany_bottom_in(sb_1__1__15_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__16_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_18_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__18_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__18_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__18_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__18_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__18_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__18_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__18_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__18_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__18_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__18_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__18_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__18_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__18_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__18_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__18_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__18_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__18_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__18_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__18_ccff_tail[0])
  );


  cby_1__1_
  cby_3__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[80]),
    .prog_clk_0_W_in(prog_clk_0_wires[79]),
    .Test_en_E_in(Test_enWires[64]),
    .Test_en_W_out(Test_enWires[61]),
    .chany_bottom_in(sb_1__1__16_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__17_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_19_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__19_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__19_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__19_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__19_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__19_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__19_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__19_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__19_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__19_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__19_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__19_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__19_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__19_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__19_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__19_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__19_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__19_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__19_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__19_ccff_tail[0])
  );


  cby_1__1_
  cby_3__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[83]),
    .prog_clk_0_W_in(prog_clk_0_wires[82]),
    .Test_en_E_in(Test_enWires[78]),
    .Test_en_W_out(Test_enWires[75]),
    .chany_bottom_in(sb_1__1__17_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__18_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_20_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__20_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__20_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__20_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__20_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__20_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__20_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__20_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__20_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__20_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__20_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__20_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__20_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__20_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__20_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__20_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__20_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__20_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__20_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__20_ccff_tail[0])
  );


  cby_1__1_
  cby_3__6_
  (
    .clk_2_S_out(clk_2_wires[25]),
    .clk_2_N_in(clk_2_wires[24]),
    .prog_clk_2_S_out(prog_clk_2_wires[25]),
    .prog_clk_2_N_in(prog_clk_2_wires[24]),
    .prog_clk_0_S_out(prog_clk_0_wires[86]),
    .prog_clk_0_W_in(prog_clk_0_wires[85]),
    .Test_en_E_in(Test_enWires[92]),
    .Test_en_W_out(Test_enWires[89]),
    .chany_bottom_in(sb_1__1__18_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__19_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_21_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__21_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__21_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__21_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__21_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__21_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__21_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__21_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__21_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__21_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__21_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__21_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__21_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__21_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__21_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__21_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__21_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__21_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__21_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__21_ccff_tail[0])
  );


  cby_1__1_
  cby_3__7_
  (
    .clk_2_N_out(clk_2_wires[23]),
    .clk_2_S_in(clk_2_wires[22]),
    .prog_clk_2_N_out(prog_clk_2_wires[23]),
    .prog_clk_2_S_in(prog_clk_2_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[89]),
    .prog_clk_0_W_in(prog_clk_0_wires[88]),
    .Test_en_E_in(Test_enWires[106]),
    .Test_en_W_out(Test_enWires[103]),
    .chany_bottom_in(sb_1__1__19_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__20_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_22_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__22_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__22_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__22_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__22_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__22_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__22_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__22_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__22_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__22_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__22_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__22_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__22_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__22_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__22_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__22_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__22_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__22_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__22_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__22_ccff_tail[0])
  );


  cby_1__1_
  cby_3__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[94]),
    .prog_clk_0_S_out(prog_clk_0_wires[92]),
    .prog_clk_0_W_in(prog_clk_0_wires[91]),
    .Test_en_E_in(Test_enWires[120]),
    .Test_en_W_out(Test_enWires[117]),
    .chany_bottom_in(sb_1__1__20_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_23_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__23_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__23_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__23_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__23_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__23_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__23_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__23_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__23_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__23_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__23_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__23_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__23_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__23_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__23_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__23_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__23_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__23_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__23_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__23_ccff_tail[0])
  );


  cby_1__1_
  cby_4__1_
  (
    .clk_3_S_in(clk_3_wires[28]),
    .clk_3_N_out(clk_3_wires[27]),
    .prog_clk_3_S_in(prog_clk_3_wires[28]),
    .prog_clk_3_N_out(prog_clk_3_wires[27]),
    .prog_clk_0_S_out(prog_clk_0_wires[97]),
    .prog_clk_0_W_in(prog_clk_0_wires[96]),
    .Test_en_E_out(Test_enWires[23]),
    .Test_en_W_out(Test_enWires[21]),
    .Test_en_N_out(Test_enWires[2]),
    .Test_en_S_in(Test_enWires[1]),
    .chany_bottom_in(sb_1__0__3_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__21_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_24_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__24_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__24_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__24_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__24_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__24_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__24_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__24_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__24_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__24_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__24_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__24_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__24_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__24_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__24_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__24_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__24_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__24_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__24_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__24_ccff_tail[0])
  );


  cby_1__1_
  cby_4__2_
  (
    .clk_3_S_in(clk_3_wires[30]),
    .clk_3_N_out(clk_3_wires[29]),
    .prog_clk_3_S_in(prog_clk_3_wires[30]),
    .prog_clk_3_N_out(prog_clk_3_wires[29]),
    .prog_clk_0_S_out(prog_clk_0_wires[100]),
    .prog_clk_0_W_in(prog_clk_0_wires[99]),
    .Test_en_E_out(Test_enWires[37]),
    .Test_en_W_out(Test_enWires[35]),
    .Test_en_N_out(Test_enWires[4]),
    .Test_en_S_in(Test_enWires[3]),
    .chany_bottom_in(sb_1__1__21_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__22_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_25_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__25_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__25_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__25_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__25_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__25_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__25_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__25_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__25_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__25_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__25_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__25_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__25_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__25_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__25_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__25_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__25_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__25_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__25_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__25_ccff_tail[0])
  );


  cby_1__1_
  cby_4__3_
  (
    .clk_3_S_in(clk_3_wires[32]),
    .clk_3_N_out(clk_3_wires[31]),
    .prog_clk_3_S_in(prog_clk_3_wires[32]),
    .prog_clk_3_N_out(prog_clk_3_wires[31]),
    .prog_clk_0_S_out(prog_clk_0_wires[103]),
    .prog_clk_0_W_in(prog_clk_0_wires[102]),
    .Test_en_E_out(Test_enWires[51]),
    .Test_en_W_out(Test_enWires[49]),
    .Test_en_N_out(Test_enWires[6]),
    .Test_en_S_in(Test_enWires[5]),
    .chany_bottom_in(sb_1__1__22_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__23_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_26_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__26_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__26_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__26_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__26_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__26_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__26_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__26_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__26_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__26_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__26_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__26_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__26_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__26_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__26_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__26_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__26_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__26_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__26_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__26_ccff_tail[0])
  );


  cby_1__1_
  cby_4__4_
  (
    .clk_3_S_in(clk_3_wires[34]),
    .clk_3_N_out(clk_3_wires[33]),
    .prog_clk_3_S_in(prog_clk_3_wires[34]),
    .prog_clk_3_N_out(prog_clk_3_wires[33]),
    .prog_clk_0_S_out(prog_clk_0_wires[106]),
    .prog_clk_0_W_in(prog_clk_0_wires[105]),
    .Test_en_E_out(Test_enWires[65]),
    .Test_en_W_out(Test_enWires[63]),
    .Test_en_N_out(Test_enWires[8]),
    .Test_en_S_in(Test_enWires[7]),
    .chany_bottom_in(sb_1__1__23_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__24_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_27_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__27_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__27_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__27_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__27_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__27_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__27_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__27_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__27_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__27_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__27_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__27_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__27_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__27_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__27_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__27_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__27_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__27_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__27_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__27_ccff_tail[0])
  );


  cby_1__1_
  cby_4__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[109]),
    .prog_clk_0_W_in(prog_clk_0_wires[108]),
    .Test_en_E_out(Test_enWires[79]),
    .Test_en_W_out(Test_enWires[77]),
    .Test_en_N_out(Test_enWires[10]),
    .Test_en_S_in(Test_enWires[9]),
    .chany_bottom_in(sb_1__1__24_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__25_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_28_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__28_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__28_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__28_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__28_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__28_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__28_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__28_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__28_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__28_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__28_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__28_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__28_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__28_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__28_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__28_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__28_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__28_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__28_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__28_ccff_tail[0])
  );


  cby_1__1_
  cby_4__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[112]),
    .prog_clk_0_W_in(prog_clk_0_wires[111]),
    .Test_en_E_out(Test_enWires[93]),
    .Test_en_W_out(Test_enWires[91]),
    .Test_en_N_out(Test_enWires[12]),
    .Test_en_S_in(Test_enWires[11]),
    .chany_bottom_in(sb_1__1__25_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__26_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_29_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__29_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__29_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__29_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__29_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__29_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__29_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__29_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__29_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__29_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__29_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__29_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__29_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__29_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__29_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__29_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__29_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__29_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__29_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__29_ccff_tail[0])
  );


  cby_1__1_
  cby_4__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[115]),
    .prog_clk_0_W_in(prog_clk_0_wires[114]),
    .Test_en_E_out(Test_enWires[107]),
    .Test_en_W_out(Test_enWires[105]),
    .Test_en_N_out(Test_enWires[14]),
    .Test_en_S_in(Test_enWires[13]),
    .chany_bottom_in(sb_1__1__26_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__27_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_30_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__30_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__30_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__30_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__30_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__30_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__30_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__30_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__30_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__30_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__30_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__30_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__30_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__30_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__30_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__30_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__30_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__30_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__30_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__30_ccff_tail[0])
  );


  cby_1__1_
  cby_4__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[120]),
    .prog_clk_0_S_out(prog_clk_0_wires[118]),
    .prog_clk_0_W_in(prog_clk_0_wires[117]),
    .Test_en_E_out(Test_enWires[121]),
    .Test_en_W_out(Test_enWires[119]),
    .Test_en_S_in(Test_enWires[15]),
    .chany_bottom_in(sb_1__1__27_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_31_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__31_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__31_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__31_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__31_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__31_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__31_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__31_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__31_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__31_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__31_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__31_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__31_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__31_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__31_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__31_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__31_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__31_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__31_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__31_ccff_tail[0])
  );


  cby_1__1_
  cby_5__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[123]),
    .prog_clk_0_W_in(prog_clk_0_wires[122]),
    .Test_en_E_out(Test_enWires[25]),
    .Test_en_W_in(Test_enWires[24]),
    .chany_bottom_in(sb_1__0__4_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__28_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_32_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__32_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__32_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__32_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__32_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__32_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__32_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__32_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__32_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__32_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__32_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__32_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__32_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__32_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__32_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__32_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__32_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__32_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__32_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__32_ccff_tail[0])
  );


  cby_1__1_
  cby_5__2_
  (
    .clk_2_S_out(clk_2_wires[34]),
    .clk_2_N_in(clk_2_wires[33]),
    .prog_clk_2_S_out(prog_clk_2_wires[34]),
    .prog_clk_2_N_in(prog_clk_2_wires[33]),
    .prog_clk_0_S_out(prog_clk_0_wires[126]),
    .prog_clk_0_W_in(prog_clk_0_wires[125]),
    .Test_en_E_out(Test_enWires[39]),
    .Test_en_W_in(Test_enWires[38]),
    .chany_bottom_in(sb_1__1__28_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__29_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_33_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__33_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__33_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__33_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__33_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__33_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__33_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__33_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__33_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__33_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__33_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__33_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__33_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__33_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__33_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__33_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__33_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__33_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__33_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__33_ccff_tail[0])
  );


  cby_1__1_
  cby_5__3_
  (
    .clk_2_N_out(clk_2_wires[32]),
    .clk_2_S_in(clk_2_wires[31]),
    .prog_clk_2_N_out(prog_clk_2_wires[32]),
    .prog_clk_2_S_in(prog_clk_2_wires[31]),
    .prog_clk_0_S_out(prog_clk_0_wires[129]),
    .prog_clk_0_W_in(prog_clk_0_wires[128]),
    .Test_en_E_out(Test_enWires[53]),
    .Test_en_W_in(Test_enWires[52]),
    .chany_bottom_in(sb_1__1__29_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__30_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_34_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__34_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__34_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__34_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__34_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__34_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__34_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__34_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__34_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__34_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__34_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__34_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__34_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__34_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__34_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__34_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__34_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__34_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__34_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__34_ccff_tail[0])
  );


  cby_1__1_
  cby_5__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[132]),
    .prog_clk_0_W_in(prog_clk_0_wires[131]),
    .Test_en_E_out(Test_enWires[67]),
    .Test_en_W_in(Test_enWires[66]),
    .chany_bottom_in(sb_1__1__30_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__31_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_35_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__35_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__35_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__35_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__35_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__35_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__35_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__35_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__35_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__35_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__35_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__35_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__35_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__35_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__35_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__35_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__35_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__35_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__35_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__35_ccff_tail[0])
  );


  cby_1__1_
  cby_5__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[135]),
    .prog_clk_0_W_in(prog_clk_0_wires[134]),
    .Test_en_E_out(Test_enWires[81]),
    .Test_en_W_in(Test_enWires[80]),
    .chany_bottom_in(sb_1__1__31_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__32_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_36_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__36_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__36_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__36_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__36_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__36_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__36_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__36_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__36_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__36_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__36_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__36_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__36_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__36_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__36_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__36_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__36_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__36_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__36_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__36_ccff_tail[0])
  );


  cby_1__1_
  cby_5__6_
  (
    .clk_2_S_out(clk_2_wires[47]),
    .clk_2_N_in(clk_2_wires[46]),
    .prog_clk_2_S_out(prog_clk_2_wires[47]),
    .prog_clk_2_N_in(prog_clk_2_wires[46]),
    .prog_clk_0_S_out(prog_clk_0_wires[138]),
    .prog_clk_0_W_in(prog_clk_0_wires[137]),
    .Test_en_E_out(Test_enWires[95]),
    .Test_en_W_in(Test_enWires[94]),
    .chany_bottom_in(sb_1__1__32_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__33_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_37_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__37_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__37_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__37_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__37_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__37_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__37_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__37_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__37_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__37_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__37_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__37_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__37_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__37_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__37_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__37_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__37_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__37_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__37_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__37_ccff_tail[0])
  );


  cby_1__1_
  cby_5__7_
  (
    .clk_2_N_out(clk_2_wires[45]),
    .clk_2_S_in(clk_2_wires[44]),
    .prog_clk_2_N_out(prog_clk_2_wires[45]),
    .prog_clk_2_S_in(prog_clk_2_wires[44]),
    .prog_clk_0_S_out(prog_clk_0_wires[141]),
    .prog_clk_0_W_in(prog_clk_0_wires[140]),
    .Test_en_E_out(Test_enWires[109]),
    .Test_en_W_in(Test_enWires[108]),
    .chany_bottom_in(sb_1__1__33_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__34_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_38_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__38_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__38_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__38_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__38_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__38_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__38_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__38_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__38_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__38_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__38_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__38_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__38_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__38_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__38_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__38_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__38_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__38_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__38_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__38_ccff_tail[0])
  );


  cby_1__1_
  cby_5__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[146]),
    .prog_clk_0_S_out(prog_clk_0_wires[144]),
    .prog_clk_0_W_in(prog_clk_0_wires[143]),
    .Test_en_E_out(Test_enWires[123]),
    .Test_en_W_in(Test_enWires[122]),
    .chany_bottom_in(sb_1__1__34_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_39_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__39_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__39_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__39_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__39_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__39_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__39_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__39_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__39_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__39_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__39_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__39_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__39_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__39_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__39_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__39_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__39_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__39_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__39_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__39_ccff_tail[0])
  );


  cby_1__1_
  cby_6__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[149]),
    .prog_clk_0_W_in(prog_clk_0_wires[148]),
    .Test_en_E_out(Test_enWires[27]),
    .Test_en_W_in(Test_enWires[26]),
    .chany_bottom_in(sb_1__0__5_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__35_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_40_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__40_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__40_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__40_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__40_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__40_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__40_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__40_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__40_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__40_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__40_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__40_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__40_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__40_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__40_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__40_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__40_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__40_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__40_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__40_ccff_tail[0])
  );


  cby_1__1_
  cby_6__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[152]),
    .prog_clk_0_W_in(prog_clk_0_wires[151]),
    .Test_en_E_out(Test_enWires[41]),
    .Test_en_W_in(Test_enWires[40]),
    .chany_bottom_in(sb_1__1__35_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__36_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_41_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__41_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__41_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__41_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__41_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__41_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__41_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__41_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__41_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__41_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__41_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__41_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__41_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__41_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__41_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__41_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__41_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__41_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__41_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__41_ccff_tail[0])
  );


  cby_1__1_
  cby_6__3_
  (
    .clk_3_S_out(clk_3_wires[25]),
    .clk_3_N_in(clk_3_wires[24]),
    .prog_clk_3_S_out(prog_clk_3_wires[25]),
    .prog_clk_3_N_in(prog_clk_3_wires[24]),
    .prog_clk_0_S_out(prog_clk_0_wires[155]),
    .prog_clk_0_W_in(prog_clk_0_wires[154]),
    .Test_en_E_out(Test_enWires[55]),
    .Test_en_W_in(Test_enWires[54]),
    .chany_bottom_in(sb_1__1__36_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__37_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_42_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__42_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__42_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__42_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__42_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__42_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__42_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__42_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__42_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__42_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__42_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__42_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__42_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__42_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__42_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__42_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__42_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__42_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__42_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__42_ccff_tail[0])
  );


  cby_1__1_
  cby_6__4_
  (
    .clk_3_S_out(clk_3_wires[21]),
    .clk_3_N_in(clk_3_wires[20]),
    .prog_clk_3_S_out(prog_clk_3_wires[21]),
    .prog_clk_3_N_in(prog_clk_3_wires[20]),
    .prog_clk_0_S_out(prog_clk_0_wires[158]),
    .prog_clk_0_W_in(prog_clk_0_wires[157]),
    .Test_en_E_out(Test_enWires[69]),
    .Test_en_W_in(Test_enWires[68]),
    .chany_bottom_in(sb_1__1__37_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__38_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_43_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__43_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__43_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__43_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__43_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__43_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__43_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__43_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__43_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__43_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__43_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__43_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__43_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__43_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__43_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__43_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__43_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__43_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__43_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__43_ccff_tail[0])
  );


  cby_1__1_
  cby_6__5_
  (
    .clk_3_N_out(clk_3_wires[19]),
    .clk_3_S_in(clk_3_wires[18]),
    .prog_clk_3_N_out(prog_clk_3_wires[19]),
    .prog_clk_3_S_in(prog_clk_3_wires[18]),
    .prog_clk_0_S_out(prog_clk_0_wires[161]),
    .prog_clk_0_W_in(prog_clk_0_wires[160]),
    .Test_en_E_out(Test_enWires[83]),
    .Test_en_W_in(Test_enWires[82]),
    .chany_bottom_in(sb_1__1__38_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__39_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_44_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__44_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__44_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__44_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__44_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__44_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__44_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__44_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__44_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__44_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__44_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__44_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__44_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__44_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__44_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__44_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__44_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__44_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__44_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__44_ccff_tail[0])
  );


  cby_1__1_
  cby_6__6_
  (
    .clk_3_N_out(clk_3_wires[23]),
    .clk_3_S_in(clk_3_wires[22]),
    .prog_clk_3_N_out(prog_clk_3_wires[23]),
    .prog_clk_3_S_in(prog_clk_3_wires[22]),
    .prog_clk_0_S_out(prog_clk_0_wires[164]),
    .prog_clk_0_W_in(prog_clk_0_wires[163]),
    .Test_en_E_out(Test_enWires[97]),
    .Test_en_W_in(Test_enWires[96]),
    .chany_bottom_in(sb_1__1__39_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__40_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_45_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__45_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__45_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__45_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__45_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__45_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__45_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__45_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__45_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__45_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__45_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__45_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__45_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__45_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__45_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__45_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__45_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__45_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__45_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__45_ccff_tail[0])
  );


  cby_1__1_
  cby_6__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[167]),
    .prog_clk_0_W_in(prog_clk_0_wires[166]),
    .Test_en_E_out(Test_enWires[111]),
    .Test_en_W_in(Test_enWires[110]),
    .chany_bottom_in(sb_1__1__40_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__41_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_46_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__46_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__46_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__46_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__46_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__46_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__46_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__46_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__46_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__46_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__46_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__46_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__46_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__46_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__46_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__46_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__46_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__46_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__46_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__46_ccff_tail[0])
  );


  cby_1__1_
  cby_6__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[172]),
    .prog_clk_0_S_out(prog_clk_0_wires[170]),
    .prog_clk_0_W_in(prog_clk_0_wires[169]),
    .Test_en_E_out(Test_enWires[125]),
    .Test_en_W_in(Test_enWires[124]),
    .chany_bottom_in(sb_1__1__41_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_47_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__47_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__47_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__47_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__47_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__47_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__47_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__47_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__47_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__47_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__47_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__47_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__47_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__47_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__47_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__47_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__47_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__47_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__47_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__47_ccff_tail[0])
  );


  cby_1__1_
  cby_7__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[175]),
    .prog_clk_0_W_in(prog_clk_0_wires[174]),
    .Test_en_E_out(Test_enWires[29]),
    .Test_en_W_in(Test_enWires[28]),
    .chany_bottom_in(sb_1__0__6_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__42_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_48_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__48_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__48_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__48_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__48_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__48_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__48_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__48_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__48_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__48_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__48_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__48_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__48_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__48_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__48_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__48_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__48_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__48_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__48_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__48_ccff_tail[0])
  );


  cby_1__1_
  cby_7__2_
  (
    .clk_2_S_out(clk_2_wires[38]),
    .clk_2_N_in(clk_2_wires[37]),
    .prog_clk_2_S_out(prog_clk_2_wires[38]),
    .prog_clk_2_N_in(prog_clk_2_wires[37]),
    .prog_clk_0_S_out(prog_clk_0_wires[178]),
    .prog_clk_0_W_in(prog_clk_0_wires[177]),
    .Test_en_E_out(Test_enWires[43]),
    .Test_en_W_in(Test_enWires[42]),
    .chany_bottom_in(sb_1__1__42_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__43_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_49_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__49_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__49_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__49_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__49_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__49_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__49_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__49_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__49_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__49_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__49_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__49_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__49_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__49_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__49_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__49_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__49_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__49_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__49_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__49_ccff_tail[0])
  );


  cby_1__1_
  cby_7__3_
  (
    .clk_2_N_out(clk_2_wires[36]),
    .clk_2_S_in(clk_2_wires[35]),
    .prog_clk_2_N_out(prog_clk_2_wires[36]),
    .prog_clk_2_S_in(prog_clk_2_wires[35]),
    .prog_clk_0_S_out(prog_clk_0_wires[181]),
    .prog_clk_0_W_in(prog_clk_0_wires[180]),
    .Test_en_E_out(Test_enWires[57]),
    .Test_en_W_in(Test_enWires[56]),
    .chany_bottom_in(sb_1__1__43_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__44_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_50_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__50_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__50_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__50_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__50_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__50_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__50_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__50_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__50_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__50_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__50_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__50_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__50_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__50_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__50_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__50_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__50_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__50_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__50_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__50_ccff_tail[0])
  );


  cby_1__1_
  cby_7__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[184]),
    .prog_clk_0_W_in(prog_clk_0_wires[183]),
    .Test_en_E_out(Test_enWires[71]),
    .Test_en_W_in(Test_enWires[70]),
    .chany_bottom_in(sb_1__1__44_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__45_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_51_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__51_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__51_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__51_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__51_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__51_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__51_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__51_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__51_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__51_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__51_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__51_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__51_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__51_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__51_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__51_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__51_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__51_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__51_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__51_ccff_tail[0])
  );


  cby_1__1_
  cby_7__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[187]),
    .prog_clk_0_W_in(prog_clk_0_wires[186]),
    .Test_en_E_out(Test_enWires[85]),
    .Test_en_W_in(Test_enWires[84]),
    .chany_bottom_in(sb_1__1__45_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__46_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_52_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__52_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__52_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__52_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__52_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__52_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__52_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__52_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__52_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__52_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__52_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__52_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__52_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__52_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__52_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__52_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__52_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__52_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__52_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__52_ccff_tail[0])
  );


  cby_1__1_
  cby_7__6_
  (
    .clk_2_S_out(clk_2_wires[51]),
    .clk_2_N_in(clk_2_wires[50]),
    .prog_clk_2_S_out(prog_clk_2_wires[51]),
    .prog_clk_2_N_in(prog_clk_2_wires[50]),
    .prog_clk_0_S_out(prog_clk_0_wires[190]),
    .prog_clk_0_W_in(prog_clk_0_wires[189]),
    .Test_en_E_out(Test_enWires[99]),
    .Test_en_W_in(Test_enWires[98]),
    .chany_bottom_in(sb_1__1__46_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__47_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_53_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__53_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__53_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__53_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__53_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__53_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__53_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__53_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__53_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__53_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__53_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__53_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__53_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__53_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__53_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__53_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__53_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__53_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__53_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__53_ccff_tail[0])
  );


  cby_1__1_
  cby_7__7_
  (
    .clk_2_N_out(clk_2_wires[49]),
    .clk_2_S_in(clk_2_wires[48]),
    .prog_clk_2_N_out(prog_clk_2_wires[49]),
    .prog_clk_2_S_in(prog_clk_2_wires[48]),
    .prog_clk_0_S_out(prog_clk_0_wires[193]),
    .prog_clk_0_W_in(prog_clk_0_wires[192]),
    .Test_en_E_out(Test_enWires[113]),
    .Test_en_W_in(Test_enWires[112]),
    .chany_bottom_in(sb_1__1__47_chany_top_out[0:19]),
    .chany_top_in(sb_1__1__48_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_54_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__54_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__54_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__54_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__54_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__54_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__54_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__54_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__54_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__54_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__54_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__54_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__54_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__54_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__54_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__54_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__54_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__54_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__54_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__54_ccff_tail[0])
  );


  cby_1__1_
  cby_7__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[198]),
    .prog_clk_0_S_out(prog_clk_0_wires[196]),
    .prog_clk_0_W_in(prog_clk_0_wires[195]),
    .Test_en_E_out(Test_enWires[127]),
    .Test_en_W_in(Test_enWires[126]),
    .chany_bottom_in(sb_1__1__48_chany_top_out[0:19]),
    .chany_top_in(sb_1__8__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_55_ccff_tail[0]),
    .chany_bottom_out(cby_1__1__55_chany_bottom_out[0:19]),
    .chany_top_out(cby_1__1__55_chany_top_out[0:19]),
    .left_grid_pin_16_(cby_1__1__55_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_1__1__55_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_1__1__55_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_1__1__55_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_1__1__55_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_1__1__55_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_1__1__55_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_1__1__55_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_1__1__55_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_1__1__55_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_1__1__55_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_1__1__55_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_1__1__55_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_1__1__55_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_1__1__55_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_1__1__55_left_grid_pin_31_[0]),
    .ccff_tail(cby_1__1__55_ccff_tail[0])
  );


  cby_2__1_
  cby_8__1_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[201]),
    .prog_clk_0_W_in(prog_clk_0_wires[200]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_7_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_7_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__0_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__0__0_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_56_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__0_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__0_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__0_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__0_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__0_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__0_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__0_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__0_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__0_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__0_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__0_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__0_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__0_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__0_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__0_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__0_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__0_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__0_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__0_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_7_ccff_tail[0])
  );


  cby_2__1_
  cby_8__2_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[204]),
    .prog_clk_0_W_in(prog_clk_0_wires[203]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_6_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_6_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__1_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__0_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__1_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_57_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__1_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__1_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__1_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__1_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__1_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__1_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__1_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__1_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__1_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__1_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__1_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__1_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__1_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__1_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__1_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__1_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__1_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__1_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__1_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_6_ccff_tail[0])
  );


  cby_2__1_
  cby_8__3_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[207]),
    .prog_clk_0_W_in(prog_clk_0_wires[206]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_5_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_5_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__2_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__1_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__2_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_58_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__2_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__2_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__2_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__2_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__2_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__2_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__2_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__2_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__2_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__2_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__2_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__2_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__2_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__2_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__2_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__2_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__2_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__2_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__2_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_5_ccff_tail[0])
  );


  cby_2__1_
  cby_8__4_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[210]),
    .prog_clk_0_W_in(prog_clk_0_wires[209]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_4_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_4_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__3_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__2_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__3_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_59_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__3_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__3_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__3_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__3_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__3_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__3_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__3_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__3_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__3_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__3_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__3_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__3_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__3_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__3_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__3_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__3_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__3_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__3_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__3_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_4_ccff_tail[0])
  );


  cby_2__1_
  cby_8__5_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[213]),
    .prog_clk_0_W_in(prog_clk_0_wires[212]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_3_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_3_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__4_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__3_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__4_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_60_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__4_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__4_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__4_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__4_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__4_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__4_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__4_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__4_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__4_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__4_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__4_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__4_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__4_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__4_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__4_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__4_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__4_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__4_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__4_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_3_ccff_tail[0])
  );


  cby_2__1_
  cby_8__6_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[216]),
    .prog_clk_0_W_in(prog_clk_0_wires[215]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_2_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_2_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__5_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__4_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__5_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_61_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__5_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__5_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__5_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__5_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__5_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__5_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__5_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__5_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__5_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__5_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__5_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__5_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__5_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__5_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__5_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__5_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__5_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__5_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__5_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_2_ccff_tail[0])
  );


  cby_2__1_
  cby_8__7_
  (
    .prog_clk_0_S_out(prog_clk_0_wires[219]),
    .prog_clk_0_W_in(prog_clk_0_wires[218]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_1_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_1_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__6_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__5_chany_top_out[0:19]),
    .chany_top_in(sb_8__1__6_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_62_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__6_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__6_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__6_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__6_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__6_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__6_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__6_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__6_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__6_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__6_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__6_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__6_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__6_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__6_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__6_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__6_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__6_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__6_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__6_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_1_ccff_tail[0])
  );


  cby_2__1_
  cby_8__8_
  (
    .prog_clk_0_N_out(prog_clk_0_wires[224]),
    .prog_clk_0_S_out(prog_clk_0_wires[222]),
    .prog_clk_0_W_in(prog_clk_0_wires[221]),
    .left_width_0_height_0__pin_1_lower(grid_io_right_0_left_width_0_height_0__pin_1_lower[0]),
    .left_width_0_height_0__pin_1_upper(grid_io_right_0_left_width_0_height_0__pin_1_upper[0]),
    .left_width_0_height_0__pin_0_(cby_8__1__7_right_grid_pin_0_[0]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]),
    .gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]),
    .IO_ISOL_N(IO_ISOL_N[0]),
    .chany_bottom_in(sb_8__1__6_chany_top_out[0:19]),
    .chany_top_in(sb_8__8__0_chany_bottom_out[0:19]),
    .ccff_head(grid_clb_63_ccff_tail[0]),
    .chany_bottom_out(cby_8__1__7_chany_bottom_out[0:19]),
    .chany_top_out(cby_8__1__7_chany_top_out[0:19]),
    .right_grid_pin_0_(cby_8__1__7_right_grid_pin_0_[0]),
    .left_grid_pin_16_(cby_8__1__7_left_grid_pin_16_[0]),
    .left_grid_pin_17_(cby_8__1__7_left_grid_pin_17_[0]),
    .left_grid_pin_18_(cby_8__1__7_left_grid_pin_18_[0]),
    .left_grid_pin_19_(cby_8__1__7_left_grid_pin_19_[0]),
    .left_grid_pin_20_(cby_8__1__7_left_grid_pin_20_[0]),
    .left_grid_pin_21_(cby_8__1__7_left_grid_pin_21_[0]),
    .left_grid_pin_22_(cby_8__1__7_left_grid_pin_22_[0]),
    .left_grid_pin_23_(cby_8__1__7_left_grid_pin_23_[0]),
    .left_grid_pin_24_(cby_8__1__7_left_grid_pin_24_[0]),
    .left_grid_pin_25_(cby_8__1__7_left_grid_pin_25_[0]),
    .left_grid_pin_26_(cby_8__1__7_left_grid_pin_26_[0]),
    .left_grid_pin_27_(cby_8__1__7_left_grid_pin_27_[0]),
    .left_grid_pin_28_(cby_8__1__7_left_grid_pin_28_[0]),
    .left_grid_pin_29_(cby_8__1__7_left_grid_pin_29_[0]),
    .left_grid_pin_30_(cby_8__1__7_left_grid_pin_30_[0]),
    .left_grid_pin_31_(cby_8__1__7_left_grid_pin_31_[0]),
    .ccff_tail(grid_io_right_0_ccff_tail[0])
  );


  direct_interc
  direct_interc_0_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_0_out[0])
  );


  direct_interc
  direct_interc_1_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_1_out[0])
  );


  direct_interc
  direct_interc_2_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_2_out[0])
  );


  direct_interc
  direct_interc_3_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_3_out[0])
  );


  direct_interc
  direct_interc_4_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_4_out[0])
  );


  direct_interc
  direct_interc_5_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_5_out[0])
  );


  direct_interc
  direct_interc_6_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_6_out[0])
  );


  direct_interc
  direct_interc_7_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_7_out[0])
  );


  direct_interc
  direct_interc_8_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_8_out[0])
  );


  direct_interc
  direct_interc_9_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_9_out[0])
  );


  direct_interc
  direct_interc_10_
  (
    .in(grid_clb_12_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_10_out[0])
  );


  direct_interc
  direct_interc_11_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_11_out[0])
  );


  direct_interc
  direct_interc_12_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_12_out[0])
  );


  direct_interc
  direct_interc_13_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_13_out[0])
  );


  direct_interc
  direct_interc_14_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_14_out[0])
  );


  direct_interc
  direct_interc_15_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_15_out[0])
  );


  direct_interc
  direct_interc_16_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_16_out[0])
  );


  direct_interc
  direct_interc_17_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_17_out[0])
  );


  direct_interc
  direct_interc_18_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_18_out[0])
  );


  direct_interc
  direct_interc_19_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_19_out[0])
  );


  direct_interc
  direct_interc_20_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_20_out[0])
  );


  direct_interc
  direct_interc_21_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_21_out[0])
  );


  direct_interc
  direct_interc_22_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_22_out[0])
  );


  direct_interc
  direct_interc_23_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_23_out[0])
  );


  direct_interc
  direct_interc_24_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_24_out[0])
  );


  direct_interc
  direct_interc_25_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_25_out[0])
  );


  direct_interc
  direct_interc_26_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_26_out[0])
  );


  direct_interc
  direct_interc_27_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_27_out[0])
  );


  direct_interc
  direct_interc_28_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_28_out[0])
  );


  direct_interc
  direct_interc_29_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_29_out[0])
  );


  direct_interc
  direct_interc_30_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_30_out[0])
  );


  direct_interc
  direct_interc_31_
  (
    .in(grid_clb_36_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_31_out[0])
  );


  direct_interc
  direct_interc_32_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_32_out[0])
  );


  direct_interc
  direct_interc_33_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_33_out[0])
  );


  direct_interc
  direct_interc_34_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_34_out[0])
  );


  direct_interc
  direct_interc_35_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_35_out[0])
  );


  direct_interc
  direct_interc_36_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_36_out[0])
  );


  direct_interc
  direct_interc_37_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_37_out[0])
  );


  direct_interc
  direct_interc_38_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_38_out[0])
  );


  direct_interc
  direct_interc_39_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_39_out[0])
  );


  direct_interc
  direct_interc_40_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_40_out[0])
  );


  direct_interc
  direct_interc_41_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_41_out[0])
  );


  direct_interc
  direct_interc_42_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_42_out[0])
  );


  direct_interc
  direct_interc_43_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_43_out[0])
  );


  direct_interc
  direct_interc_44_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_44_out[0])
  );


  direct_interc
  direct_interc_45_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_45_out[0])
  );


  direct_interc
  direct_interc_46_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_46_out[0])
  );


  direct_interc
  direct_interc_47_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_47_out[0])
  );


  direct_interc
  direct_interc_48_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_48_out[0])
  );


  direct_interc
  direct_interc_49_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_49_out[0])
  );


  direct_interc
  direct_interc_50_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_50_out[0])
  );


  direct_interc
  direct_interc_51_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_51_out[0])
  );


  direct_interc
  direct_interc_52_
  (
    .in(grid_clb_60_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_52_out[0])
  );


  direct_interc
  direct_interc_53_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_53_out[0])
  );


  direct_interc
  direct_interc_54_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_54_out[0])
  );


  direct_interc
  direct_interc_55_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_50_[0]),
    .out(direct_interc_55_out[0])
  );


  direct_interc
  direct_interc_56_
  (
    .in(grid_clb_1_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_56_out[0])
  );


  direct_interc
  direct_interc_57_
  (
    .in(grid_clb_2_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_57_out[0])
  );


  direct_interc
  direct_interc_58_
  (
    .in(grid_clb_3_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_58_out[0])
  );


  direct_interc
  direct_interc_59_
  (
    .in(grid_clb_4_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_59_out[0])
  );


  direct_interc
  direct_interc_60_
  (
    .in(grid_clb_5_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_60_out[0])
  );


  direct_interc
  direct_interc_61_
  (
    .in(grid_clb_6_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_61_out[0])
  );


  direct_interc
  direct_interc_62_
  (
    .in(grid_clb_7_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_62_out[0])
  );


  direct_interc
  direct_interc_63_
  (
    .in(grid_clb_9_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_63_out[0])
  );


  direct_interc
  direct_interc_64_
  (
    .in(grid_clb_10_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_64_out[0])
  );


  direct_interc
  direct_interc_65_
  (
    .in(grid_clb_11_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_65_out[0])
  );


  direct_interc
  direct_interc_66_
  (
    .in(grid_clb_12_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_66_out[0])
  );


  direct_interc
  direct_interc_67_
  (
    .in(grid_clb_13_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_67_out[0])
  );


  direct_interc
  direct_interc_68_
  (
    .in(grid_clb_14_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_68_out[0])
  );


  direct_interc
  direct_interc_69_
  (
    .in(grid_clb_15_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_69_out[0])
  );


  direct_interc
  direct_interc_70_
  (
    .in(grid_clb_17_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_70_out[0])
  );


  direct_interc
  direct_interc_71_
  (
    .in(grid_clb_18_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_71_out[0])
  );


  direct_interc
  direct_interc_72_
  (
    .in(grid_clb_19_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_72_out[0])
  );


  direct_interc
  direct_interc_73_
  (
    .in(grid_clb_20_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_73_out[0])
  );


  direct_interc
  direct_interc_74_
  (
    .in(grid_clb_21_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_74_out[0])
  );


  direct_interc
  direct_interc_75_
  (
    .in(grid_clb_22_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_75_out[0])
  );


  direct_interc
  direct_interc_76_
  (
    .in(grid_clb_23_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_76_out[0])
  );


  direct_interc
  direct_interc_77_
  (
    .in(grid_clb_25_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_77_out[0])
  );


  direct_interc
  direct_interc_78_
  (
    .in(grid_clb_26_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_78_out[0])
  );


  direct_interc
  direct_interc_79_
  (
    .in(grid_clb_27_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_79_out[0])
  );


  direct_interc
  direct_interc_80_
  (
    .in(grid_clb_28_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_80_out[0])
  );


  direct_interc
  direct_interc_81_
  (
    .in(grid_clb_29_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_81_out[0])
  );


  direct_interc
  direct_interc_82_
  (
    .in(grid_clb_30_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_82_out[0])
  );


  direct_interc
  direct_interc_83_
  (
    .in(grid_clb_31_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_83_out[0])
  );


  direct_interc
  direct_interc_84_
  (
    .in(grid_clb_33_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_84_out[0])
  );


  direct_interc
  direct_interc_85_
  (
    .in(grid_clb_34_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_85_out[0])
  );


  direct_interc
  direct_interc_86_
  (
    .in(grid_clb_35_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_86_out[0])
  );


  direct_interc
  direct_interc_87_
  (
    .in(grid_clb_36_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_87_out[0])
  );


  direct_interc
  direct_interc_88_
  (
    .in(grid_clb_37_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_88_out[0])
  );


  direct_interc
  direct_interc_89_
  (
    .in(grid_clb_38_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_89_out[0])
  );


  direct_interc
  direct_interc_90_
  (
    .in(grid_clb_39_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_90_out[0])
  );


  direct_interc
  direct_interc_91_
  (
    .in(grid_clb_41_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_91_out[0])
  );


  direct_interc
  direct_interc_92_
  (
    .in(grid_clb_42_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_92_out[0])
  );


  direct_interc
  direct_interc_93_
  (
    .in(grid_clb_43_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_93_out[0])
  );


  direct_interc
  direct_interc_94_
  (
    .in(grid_clb_44_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_94_out[0])
  );


  direct_interc
  direct_interc_95_
  (
    .in(grid_clb_45_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_95_out[0])
  );


  direct_interc
  direct_interc_96_
  (
    .in(grid_clb_46_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_96_out[0])
  );


  direct_interc
  direct_interc_97_
  (
    .in(grid_clb_47_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_97_out[0])
  );


  direct_interc
  direct_interc_98_
  (
    .in(grid_clb_49_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_98_out[0])
  );


  direct_interc
  direct_interc_99_
  (
    .in(grid_clb_50_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_99_out[0])
  );


  direct_interc
  direct_interc_100_
  (
    .in(grid_clb_51_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_100_out[0])
  );


  direct_interc
  direct_interc_101_
  (
    .in(grid_clb_52_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_101_out[0])
  );


  direct_interc
  direct_interc_102_
  (
    .in(grid_clb_53_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_102_out[0])
  );


  direct_interc
  direct_interc_103_
  (
    .in(grid_clb_54_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_103_out[0])
  );


  direct_interc
  direct_interc_104_
  (
    .in(grid_clb_55_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_104_out[0])
  );


  direct_interc
  direct_interc_105_
  (
    .in(grid_clb_57_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_105_out[0])
  );


  direct_interc
  direct_interc_106_
  (
    .in(grid_clb_58_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_106_out[0])
  );


  direct_interc
  direct_interc_107_
  (
    .in(grid_clb_59_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_107_out[0])
  );


  direct_interc
  direct_interc_108_
  (
    .in(grid_clb_60_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_108_out[0])
  );


  direct_interc
  direct_interc_109_
  (
    .in(grid_clb_61_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_109_out[0])
  );


  direct_interc
  direct_interc_110_
  (
    .in(grid_clb_62_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_110_out[0])
  );


  direct_interc
  direct_interc_111_
  (
    .in(grid_clb_63_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_111_out[0])
  );


  direct_interc
  direct_interc_112_
  (
    .in(grid_clb_0_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_112_out[0])
  );


  direct_interc
  direct_interc_113_
  (
    .in(grid_clb_8_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_113_out[0])
  );


  direct_interc
  direct_interc_114_
  (
    .in(grid_clb_16_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_114_out[0])
  );


  direct_interc
  direct_interc_115_
  (
    .in(grid_clb_24_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_115_out[0])
  );


  direct_interc
  direct_interc_116_
  (
    .in(grid_clb_32_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_116_out[0])
  );


  direct_interc
  direct_interc_117_
  (
    .in(grid_clb_40_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_117_out[0])
  );


  direct_interc
  direct_interc_118_
  (
    .in(grid_clb_48_bottom_width_0_height_0__pin_51_[0]),
    .out(direct_interc_118_out[0])
  );


endmodule

