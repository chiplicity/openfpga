* NGSPICE file created from cby_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

.subckt cby_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_grid_pin_0_ left_grid_pin_10_ left_grid_pin_12_ left_grid_pin_14_ left_grid_pin_2_
+ left_grid_pin_4_ left_grid_pin_6_ left_grid_pin_8_ right_grid_pin_3_ right_grid_pin_7_
+ vpwr vgnd
XFILLER_3_23 vpwr vgnd scs8hd_fill_2
XFILLER_3_12 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_114 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vpwr vgnd scs8hd_fill_2
XFILLER_12_43 vpwr vgnd scs8hd_fill_2
XFILLER_12_87 vgnd vpwr scs8hd_decap_4
XANTENNA__108__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _116_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_131_ _139_/A _133_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_42 vpwr vgnd scs8hd_fill_2
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_23_75 vpwr vgnd scs8hd_fill_2
XFILLER_23_97 vpwr vgnd scs8hd_fill_2
X_062_ address[1] address[2] address[0] _062_/X vgnd vpwr scs8hd_or3_4
XFILLER_2_132 vgnd vpwr scs8hd_decap_12
XANTENNA__110__C _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
XFILLER_9_66 vgnd vpwr scs8hd_decap_3
XANTENNA__119__A _119_/A vgnd vpwr scs8hd_diode_2
XFILLER_50_3 vgnd vpwr scs8hd_decap_12
XFILLER_47_117 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_0_.latch/Q mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_50_84 vgnd vpwr scs8hd_decap_3
X_114_ _073_/X _115_/B _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_117 vgnd vpwr scs8hd_decap_8
XFILLER_38_128 vgnd vpwr scs8hd_decap_12
XANTENNA__121__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_61_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_19 vpwr vgnd scs8hd_fill_2
XFILLER_29_117 vgnd vpwr scs8hd_decap_4
XFILLER_52_131 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_2.LATCH_1_.latch data_in mem_right_ipin_2.LATCH_1_.latch/Q _097_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_54 vgnd vpwr scs8hd_decap_8
XFILLER_20_65 vpwr vgnd scs8hd_fill_2
XFILLER_29_85 vpwr vgnd scs8hd_fill_2
XFILLER_35_109 vpwr vgnd scs8hd_fill_2
XANTENNA__116__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _132_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_4.LATCH_4_.latch data_in mem_right_ipin_4.LATCH_4_.latch/Q _113_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XFILLER_31_86 vpwr vgnd scs8hd_fill_2
XFILLER_56_83 vpwr vgnd scs8hd_fill_2
XFILLER_56_72 vpwr vgnd scs8hd_fill_2
XFILLER_16_131 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_145 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_42_52 vgnd vpwr scs8hd_decap_6
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XFILLER_6_108 vgnd vpwr scs8hd_decap_12
XFILLER_10_126 vgnd vpwr scs8hd_decap_12
XFILLER_12_55 vpwr vgnd scs8hd_fill_2
XFILLER_37_30 vpwr vgnd scs8hd_fill_2
XFILLER_53_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _175_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__124__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _132_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_130_ _138_/A _133_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_48_51 vgnd vpwr scs8hd_decap_3
XFILLER_2_144 vpwr vgnd scs8hd_fill_2
XFILLER_64_94 vgnd vpwr scs8hd_decap_12
XFILLER_0_36 vgnd vpwr scs8hd_decap_3
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__135__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_43_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_6
XFILLER_18_54 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _145_/A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_42 vgnd vpwr scs8hd_decap_12
X_113_ _071_/X _115_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_5.LATCH_0_.latch data_in mem_right_ipin_5.LATCH_0_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_61_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_20_88 vgnd vpwr scs8hd_decap_4
XFILLER_45_52 vgnd vpwr scs8hd_decap_3
XFILLER_43_132 vpwr vgnd scs8hd_fill_2
XFILLER_61_95 vpwr vgnd scs8hd_fill_2
XFILLER_61_51 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_7.LATCH_3_.latch data_in mem_right_ipin_7.LATCH_3_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_24 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__B _133_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_6_79 vgnd vpwr scs8hd_decap_8
XFILLER_34_143 vgnd vpwr scs8hd_decap_3
XFILLER_15_11 vgnd vpwr scs8hd_decap_3
XFILLER_15_55 vgnd vpwr scs8hd_fill_1
XFILLER_15_66 vgnd vpwr scs8hd_fill_1
XFILLER_31_54 vgnd vpwr scs8hd_decap_4
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_143 vgnd vpwr scs8hd_decap_3
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_31_135 vgnd vpwr scs8hd_decap_8
XANTENNA__143__A _067_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_36 vgnd vpwr scs8hd_decap_3
XANTENNA__138__A _138_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_0_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_138 vgnd vpwr scs8hd_decap_8
XFILLER_37_53 vgnd vpwr scs8hd_decap_4
XFILLER_37_75 vgnd vpwr scs8hd_fill_1
XFILLER_53_52 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_127 vpwr vgnd scs8hd_fill_2
XFILLER_23_11 vgnd vpwr scs8hd_fill_1
XFILLER_23_88 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vpwr vgnd scs8hd_fill_2
XFILLER_48_63 vpwr vgnd scs8hd_fill_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
X_189_ chany_bottom_in[8] chany_top_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__135__B _127_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vpwr scs8hd_fill_1
XFILLER_34_54 vpwr vgnd scs8hd_fill_2
X_112_ _156_/A _115_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_95 vpwr vgnd scs8hd_fill_2
XFILLER_59_62 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_46_130 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _146_/A vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_7_ vgnd vpwr scs8hd_inv_1
XFILLER_37_130 vgnd vpwr scs8hd_decap_4
XFILLER_37_141 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_23 vgnd vpwr scs8hd_decap_4
XFILLER_29_98 vpwr vgnd scs8hd_fill_2
XFILLER_45_86 vpwr vgnd scs8hd_fill_2
XFILLER_45_75 vgnd vpwr scs8hd_decap_4
XFILLER_43_144 vpwr vgnd scs8hd_fill_2
XFILLER_61_74 vgnd vpwr scs8hd_decap_3
XFILLER_6_58 vgnd vpwr scs8hd_decap_8
XFILLER_6_47 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _154_/C vgnd vpwr scs8hd_diode_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_103 vpwr vgnd scs8hd_fill_2
XANTENNA__143__B _101_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_87 vgnd vpwr scs8hd_decap_4
XFILLER_42_76 vpwr vgnd scs8hd_fill_2
XFILLER_42_32 vpwr vgnd scs8hd_fill_2
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_0.LATCH_4_.latch data_in mem_right_ipin_0.LATCH_4_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__138__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_ipin_0.LATCH_3_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__A _166_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_68 vpwr vgnd scs8hd_fill_2
XFILLER_12_79 vpwr vgnd scs8hd_fill_2
XFILLER_53_75 vgnd vpwr scs8hd_decap_4
XFILLER_5_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _176_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_86 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_64_63 vgnd vpwr scs8hd_decap_12
X_188_ chany_top_in[0] chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__135__C _066_/C vgnd vpwr scs8hd_diode_2
XFILLER_29_3 vgnd vpwr scs8hd_decap_6
XFILLER_55_131 vgnd vpwr scs8hd_decap_12
XFILLER_47_109 vpwr vgnd scs8hd_fill_2
XFILLER_18_23 vgnd vpwr scs8hd_decap_4
XFILLER_18_67 vgnd vpwr scs8hd_decap_4
XFILLER_50_32 vgnd vpwr scs8hd_decap_12
X_111_ _110_/X _115_/B vgnd vpwr scs8hd_buf_1
XFILLER_61_123 vgnd vpwr scs8hd_decap_12
XFILLER_46_142 vgnd vpwr scs8hd_decap_4
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_109 vpwr vgnd scs8hd_fill_2
XFILLER_1_70 vgnd vpwr scs8hd_decap_4
XANTENNA__072__A _071_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_35 vpwr vgnd scs8hd_fill_2
XFILLER_29_11 vgnd vpwr scs8hd_decap_3
XFILLER_29_22 vgnd vpwr scs8hd_decap_3
XFILLER_43_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_55 vgnd vpwr scs8hd_decap_4
XFILLER_29_77 vpwr vgnd scs8hd_fill_2
XFILLER_61_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_0_.latch/Q mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_34_123 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_0_.latch data_in mem_right_ipin_1.LATCH_0_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_104 vpwr vgnd scs8hd_fill_2
XFILLER_15_24 vgnd vpwr scs8hd_fill_1
XFILLER_25_134 vgnd vpwr scs8hd_fill_1
XFILLER_25_145 vgnd vpwr scs8hd_fill_1
XANTENNA__067__A _066_/X vgnd vpwr scs8hd_diode_2
XFILLER_31_45 vgnd vpwr scs8hd_decap_3
XFILLER_56_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_115 vgnd vpwr scs8hd_decap_6
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _161_/C vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_104 vgnd vpwr scs8hd_decap_8
XFILLER_22_115 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_3.LATCH_3_.latch data_in mem_right_ipin_3.LATCH_3_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_67 vgnd vpwr scs8hd_decap_3
XFILLER_42_11 vgnd vpwr scs8hd_decap_3
XFILLER_59_3 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__064__B _134_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_47 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.INVTX1_3_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_22 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_88 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _164_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_46 vpwr vgnd scs8hd_fill_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A _132_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_43 vpwr vgnd scs8hd_fill_2
XFILLER_48_32 vgnd vpwr scs8hd_decap_8
XFILLER_64_75 vgnd vpwr scs8hd_decap_12
XFILLER_9_15 vgnd vpwr scs8hd_decap_4
X_187_ chany_top_in[1] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_13_90 vgnd vpwr scs8hd_decap_3
XANTENNA__135__D _101_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_4_.latch data_in mem_left_ipin_0.LATCH_4_.latch/Q _159_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_143 vgnd vpwr scs8hd_decap_3
X_110_ _065_/Y address[3] _099_/X _110_/X vgnd vpwr scs8hd_or3_4
XFILLER_34_89 vgnd vpwr scs8hd_fill_1
XFILLER_59_53 vpwr vgnd scs8hd_fill_2
XFILLER_61_135 vgnd vpwr scs8hd_decap_8
XFILLER_41_3 vgnd vpwr scs8hd_decap_8
XFILLER_37_121 vgnd vpwr scs8hd_fill_1
XFILLER_52_102 vpwr vgnd scs8hd_fill_2
XANTENNA__072__B _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_20_69 vpwr vgnd scs8hd_fill_2
XFILLER_29_34 vgnd vpwr scs8hd_decap_3
XFILLER_6_16 vgnd vpwr scs8hd_decap_8
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_34_102 vpwr vgnd scs8hd_fill_2
XFILLER_34_135 vgnd vpwr scs8hd_decap_8
XANTENNA__157__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_47 vpwr vgnd scs8hd_fill_2
XFILLER_15_58 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_6.LATCH_2_.latch data_in mem_right_ipin_6.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_56_32 vgnd vpwr scs8hd_decap_12
XFILLER_56_87 vpwr vgnd scs8hd_fill_2
XFILLER_56_76 vpwr vgnd scs8hd_fill_2
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_102 vgnd vpwr scs8hd_decap_8
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_127 vgnd vpwr scs8hd_decap_12
XANTENNA__078__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_79 vgnd vpwr scs8hd_decap_3
XFILLER_42_23 vgnd vpwr scs8hd_decap_8
XANTENNA__154__C _154_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA__080__B _076_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_34 vpwr vgnd scs8hd_fill_2
XFILLER_37_78 vgnd vpwr scs8hd_fill_1
XFILLER_53_99 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
Xmem_left_ipin_1.LATCH_0_.latch data_in _146_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _177_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__149__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_59_108 vpwr vgnd scs8hd_fill_2
XANTENNA__181__A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _090_/Y vgnd vpwr scs8hd_diode_2
XFILLER_64_87 vgnd vpwr scs8hd_decap_6
XFILLER_64_32 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_0_.latch/Q mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_186_ chany_top_in[2] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
Xmux_right_ipin_3.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__086__A _073_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_68 vpwr vgnd scs8hd_fill_2
XFILLER_34_79 vpwr vgnd scs8hd_fill_2
XFILLER_50_89 vgnd vpwr scs8hd_decap_3
XFILLER_50_67 vpwr vgnd scs8hd_fill_2
XFILLER_1_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_169_ _166_/A _133_/A _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_43_136 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_144 vpwr vgnd scs8hd_fill_2
XFILLER_61_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_90 vgnd vpwr scs8hd_decap_4
XFILLER_19_111 vgnd vpwr scs8hd_fill_1
XANTENNA__157__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_117 vpwr vgnd scs8hd_fill_2
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XFILLER_40_128 vgnd vpwr scs8hd_decap_12
XFILLER_31_58 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_56_44 vgnd vpwr scs8hd_decap_6
XPHY_120 vgnd vpwr scs8hd_decap_3
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_91 vpwr vgnd scs8hd_fill_2
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_139 vgnd vpwr scs8hd_decap_6
XANTENNA__078__B _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _071_/X vgnd vpwr scs8hd_diode_2
XFILLER_26_47 vgnd vpwr scs8hd_decap_4
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _146_/A mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__089__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_56 vgnd vpwr scs8hd_decap_3
XFILLER_5_135 vgnd vpwr scs8hd_decap_8
XFILLER_5_102 vgnd vpwr scs8hd_decap_12
XFILLER_64_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_50 vpwr vgnd scs8hd_fill_2
XANTENNA__091__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_48_67 vpwr vgnd scs8hd_fill_2
XFILLER_64_44 vgnd vpwr scs8hd_decap_12
X_185_ chany_top_in[3] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_64_145 vgnd vpwr scs8hd_fill_1
XANTENNA__192__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__086__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_50_46 vgnd vpwr scs8hd_decap_12
XFILLER_34_58 vgnd vpwr scs8hd_fill_1
XFILLER_59_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_7.LATCH_3_.latch/Q mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
X_168_ _168_/A _133_/A vgnd vpwr scs8hd_buf_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_099_ _090_/Y address[6] _066_/C _099_/X vgnd vpwr scs8hd_or3_4
XANTENNA__187__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_37_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_1.INVTX1_3_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XFILLER_45_57 vpwr vgnd scs8hd_fill_2
XFILLER_45_35 vpwr vgnd scs8hd_fill_2
XFILLER_45_24 vpwr vgnd scs8hd_fill_2
XANTENNA__097__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XFILLER_25_126 vgnd vpwr scs8hd_decap_8
XFILLER_25_137 vgnd vpwr scs8hd_decap_8
XFILLER_31_26 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_121 vgnd vpwr scs8hd_decap_3
XPHY_110 vgnd vpwr scs8hd_decap_3
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_107 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_0_.latch/Q mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_58 vgnd vpwr scs8hd_fill_1
XFILLER_42_36 vgnd vpwr scs8hd_decap_3
XFILLER_13_107 vgnd vpwr scs8hd_decap_12
XANTENNA__094__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_19 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_2.LATCH_2_.latch data_in mem_right_ipin_2.LATCH_2_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_80 vgnd vpwr scs8hd_decap_8
XANTENNA__195__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_53_79 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_114 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_4.LATCH_5_.latch data_in mem_right_ipin_4.LATCH_5_.latch/Q _112_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _178_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_57_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_27 vpwr vgnd scs8hd_fill_2
XFILLER_3_8 vpwr vgnd scs8hd_fill_2
XANTENNA__091__C _154_/C vgnd vpwr scs8hd_diode_2
XFILLER_58_121 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_1_.latch/Q mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_64_56 vgnd vpwr scs8hd_decap_6
X_184_ chany_top_in[4] chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_13_71 vgnd vpwr scs8hd_decap_4
XFILLER_13_82 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_49_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_113 vpwr vgnd scs8hd_fill_2
XFILLER_18_38 vgnd vpwr scs8hd_fill_1
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XFILLER_46_102 vgnd vpwr scs8hd_decap_8
XFILLER_24_70 vpwr vgnd scs8hd_fill_2
X_098_ _117_/A _094_/B _098_/Y vgnd vpwr scs8hd_nor2_4
X_167_ address[1] address[2] _161_/C _168_/A vgnd vpwr scs8hd_or3_4
XFILLER_37_113 vpwr vgnd scs8hd_fill_2
XFILLER_1_85 vpwr vgnd scs8hd_fill_2
XFILLER_20_39 vpwr vgnd scs8hd_fill_2
XFILLER_43_116 vgnd vpwr scs8hd_decap_4
XANTENNA__097__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_50 vgnd vpwr scs8hd_decap_8
XFILLER_19_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_28 vpwr vgnd scs8hd_fill_2
XFILLER_56_57 vgnd vpwr scs8hd_decap_4
XPHY_100 vgnd vpwr scs8hd_decap_3
XPHY_122 vgnd vpwr scs8hd_decap_3
XPHY_111 vgnd vpwr scs8hd_decap_3
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_82 vgnd vpwr scs8hd_decap_3
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_84 vpwr vgnd scs8hd_fill_2
XFILLER_7_62 vgnd vpwr scs8hd_decap_4
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_5.LATCH_1_.latch data_in mem_right_ipin_5.LATCH_1_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_119 vgnd vpwr scs8hd_decap_3
XFILLER_16_82 vgnd vpwr scs8hd_decap_8
XFILLER_12_141 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_7.LATCH_4_.latch data_in mem_right_ipin_7.LATCH_4_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_ipin_6.LATCH_3_.latch/Q mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_4
XFILLER_53_47 vgnd vpwr scs8hd_decap_3
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_96 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_58_133 vgnd vpwr scs8hd_decap_12
XFILLER_48_47 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _171_/HI _145_/Y mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_19 vgnd vpwr scs8hd_fill_1
X_183_ chany_top_in[5] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_64_125 vgnd vpwr scs8hd_decap_12
XFILLER_38_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_50_15 vgnd vpwr scs8hd_decap_12
XFILLER_59_79 vpwr vgnd scs8hd_fill_2
XFILLER_59_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
X_166_ _166_/A _132_/A _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _116_/A _094_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_0_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_52_106 vgnd vpwr scs8hd_decap_4
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XFILLER_45_15 vgnd vpwr scs8hd_decap_6
XFILLER_28_136 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_73 vpwr vgnd scs8hd_fill_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_6
XFILLER_19_114 vgnd vpwr scs8hd_decap_8
XFILLER_34_106 vgnd vpwr scs8hd_decap_4
XFILLER_35_92 vpwr vgnd scs8hd_fill_2
XFILLER_51_91 vpwr vgnd scs8hd_fill_2
XFILLER_51_80 vpwr vgnd scs8hd_fill_2
X_149_ address[1] _149_/B _161_/C _149_/X vgnd vpwr scs8hd_or3_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XPHY_123 vgnd vpwr scs8hd_decap_3
XPHY_112 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_decap_3
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_46_91 vgnd vpwr scs8hd_fill_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_131 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_1_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_102 vgnd vpwr scs8hd_decap_12
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_49 vpwr vgnd scs8hd_fill_2
XFILLER_53_15 vgnd vpwr scs8hd_decap_12
XFILLER_43_70 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_86 vgnd vpwr scs8hd_decap_6
XFILLER_4_64 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_48_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_108 vgnd vpwr scs8hd_decap_12
XFILLER_58_145 vgnd vpwr scs8hd_fill_1
X_182_ chany_top_in[6] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vgnd vpwr scs8hd_decap_12
XFILLER_49_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_137 vgnd vpwr scs8hd_decap_8
XFILLER_54_80 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_62_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_0.LATCH_5_.latch data_in mem_right_ipin_0.LATCH_5_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_55_126 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_29 vpwr vgnd scs8hd_fill_2
XFILLER_50_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_59_47 vpwr vgnd scs8hd_fill_2
XFILLER_24_83 vpwr vgnd scs8hd_fill_2
X_165_ _164_/X _132_/A vgnd vpwr scs8hd_buf_1
X_096_ _115_/A _094_/B _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_60 vpwr vgnd scs8hd_fill_2
XFILLER_37_126 vpwr vgnd scs8hd_fill_2
XFILLER_37_137 vpwr vgnd scs8hd_fill_2
XFILLER_20_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_17 vgnd vpwr scs8hd_decap_3
XFILLER_29_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XFILLER_61_59 vpwr vgnd scs8hd_fill_2
XFILLER_61_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_94 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
X_148_ address[0] _161_/C vgnd vpwr scs8hd_inv_8
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_079_ _134_/A _117_/A vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_5.LATCH_3_.latch/Q mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_118 vgnd vpwr scs8hd_decap_4
XFILLER_56_15 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_decap_3
XPHY_113 vgnd vpwr scs8hd_decap_3
XPHY_102 vgnd vpwr scs8hd_decap_3
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_30_143 vgnd vpwr scs8hd_decap_3
XFILLER_7_97 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_left_ipin_0.LATCH_4_.latch/Q mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_21_143 vgnd vpwr scs8hd_decap_3
XFILLER_8_114 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_53_27 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_1.LATCH_1_.latch data_in mem_right_ipin_1.LATCH_1_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_0_.latch/Q mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_93 vpwr vgnd scs8hd_fill_2
XFILLER_43_60 vgnd vpwr scs8hd_fill_1
XFILLER_4_54 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vpwr vgnd scs8hd_fill_2
XFILLER_48_27 vgnd vpwr scs8hd_decap_4
XFILLER_64_15 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_3.LATCH_4_.latch data_in mem_right_ipin_3.LATCH_4_.latch/Q _105_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_181_ chany_top_in[7] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_49_135 vgnd vpwr scs8hd_decap_8
XFILLER_49_102 vpwr vgnd scs8hd_fill_2
XANTENNA__100__B _100_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_19 vgnd vpwr scs8hd_fill_1
XFILLER_59_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_8 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_61_108 vgnd vpwr scs8hd_decap_12
X_095_ _073_/X _094_/B _095_/Y vgnd vpwr scs8hd_nor2_4
X_164_ _161_/A address[2] address[0] _164_/X vgnd vpwr scs8hd_or3_4
XFILLER_40_50 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XFILLER_52_119 vgnd vpwr scs8hd_decap_12
XFILLER_1_44 vpwr vgnd scs8hd_fill_2
XFILLER_1_66 vpwr vgnd scs8hd_fill_2
XANTENNA__111__A _110_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_1_.latch/Q mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_45_39 vpwr vgnd scs8hd_fill_2
XFILLER_45_28 vgnd vpwr scs8hd_decap_4
XFILLER_43_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_61_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_40 vpwr vgnd scs8hd_fill_2
XFILLER_19_73 vpwr vgnd scs8hd_fill_2
XFILLER_34_119 vpwr vgnd scs8hd_fill_2
X_078_ _116_/A _076_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _073_/X vgnd vpwr scs8hd_diode_2
X_147_ address[2] _149_/B vgnd vpwr scs8hd_inv_8
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_56_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_119 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_decap_3
XPHY_114 vgnd vpwr scs8hd_decap_3
XPHY_103 vgnd vpwr scs8hd_decap_3
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_5_.latch data_in mem_left_ipin_0.LATCH_5_.latch/Q _156_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_46_82 vgnd vpwr scs8hd_decap_6
XFILLER_46_71 vgnd vpwr scs8hd_decap_8
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_21 vpwr vgnd scs8hd_fill_2
XFILLER_8_126 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_4.LATCH_0_.latch data_in mem_right_ipin_4.LATCH_0_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_53_39 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_0_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_51 vgnd vpwr scs8hd_decap_4
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_27_95 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_6.LATCH_3_.latch data_in mem_right_ipin_6.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__114__A _073_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_64_27 vgnd vpwr scs8hd_decap_4
X_180_ chany_top_in[8] chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_86 vpwr vgnd scs8hd_fill_2
XFILLER_1_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_4.LATCH_3_.latch/Q mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_64_106 vgnd vpwr scs8hd_decap_12
XFILLER_38_72 vpwr vgnd scs8hd_fill_2
XFILLER_38_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_48_3 vgnd vpwr scs8hd_decap_12
XFILLER_55_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_59_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_163_ _166_/A _139_/A _163_/Y vgnd vpwr scs8hd_nor2_4
X_094_ _071_/X _094_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_73 vgnd vpwr scs8hd_decap_8
XFILLER_40_84 vpwr vgnd scs8hd_fill_2
XFILLER_49_60 vgnd vpwr scs8hd_fill_1
XFILLER_1_12 vpwr vgnd scs8hd_fill_2
XFILLER_1_89 vpwr vgnd scs8hd_fill_2
XFILLER_37_117 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_1.LATCH_1_.latch data_in _145_/A _143_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_106 vgnd vpwr scs8hd_decap_4
XFILLER_61_39 vgnd vpwr scs8hd_decap_12
XFILLER_10_21 vgnd vpwr scs8hd_fill_1
XFILLER_10_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_146_ _146_/A _146_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__106__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _073_/X vgnd vpwr scs8hd_diode_2
X_077_ _133_/A _116_/A vgnd vpwr scs8hd_buf_1
XFILLER_33_120 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_126 vgnd vpwr scs8hd_decap_3
XPHY_115 vgnd vpwr scs8hd_decap_3
XPHY_104 vgnd vpwr scs8hd_decap_3
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_53 vgnd vpwr scs8hd_decap_3
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_120 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_66 vgnd vpwr scs8hd_fill_1
XFILLER_7_11 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_129_ _129_/A _133_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_30_3 vgnd vpwr scs8hd_decap_6
XFILLER_21_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_138 vgnd vpwr scs8hd_decap_8
XFILLER_12_145 vgnd vpwr scs8hd_fill_1
XFILLER_32_41 vpwr vgnd scs8hd_fill_2
XFILLER_57_82 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_37_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_1_.latch/Q mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_30 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_74 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__114__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__130__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_78 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_58_104 vpwr vgnd scs8hd_fill_2
XFILLER_49_115 vgnd vpwr scs8hd_fill_1
XFILLER_8_3 vgnd vpwr scs8hd_decap_8
XFILLER_64_118 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__109__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _117_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_59_39 vgnd vpwr scs8hd_decap_8
X_162_ _162_/A _139_/A vgnd vpwr scs8hd_buf_1
X_093_ _156_/A _094_/B _093_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_41 vgnd vpwr scs8hd_decap_3
XFILLER_40_96 vpwr vgnd scs8hd_fill_2
XFILLER_49_83 vpwr vgnd scs8hd_fill_2
XFILLER_60_121 vgnd vpwr scs8hd_decap_8
XFILLER_60_110 vgnd vpwr scs8hd_decap_8
XFILLER_1_57 vgnd vpwr scs8hd_decap_4
XFILLER_60_3 vgnd vpwr scs8hd_decap_12
XFILLER_51_143 vgnd vpwr scs8hd_decap_3
XFILLER_19_53 vpwr vgnd scs8hd_fill_2
XFILLER_19_107 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_97 vgnd vpwr scs8hd_fill_1
XFILLER_35_30 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_51_62 vgnd vpwr scs8hd_decap_3
XFILLER_51_51 vgnd vpwr scs8hd_decap_8
X_145_ _145_/A _145_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_076_ _115_/A _076_/B _076_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_33_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_0_.latch/Q mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_decap_3
XPHY_105 vgnd vpwr scs8hd_decap_3
XFILLER_24_110 vgnd vpwr scs8hd_decap_4
XFILLER_24_143 vgnd vpwr scs8hd_decap_3
XPHY_127 vgnd vpwr scs8hd_decap_3
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_87 vpwr vgnd scs8hd_fill_2
XFILLER_62_72 vgnd vpwr scs8hd_decap_4
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_143 vgnd vpwr scs8hd_decap_3
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XANTENNA__133__A _133_/A vgnd vpwr scs8hd_diode_2
X_128_ _128_/A _133_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_34 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_8
XFILLER_21_135 vgnd vpwr scs8hd_decap_8
Xmux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _146_/Y mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_3.LATCH_3_.latch/Q mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_16_32 vpwr vgnd scs8hd_fill_2
XFILLER_32_64 vgnd vpwr scs8hd_decap_3
XANTENNA__128__A _128_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_43_74 vpwr vgnd scs8hd_fill_2
XFILLER_43_30 vpwr vgnd scs8hd_fill_2
XFILLER_4_131 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__130__B _133_/B vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ right_grid_pin_3_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_0_.latch data_in mem_right_ipin_0.LATCH_0_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_13_22 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_77 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_7.LATCH_4_.latch/Q mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_1_101 vgnd vpwr scs8hd_decap_4
XFILLER_1_112 vpwr vgnd scs8hd_fill_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XFILLER_54_84 vgnd vpwr scs8hd_decap_8
XFILLER_38_96 vpwr vgnd scs8hd_fill_2
XANTENNA__125__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA__141__A _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_3_.latch data_in mem_right_ipin_2.LATCH_3_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_141 vgnd vpwr scs8hd_decap_4
XFILLER_46_119 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB _064_/Y vgnd vpwr scs8hd_diode_2
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XFILLER_24_87 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_5.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_161_ _161_/A address[2] _161_/C _162_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
X_092_ _091_/X _094_/B vgnd vpwr scs8hd_buf_1
XFILLER_49_62 vgnd vpwr scs8hd_decap_4
XFILLER_1_25 vpwr vgnd scs8hd_fill_2
XFILLER_60_133 vgnd vpwr scs8hd_decap_12
XFILLER_45_141 vgnd vpwr scs8hd_decap_4
XFILLER_45_130 vpwr vgnd scs8hd_fill_2
XFILLER_53_3 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _135_/X vgnd vpwr scs8hd_diode_2
XFILLER_28_119 vgnd vpwr scs8hd_decap_8
XFILLER_10_67 vgnd vpwr scs8hd_decap_4
XFILLER_35_53 vpwr vgnd scs8hd_fill_2
XFILLER_35_75 vpwr vgnd scs8hd_fill_2
X_144_ _067_/X _101_/X address[0] _144_/Y vgnd vpwr scs8hd_nor3_4
X_075_ _132_/A _115_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_1_.latch/Q mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_128 vgnd vpwr scs8hd_decap_3
XPHY_117 vgnd vpwr scs8hd_decap_3
XPHY_106 vgnd vpwr scs8hd_decap_3
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_84 vgnd vpwr scs8hd_decap_8
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__133__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_127_ address[5] _127_/B _154_/C _128_/A vgnd vpwr scs8hd_or3_4
XFILLER_16_3 vgnd vpwr scs8hd_decap_8
XFILLER_21_114 vgnd vpwr scs8hd_decap_8
XFILLER_16_11 vgnd vpwr scs8hd_decap_3
XFILLER_16_55 vgnd vpwr scs8hd_fill_1
XFILLER_32_32 vpwr vgnd scs8hd_fill_2
XFILLER_32_76 vpwr vgnd scs8hd_fill_2
XFILLER_57_62 vgnd vpwr scs8hd_decap_4
XANTENNA__144__A _067_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_2_.latch/Q mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_43 vpwr vgnd scs8hd_fill_2
XFILLER_43_53 vgnd vpwr scs8hd_fill_1
XFILLER_4_143 vgnd vpwr scs8hd_decap_3
XFILLER_4_58 vgnd vpwr scs8hd_decap_6
XFILLER_4_36 vgnd vpwr scs8hd_decap_3
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_135 vgnd vpwr scs8hd_decap_8
Xmem_right_ipin_5.LATCH_2_.latch data_in mem_right_ipin_5.LATCH_2_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_54_63 vpwr vgnd scs8hd_fill_2
XFILLER_54_52 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_0_.latch/Q mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__141__B _140_/B vgnd vpwr scs8hd_diode_2
XFILLER_55_109 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_7.LATCH_5_.latch data_in mem_right_ipin_7.LATCH_5_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_66 vpwr vgnd scs8hd_fill_2
X_091_ _090_/Y address[6] _154_/C _091_/X vgnd vpwr scs8hd_or3_4
X_160_ address[1] _161_/A vgnd vpwr scs8hd_inv_8
XFILLER_45_120 vpwr vgnd scs8hd_fill_2
XFILLER_1_48 vgnd vpwr scs8hd_decap_3
XFILLER_37_109 vpwr vgnd scs8hd_fill_2
XFILLER_60_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_1_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__152__A enable vgnd vpwr scs8hd_diode_2
XFILLER_46_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_right_ipin_2.LATCH_3_.latch/Q mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_51_123 vgnd vpwr scs8hd_decap_12
XFILLER_51_112 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_24 vgnd vpwr scs8hd_decap_3
XANTENNA__062__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_19_22 vgnd vpwr scs8hd_decap_3
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_35_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_0_.latch data_in mem_left_ipin_0.LATCH_0_.latch/Q _064_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_074_ _073_/X _076_/B _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ _067_/X _101_/X _161_/C _143_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_5_.scs8hd_inv_1 chany_top_in[5] mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_33_112 vpwr vgnd scs8hd_fill_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A address[2] vgnd vpwr scs8hd_diode_2
XPHY_129 vgnd vpwr scs8hd_decap_3
XPHY_118 vgnd vpwr scs8hd_decap_3
XPHY_107 vgnd vpwr scs8hd_decap_3
XFILLER_24_123 vgnd vpwr scs8hd_decap_12
XFILLER_21_23 vpwr vgnd scs8hd_fill_2
XFILLER_21_78 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_112 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XFILLER_62_96 vgnd vpwr scs8hd_decap_3
X_126_ address[6] _127_/B vgnd vpwr scs8hd_inv_8
XFILLER_21_104 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_ipin_6.LATCH_4_.latch/Q mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_16_23 vgnd vpwr scs8hd_decap_3
XFILLER_16_45 vpwr vgnd scs8hd_fill_2
XFILLER_16_78 vpwr vgnd scs8hd_fill_2
XFILLER_32_88 vpwr vgnd scs8hd_fill_2
XFILLER_57_85 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _101_/X vgnd vpwr scs8hd_diode_2
X_109_ _117_/A _106_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_22 vgnd vpwr scs8hd_decap_6
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XFILLER_43_65 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_4
XANTENNA__139__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _171_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XANTENNA__065__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_49_118 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vpwr vgnd scs8hd_fill_2
XFILLER_38_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_1_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_143 vgnd vpwr scs8hd_decap_3
XFILLER_24_23 vgnd vpwr scs8hd_decap_8
X_090_ address[5] _090_/Y vgnd vpwr scs8hd_inv_8
XFILLER_49_53 vgnd vpwr scs8hd_decap_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_8
XFILLER_40_88 vgnd vpwr scs8hd_decap_4
XFILLER_39_3 vgnd vpwr scs8hd_decap_8
XFILLER_51_135 vgnd vpwr scs8hd_decap_8
XFILLER_10_36 vgnd vpwr scs8hd_decap_3
XANTENNA__062__B address[2] vgnd vpwr scs8hd_diode_2
X_142_ _134_/A _140_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_35_88 vpwr vgnd scs8hd_fill_2
XFILLER_51_87 vpwr vgnd scs8hd_fill_2
XFILLER_51_76 vpwr vgnd scs8hd_fill_2
X_073_ _139_/A _073_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_135 vgnd vpwr scs8hd_decap_8
XANTENNA__163__A _166_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_2_.latch/Q mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_119 vgnd vpwr scs8hd_decap_3
XPHY_108 vgnd vpwr scs8hd_decap_3
XFILLER_24_135 vgnd vpwr scs8hd_decap_8
XANTENNA__073__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_46_54 vpwr vgnd scs8hd_fill_2
XFILLER_46_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_135 vgnd vpwr scs8hd_decap_8
X_125_ _117_/A _120_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_90 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__158__A _157_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.INVTX1_5_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _065_/Y vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_0_.latch/Q mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_23 vgnd vpwr scs8hd_decap_8
XFILLER_32_45 vgnd vpwr scs8hd_decap_3
XFILLER_57_53 vpwr vgnd scs8hd_fill_2
XFILLER_57_42 vpwr vgnd scs8hd_fill_2
X_108_ _116_/A _106_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__144__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_80 vpwr vgnd scs8hd_fill_2
XANTENNA__070__B _076_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_1.LATCH_3_.latch/Q mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_58_108 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_54_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_63_111 vgnd vpwr scs8hd_decap_8
XANTENNA__166__A _166_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_70 vpwr vgnd scs8hd_fill_2
XANTENNA__076__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_23 vgnd vpwr scs8hd_decap_4
XFILLER_40_56 vpwr vgnd scs8hd_fill_2
XFILLER_49_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_1.LATCH_2_.latch data_in mem_right_ipin_1.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_90 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_5.LATCH_4_.latch/Q mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_6
XANTENNA__062__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_133 vpwr vgnd scs8hd_fill_2
X_141_ _133_/A _140_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_072_ _071_/X _076_/B _072_/Y vgnd vpwr scs8hd_nor2_4
Xmem_right_ipin_3.LATCH_5_.latch data_in mem_right_ipin_3.LATCH_5_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__163__B _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_51_3 vgnd vpwr scs8hd_decap_12
Xmux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _170_/HI mem_left_ipin_0.LATCH_5_.latch/Q
+ mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XFILLER_2_60 vgnd vpwr scs8hd_decap_4
XPHY_109 vgnd vpwr scs8hd_decap_3
XFILLER_21_36 vpwr vgnd scs8hd_fill_2
XFILLER_21_58 vgnd vpwr scs8hd_decap_3
XFILLER_62_32 vgnd vpwr scs8hd_decap_12
XFILLER_46_88 vgnd vpwr scs8hd_fill_1
XFILLER_30_106 vgnd vpwr scs8hd_decap_4
XFILLER_62_76 vgnd vpwr scs8hd_fill_1
XFILLER_7_38 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
X_124_ _116_/A _120_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_117 vgnd vpwr scs8hd_decap_12
XANTENNA__068__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__084__A _156_/A vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_1_.latch/Q mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_143 vgnd vpwr scs8hd_decap_3
XFILLER_7_121 vgnd vpwr scs8hd_fill_1
X_107_ _115_/A _106_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A _166_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_43_89 vpwr vgnd scs8hd_fill_2
XFILLER_43_56 vpwr vgnd scs8hd_fill_2
XFILLER_43_45 vpwr vgnd scs8hd_fill_2
XFILLER_27_79 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XFILLER_13_15 vgnd vpwr scs8hd_decap_4
XFILLER_13_26 vgnd vpwr scs8hd_fill_1
XFILLER_49_109 vgnd vpwr scs8hd_decap_6
XFILLER_1_116 vgnd vpwr scs8hd_decap_6
XFILLER_38_23 vgnd vpwr scs8hd_decap_4
XFILLER_54_44 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_2_.latch/Q mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_5.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_63_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__166__B _132_/A vgnd vpwr scs8hd_diode_2
XANTENNA__182__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_54_145 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_4.LATCH_1_.latch data_in mem_right_ipin_4.LATCH_1_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__076__B _076_/B vgnd vpwr scs8hd_diode_2
XFILLER_24_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _091_/X vgnd vpwr scs8hd_diode_2
XFILLER_40_46 vpwr vgnd scs8hd_fill_2
XFILLER_45_101 vpwr vgnd scs8hd_fill_2
XFILLER_1_29 vpwr vgnd scs8hd_fill_2
XFILLER_45_145 vgnd vpwr scs8hd_fill_1
XFILLER_45_112 vpwr vgnd scs8hd_fill_2
XFILLER_36_145 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_0_.latch/Q mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_ipin_6.LATCH_4_.latch data_in mem_right_ipin_6.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_36 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_112 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_decap_4
XFILLER_27_145 vgnd vpwr scs8hd_fill_1
XFILLER_35_57 vpwr vgnd scs8hd_fill_2
X_140_ _132_/A _140_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ _138_/A _071_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_145 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_44_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_15 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_0.LATCH_3_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_62_44 vgnd vpwr scs8hd_decap_12
XFILLER_7_17 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_123_ _115_/A _120_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__190__A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_129 vgnd vpwr scs8hd_decap_12
XFILLER_16_59 vgnd vpwr scs8hd_decap_8
XANTENNA__068__C _067_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_1_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__084__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_57_66 vgnd vpwr scs8hd_fill_1
X_106_ _073_/X _106_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__B _133_/A vgnd vpwr scs8hd_diode_2
XANTENNA__185__A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _146_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_60 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_47 vpwr vgnd scs8hd_fill_2
XANTENNA__095__A _073_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_29 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_4.LATCH_4_.latch/Q mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_57_132 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vpwr vgnd scs8hd_fill_2
XFILLER_38_79 vpwr vgnd scs8hd_fill_2
XFILLER_54_67 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_7.LATCH_0_.latch data_in mem_right_ipin_7.LATCH_0_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_63_135 vgnd vpwr scs8hd_decap_8
XFILLER_39_121 vgnd vpwr scs8hd_fill_1
XFILLER_54_113 vpwr vgnd scs8hd_fill_2
XFILLER_54_102 vpwr vgnd scs8hd_fill_2
XFILLER_24_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_4
XFILLER_30_91 vgnd vpwr scs8hd_fill_1
XFILLER_51_116 vgnd vpwr scs8hd_decap_6
XANTENNA__193__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_3.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_15 vgnd vpwr scs8hd_decap_4
XFILLER_42_138 vgnd vpwr scs8hd_decap_8
XFILLER_42_127 vpwr vgnd scs8hd_fill_2
XANTENNA__087__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_35_47 vgnd vpwr scs8hd_decap_4
X_070_ _156_/A _076_/B _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_102 vpwr vgnd scs8hd_fill_2
XFILLER_18_113 vgnd vpwr scs8hd_decap_12
XFILLER_33_105 vgnd vpwr scs8hd_decap_4
XFILLER_33_116 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_decap_3
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_2_84 vgnd vpwr scs8hd_decap_8
XANTENNA__188__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_116 vpwr vgnd scs8hd_fill_2
XFILLER_62_56 vgnd vpwr scs8hd_decap_12
XFILLER_30_119 vgnd vpwr scs8hd_decap_12
X_122_ _073_/X _120_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_108 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_49 vgnd vpwr scs8hd_decap_6
XFILLER_32_15 vgnd vpwr scs8hd_decap_4
XFILLER_32_37 vpwr vgnd scs8hd_fill_2
XFILLER_32_59 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_57_78 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_2_.latch/Q mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
X_105_ _071_/X _106_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_4
XANTENNA__095__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_0_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_57_144 vpwr vgnd scs8hd_fill_2
XFILLER_57_100 vpwr vgnd scs8hd_fill_2
XFILLER_38_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_91 vgnd vpwr scs8hd_fill_1
XFILLER_5_40 vpwr vgnd scs8hd_fill_2
XFILLER_39_111 vpwr vgnd scs8hd_fill_2
XFILLER_24_49 vgnd vpwr scs8hd_decap_6
XFILLER_40_15 vgnd vpwr scs8hd_decap_4
XFILLER_49_79 vpwr vgnd scs8hd_fill_2
XFILLER_49_57 vgnd vpwr scs8hd_fill_1
XFILLER_14_71 vpwr vgnd scs8hd_fill_2
XFILLER_39_90 vpwr vgnd scs8hd_fill_2
XFILLER_51_106 vgnd vpwr scs8hd_decap_4
XFILLER_36_125 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_1_.latch/Q mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_29 vpwr vgnd scs8hd_fill_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_1_.latch data_in mem_right_ipin_0.LATCH_1_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_125 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_decap_3
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_106 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_3.LATCH_4_.latch/Q mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_46_58 vpwr vgnd scs8hd_fill_2
XANTENNA__098__B _094_/B vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_4_.latch data_in mem_right_ipin_2.LATCH_4_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_62_79 vgnd vpwr scs8hd_fill_1
XFILLER_62_68 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_1.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_121_ _071_/X _120_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_28 vgnd vpwr scs8hd_decap_3
XFILLER_57_57 vpwr vgnd scs8hd_fill_2
XFILLER_57_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_135 vgnd vpwr scs8hd_decap_8
XFILLER_22_82 vpwr vgnd scs8hd_fill_2
X_104_ _156_/A _106_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_43_15 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_right_ipin_7.LATCH_5_.latch/Q
+ mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_left_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[1] mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_33_92 vgnd vpwr scs8hd_fill_1
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_29 vpwr vgnd scs8hd_fill_2
XFILLER_1_108 vpwr vgnd scs8hd_fill_2
XFILLER_57_112 vpwr vgnd scs8hd_fill_2
XFILLER_38_15 vgnd vpwr scs8hd_decap_4
XFILLER_48_145 vgnd vpwr scs8hd_fill_1
XFILLER_5_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_145 vgnd vpwr scs8hd_fill_1
XFILLER_39_123 vpwr vgnd scs8hd_fill_2
XFILLER_45_137 vpwr vgnd scs8hd_fill_2
XFILLER_45_126 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_3.LATCH_0_.latch data_in mem_right_ipin_3.LATCH_0_.latch/Q _109_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_137 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_2_.latch/Q mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_137 vgnd vpwr scs8hd_decap_8
XFILLER_35_27 vgnd vpwr scs8hd_fill_1
XFILLER_51_59 vpwr vgnd scs8hd_fill_2
XFILLER_51_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XFILLER_18_137 vgnd vpwr scs8hd_decap_8
XFILLER_25_71 vpwr vgnd scs8hd_fill_2
XPHY_60 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
X_197_ chany_bottom_in[0] chany_top_out[0] vgnd vpwr scs8hd_buf_2
XPHY_93 vgnd vpwr scs8hd_decap_3
XFILLER_41_92 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_5.LATCH_3_.latch data_in mem_right_ipin_5.LATCH_3_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_97 vgnd vpwr scs8hd_decap_8
XFILLER_2_64 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_15 vgnd vpwr scs8hd_decap_12
XFILLER_46_37 vpwr vgnd scs8hd_fill_2
X_120_ _129_/A _120_/B _120_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_0_.latch/Q mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_40 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_143 vgnd vpwr scs8hd_decap_3
XFILLER_22_50 vgnd vpwr scs8hd_decap_4
X_103_ _102_/X _106_/B vgnd vpwr scs8hd_buf_1
Xmem_left_ipin_0.LATCH_1_.latch data_in mem_left_ipin_0.LATCH_1_.latch/Q _169_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_43_49 vgnd vpwr scs8hd_decap_4
XFILLER_43_27 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_1_.latch/Q mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_71 vpwr vgnd scs8hd_fill_2
XFILLER_13_19 vgnd vpwr scs8hd_fill_1
XFILLER_54_15 vgnd vpwr scs8hd_decap_12
XFILLER_38_49 vgnd vpwr scs8hd_decap_6
XFILLER_48_113 vgnd vpwr scs8hd_decap_12
XFILLER_48_102 vgnd vpwr scs8hd_decap_8
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_2_.latch/Q mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_2.LATCH_4_.latch/Q mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.INVTX1_3_.scs8hd_inv_1 chany_top_in[7] mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_49_15 vgnd vpwr scs8hd_decap_12
XFILLER_45_116 vpwr vgnd scs8hd_fill_2
XFILLER_45_105 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__101__A _100_/X vgnd vpwr scs8hd_diode_2
XFILLER_42_108 vgnd vpwr scs8hd_decap_8
XFILLER_27_116 vgnd vpwr scs8hd_decap_6
XFILLER_51_27 vgnd vpwr scs8hd_decap_12
XPHY_94 vgnd vpwr scs8hd_decap_3
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
X_196_ chany_bottom_in[1] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_2_43 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _145_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _178_/HI mem_right_ipin_6.LATCH_5_.latch/Q
+ mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_46_27 vgnd vpwr scs8hd_decap_4
XFILLER_62_15 vgnd vpwr scs8hd_decap_12
XFILLER_15_108 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_93 vpwr vgnd scs8hd_fill_2
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_57_15 vgnd vpwr scs8hd_decap_12
X_102_ _099_/X _101_/X _102_/X vgnd vpwr scs8hd_or2_4
XFILLER_47_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_4_107 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vpwr vgnd scs8hd_fill_2
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_2_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__104__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_57_136 vgnd vpwr scs8hd_decap_8
XFILLER_54_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_48_125 vgnd vpwr scs8hd_decap_12
XFILLER_44_82 vgnd vpwr scs8hd_decap_4
XFILLER_44_71 vpwr vgnd scs8hd_fill_2
XFILLER_5_98 vpwr vgnd scs8hd_fill_2
XFILLER_5_87 vgnd vpwr scs8hd_decap_6
XFILLER_54_117 vgnd vpwr scs8hd_decap_12
XFILLER_54_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_0_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_19 vgnd vpwr scs8hd_fill_1
XFILLER_49_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_41 vpwr vgnd scs8hd_fill_2
XFILLER_14_96 vgnd vpwr scs8hd_decap_12
XFILLER_30_40 vpwr vgnd scs8hd_fill_2
XFILLER_30_84 vgnd vpwr scs8hd_fill_1
XFILLER_55_92 vpwr vgnd scs8hd_fill_2
XFILLER_19_19 vgnd vpwr scs8hd_fill_1
XFILLER_51_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_106 vgnd vpwr scs8hd_decap_4
XFILLER_33_109 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_4.INVTX1_3_.scs8hd_inv_1 chany_top_in[5] mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_95 vgnd vpwr scs8hd_decap_3
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
X_195_ chany_bottom_in[2] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA__112__A _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_27 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_1_.latch/Q mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_120 vgnd vpwr scs8hd_decap_12
XANTENNA__107__A _115_/A vgnd vpwr scs8hd_diode_2
X_178_ _178_/HI _178_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_3 vgnd vpwr scs8hd_decap_8
XFILLER_32_19 vgnd vpwr scs8hd_fill_1
Xmem_right_ipin_1.LATCH_3_.latch data_in mem_right_ipin_1.LATCH_3_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_145 vgnd vpwr scs8hd_fill_1
XFILLER_57_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_105 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_ipin_1.LATCH_4_.latch/Q mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
X_101_ _100_/X _101_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_22_63 vpwr vgnd scs8hd_fill_2
XFILLER_8_43 vpwr vgnd scs8hd_fill_2
XFILLER_8_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_27_19 vgnd vpwr scs8hd_fill_1
XFILLER_4_119 vgnd vpwr scs8hd_decap_12
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_95 vgnd vpwr scs8hd_fill_1
XANTENNA__104__B _106_/B vgnd vpwr scs8hd_diode_2
XFILLER_58_81 vgnd vpwr scs8hd_decap_8
XANTENNA__120__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_57_104 vpwr vgnd scs8hd_fill_2
XFILLER_38_29 vpwr vgnd scs8hd_fill_2
XFILLER_48_137 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_73 vpwr vgnd scs8hd_fill_2
XFILLER_28_84 vgnd vpwr scs8hd_decap_4
XFILLER_44_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_60_93 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _177_/HI mem_right_ipin_5.LATCH_5_.latch/Q
+ mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_115 vgnd vpwr scs8hd_decap_6
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_54_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_19 vgnd vpwr scs8hd_fill_1
XFILLER_49_39 vgnd vpwr scs8hd_decap_3
XFILLER_39_94 vpwr vgnd scs8hd_fill_2
XFILLER_58_3 vgnd vpwr scs8hd_decap_12
XFILLER_27_129 vpwr vgnd scs8hd_fill_2
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_25_30 vpwr vgnd scs8hd_fill_2
XPHY_96 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_132 vgnd vpwr scs8hd_decap_3
XFILLER_41_40 vgnd vpwr scs8hd_fill_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_decap_3
X_194_ chany_bottom_in[3] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_41_62 vgnd vpwr scs8hd_decap_3
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vgnd vpwr scs8hd_decap_4
XFILLER_2_12 vgnd vpwr scs8hd_decap_4
XANTENNA__112__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_143 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_2_.latch/Q mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_4.LATCH_2_.latch data_in mem_right_ipin_4.LATCH_2_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_132 vgnd vpwr scs8hd_decap_12
XFILLER_36_73 vpwr vgnd scs8hd_fill_2
XFILLER_36_84 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_177_ _177_/HI _177_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__107__B _106_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.INVTX1_3_.scs8hd_inv_1 chany_top_in[4] mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_117 vgnd vpwr scs8hd_decap_4
XFILLER_11_102 vgnd vpwr scs8hd_decap_12
XFILLER_11_135 vgnd vpwr scs8hd_decap_8
X_100_ address[4] _100_/B _100_/X vgnd vpwr scs8hd_or2_4
Xmem_right_ipin_6.LATCH_5_.latch data_in mem_right_ipin_6.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_86 vgnd vpwr scs8hd_decap_4
XFILLER_8_11 vgnd vpwr scs8hd_decap_3
XANTENNA__118__A _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_86 vpwr vgnd scs8hd_fill_2
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_71 vgnd vpwr scs8hd_fill_1
XANTENNA__120__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_57_116 vgnd vpwr scs8hd_decap_4
XFILLER_38_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_145 vgnd vpwr scs8hd_fill_1
XFILLER_63_119 vgnd vpwr scs8hd_decap_3
XFILLER_28_52 vpwr vgnd scs8hd_fill_2
XFILLER_60_72 vgnd vpwr scs8hd_decap_3
XFILLER_5_23 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_127 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_1_.latch/Q mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_54 vgnd vpwr scs8hd_decap_8
XFILLER_14_65 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _146_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_30_64 vgnd vpwr scs8hd_decap_3
XFILLER_36_108 vgnd vpwr scs8hd_decap_8
XFILLER_39_40 vpwr vgnd scs8hd_fill_2
XFILLER_39_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_130 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_right_ipin_0.LATCH_4_.latch/Q mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XPHY_64 vgnd vpwr scs8hd_decap_3
X_193_ chany_bottom_in[4] chany_top_out[4] vgnd vpwr scs8hd_buf_2
XPHY_97 vgnd vpwr scs8hd_decap_3
XPHY_86 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vpwr vgnd scs8hd_fill_2
XFILLER_25_75 vgnd vpwr scs8hd_decap_4
XPHY_75 vgnd vpwr scs8hd_decap_3
Xmem_right_ipin_7.LATCH_1_.latch data_in mem_right_ipin_7.LATCH_1_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_7.LATCH_2_.latch/Q mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_144 vpwr vgnd scs8hd_fill_2
XFILLER_52_84 vgnd vpwr scs8hd_decap_6
XFILLER_52_73 vpwr vgnd scs8hd_fill_2
X_176_ _176_/HI _176_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__123__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vgnd vpwr scs8hd_decap_8
XFILLER_22_32 vgnd vpwr scs8hd_decap_4
Xmux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _176_/HI mem_right_ipin_4.LATCH_5_.latch/Q
+ mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_73 vpwr vgnd scs8hd_fill_2
XFILLER_47_51 vgnd vpwr scs8hd_decap_3
XFILLER_8_56 vpwr vgnd scs8hd_fill_2
XFILLER_8_23 vgnd vpwr scs8hd_decap_8
XANTENNA__118__B _100_/B vgnd vpwr scs8hd_diode_2
XANTENNA__134__A _134_/A vgnd vpwr scs8hd_diode_2
X_159_ _166_/A _138_/A _159_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_12_ vgnd vpwr scs8hd_inv_1
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_3_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_31 vpwr vgnd scs8hd_fill_2
XFILLER_33_75 vpwr vgnd scs8hd_fill_2
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_143 vgnd vpwr scs8hd_decap_3
XFILLER_3_121 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_135 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_44_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_60_84 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _133_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XFILLER_39_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[4] mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_2_.latch/Q mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_32 vpwr vgnd scs8hd_fill_2
XFILLER_30_76 vpwr vgnd scs8hd_fill_2
XFILLER_30_87 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_7.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_73 vpwr vgnd scs8hd_fill_2
XANTENNA__142__A _134_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_142 vgnd vpwr scs8hd_decap_4
XFILLER_50_145 vgnd vpwr scs8hd_fill_1
XPHY_98 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_decap_3
XFILLER_41_145 vgnd vpwr scs8hd_fill_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_21 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_26_131 vgnd vpwr scs8hd_decap_4
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_76 vgnd vpwr scs8hd_decap_3
X_192_ chany_bottom_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_41_53 vpwr vgnd scs8hd_fill_2
XFILLER_41_20 vgnd vpwr scs8hd_decap_4
XFILLER_2_47 vpwr vgnd scs8hd_fill_2
XANTENNA__137__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_145 vgnd vpwr scs8hd_fill_1
XFILLER_63_3 vgnd vpwr scs8hd_decap_12
XFILLER_23_101 vpwr vgnd scs8hd_fill_2
XFILLER_23_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_23 vpwr vgnd scs8hd_fill_2
XFILLER_11_78 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_175_ _175_/HI _175_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_104 vgnd vpwr scs8hd_decap_8
XFILLER_20_115 vgnd vpwr scs8hd_decap_12
XFILLER_22_11 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_63_51 vgnd vpwr scs8hd_decap_8
XFILLER_47_85 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_1_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_63_95 vpwr vgnd scs8hd_fill_2
XFILLER_63_62 vgnd vpwr scs8hd_decap_12
XFILLER_8_68 vgnd vpwr scs8hd_fill_1
XANTENNA__118__C _099_/X vgnd vpwr scs8hd_diode_2
XANTENNA__134__B _133_/B vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_2_.latch data_in mem_right_ipin_0.LATCH_2_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_089_ _117_/A _083_/X _089_/Y vgnd vpwr scs8hd_nor2_4
X_158_ _157_/X _138_/A vgnd vpwr scs8hd_buf_1
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A _149_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_22 vpwr vgnd scs8hd_fill_2
XFILLER_17_66 vgnd vpwr scs8hd_decap_3
XFILLER_17_99 vpwr vgnd scs8hd_fill_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_54 vgnd vpwr scs8hd_fill_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__129__B _133_/B vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_5_.latch data_in mem_right_ipin_2.LATCH_5_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_6
XFILLER_39_107 vpwr vgnd scs8hd_fill_2
XFILLER_5_36 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_6.LATCH_2_.latch/Q mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_53_143 vgnd vpwr scs8hd_decap_3
XFILLER_38_140 vgnd vpwr scs8hd_decap_6
XFILLER_14_23 vgnd vpwr scs8hd_decap_8
XFILLER_30_44 vpwr vgnd scs8hd_fill_2
XFILLER_55_52 vgnd vpwr scs8hd_decap_3
XFILLER_39_53 vpwr vgnd scs8hd_fill_2
XFILLER_55_96 vpwr vgnd scs8hd_fill_2
XANTENNA__142__B _140_/B vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _175_/HI mem_right_ipin_3.LATCH_5_.latch/Q
+ mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_6_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_99 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_decap_3
XFILLER_41_113 vgnd vpwr scs8hd_decap_3
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_25_55 vgnd vpwr scs8hd_decap_4
XFILLER_25_99 vgnd vpwr scs8hd_decap_4
XPHY_55 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_77 vgnd vpwr scs8hd_decap_3
X_191_ chany_bottom_in[6] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_41_98 vpwr vgnd scs8hd_fill_2
XFILLER_41_43 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_110 vpwr vgnd scs8hd_fill_2
XFILLER_17_143 vgnd vpwr scs8hd_decap_3
XANTENNA__137__B _140_/B vgnd vpwr scs8hd_diode_2
XFILLER_56_3 vgnd vpwr scs8hd_decap_12
XANTENNA__153__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_5.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _062_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vpwr vgnd scs8hd_fill_2
XFILLER_36_65 vpwr vgnd scs8hd_fill_2
X_174_ _174_/HI _174_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__148__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_127 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _170_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_right_ipin_3.LATCH_1_.latch data_in mem_right_ipin_3.LATCH_1_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_78 vpwr vgnd scs8hd_fill_2
XFILLER_63_74 vgnd vpwr scs8hd_decap_12
XFILLER_6_120 vgnd vpwr scs8hd_decap_12
X_157_ address[1] _149_/B address[0] _157_/X vgnd vpwr scs8hd_or3_4
X_088_ _116_/A _083_/X _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_left_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_5.LATCH_4_.latch data_in mem_right_ipin_5.LATCH_4_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_56 vpwr vgnd scs8hd_fill_2
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_88 vgnd vpwr scs8hd_decap_4
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_104 vpwr vgnd scs8hd_fill_2
XANTENNA__071__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_11 vgnd vpwr scs8hd_decap_3
XFILLER_28_88 vgnd vpwr scs8hd_fill_1
XFILLER_44_32 vgnd vpwr scs8hd_decap_3
XFILLER_5_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA__066__A address[5] vgnd vpwr scs8hd_diode_2
Xmem_left_ipin_0.LATCH_2_.latch data_in mem_left_ipin_0.LATCH_2_.latch/Q _166_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_30_12 vgnd vpwr scs8hd_decap_4
XFILLER_30_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_44_144 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_130 vgnd vpwr scs8hd_decap_12
XFILLER_50_125 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_1_.latch/Q mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_190_ chany_bottom_in[7] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XPHY_89 vgnd vpwr scs8hd_decap_3
XFILLER_41_11 vgnd vpwr scs8hd_decap_3
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_25_23 vpwr vgnd scs8hd_fill_2
XFILLER_25_34 vpwr vgnd scs8hd_fill_2
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_78 vgnd vpwr scs8hd_decap_3
XANTENNA__153__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_49_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_36 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_52_32 vgnd vpwr scs8hd_decap_12
X_173_ _173_/HI _173_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_6.LATCH_0_.latch data_in mem_right_ipin_6.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_139 vgnd vpwr scs8hd_decap_6
XANTENNA__164__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _073_/X vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[5] mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_46 vpwr vgnd scs8hd_fill_2
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_47_98 vpwr vgnd scs8hd_fill_2
XFILLER_63_86 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_5.LATCH_2_.latch/Q mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_37 vgnd vpwr scs8hd_decap_4
XFILLER_6_132 vgnd vpwr scs8hd_decap_12
X_087_ _115_/A _083_/X _087_/Y vgnd vpwr scs8hd_nor2_4
X_156_ _156_/A _166_/A _156_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__159__A _166_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _145_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_23 vgnd vpwr scs8hd_decap_3
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_64 vgnd vpwr scs8hd_decap_4
XFILLER_3_135 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _174_/HI mem_right_ipin_2.LATCH_5_.latch/Q
+ mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_139_ _139_/A _140_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_28_23 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vpwr vgnd scs8hd_fill_2
XFILLER_44_88 vpwr vgnd scs8hd_fill_2
XFILLER_60_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_62_145 vgnd vpwr scs8hd_fill_1
XFILLER_62_101 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _166_/A vgnd vpwr scs8hd_diode_2
XFILLER_53_123 vgnd vpwr scs8hd_decap_12
XFILLER_53_112 vpwr vgnd scs8hd_fill_2
XANTENNA__066__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_11 vgnd vpwr scs8hd_decap_3
XFILLER_39_77 vpwr vgnd scs8hd_fill_2
XFILLER_29_142 vgnd vpwr scs8hd_decap_4
XFILLER_50_137 vgnd vpwr scs8hd_decap_8
XANTENNA__167__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _133_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_137 vgnd vpwr scs8hd_decap_8
XPHY_79 vgnd vpwr scs8hd_decap_3
XFILLER_25_79 vgnd vpwr scs8hd_fill_1
XPHY_57 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XFILLER_41_78 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_32_104 vgnd vpwr scs8hd_decap_8
XFILLER_32_115 vgnd vpwr scs8hd_decap_12
XANTENNA__153__C _066_/C vgnd vpwr scs8hd_diode_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_44 vgnd vpwr scs8hd_decap_12
X_172_ _172_/HI _172_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__164__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_61_3 vgnd vpwr scs8hd_decap_12
XANTENNA__180__A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_93 vpwr vgnd scs8hd_fill_2
XANTENNA__074__B _076_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_36 vgnd vpwr scs8hd_fill_1
XANTENNA__090__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_47_77 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_0.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_144 vpwr vgnd scs8hd_fill_2
X_086_ _073_/X _083_/X _086_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
X_155_ _155_/A _166_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__159__B _138_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__A _071_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_35 vpwr vgnd scs8hd_fill_2
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_32 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
X_138_ _138_/A _140_/B _138_/Y vgnd vpwr scs8hd_nor2_4
X_069_ _068_/X _076_/B vgnd vpwr scs8hd_buf_1
XANTENNA__161__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_ipin_0.LATCH_1_.latch/Q mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_50 vpwr vgnd scs8hd_fill_2
XFILLER_0_72 vgnd vpwr scs8hd_decap_3
XFILLER_0_94 vgnd vpwr scs8hd_decap_6
XFILLER_0_139 vgnd vpwr scs8hd_decap_6
XFILLER_56_132 vgnd vpwr scs8hd_decap_12
XFILLER_56_121 vpwr vgnd scs8hd_fill_2
XFILLER_28_35 vpwr vgnd scs8hd_fill_2
XFILLER_60_55 vgnd vpwr scs8hd_decap_8
XFILLER_60_44 vgnd vpwr scs8hd_decap_8
XFILLER_44_67 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.LATCH_4_.latch data_in mem_right_ipin_1.LATCH_4_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_60_88 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_47_143 vgnd vpwr scs8hd_decap_3
XFILLER_47_121 vgnd vpwr scs8hd_fill_1
XFILLER_62_113 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_7.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_53_135 vgnd vpwr scs8hd_decap_8
XFILLER_14_15 vgnd vpwr scs8hd_decap_4
XFILLER_14_37 vpwr vgnd scs8hd_fill_2
XANTENNA__066__C _066_/C vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _100_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_36 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_121 vgnd vpwr scs8hd_fill_1
XFILLER_39_23 vpwr vgnd scs8hd_fill_2
XFILLER_55_77 vpwr vgnd scs8hd_fill_2
XFILLER_44_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_113 vgnd vpwr scs8hd_decap_3
XANTENNA__183__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__167__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_4.LATCH_2_.latch/Q mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_26_102 vpwr vgnd scs8hd_fill_2
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_decap_3
XFILLER_41_57 vpwr vgnd scs8hd_fill_2
XFILLER_41_24 vgnd vpwr scs8hd_fill_1
XANTENNA__093__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_29 vpwr vgnd scs8hd_fill_2
XFILLER_2_18 vpwr vgnd scs8hd_fill_2
XFILLER_17_135 vgnd vpwr scs8hd_decap_8
XFILLER_15_80 vpwr vgnd scs8hd_fill_2
XFILLER_32_127 vgnd vpwr scs8hd_decap_12
XFILLER_31_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__088__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_52_56 vgnd vpwr scs8hd_decap_6
Xmux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _173_/HI mem_right_ipin_1.LATCH_5_.latch/Q
+ mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_52_67 vgnd vpwr scs8hd_decap_4
X_171_ _171_/HI _171_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__164__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_54_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_22_59 vpwr vgnd scs8hd_fill_2
XFILLER_47_56 vgnd vpwr scs8hd_decap_3
XFILLER_47_34 vpwr vgnd scs8hd_fill_2
XFILLER_63_99 vgnd vpwr scs8hd_decap_12
X_085_ _071_/X _083_/X _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ address[5] address[6] _154_/C _155_/A vgnd vpwr scs8hd_or3_4
XANTENNA__191__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_2.LATCH_0_.latch data_in mem_right_ipin_2.LATCH_0_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_4
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _083_/X vgnd vpwr scs8hd_diode_2
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_137_ _129_/A _140_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_068_ _065_/Y address[3] _067_/X _068_/X vgnd vpwr scs8hd_or3_4
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
Xmem_right_ipin_4.LATCH_3_.latch data_in mem_right_ipin_4.LATCH_3_.latch/Q _114_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_60 vgnd vpwr scs8hd_fill_1
XANTENNA__186__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_84 vpwr vgnd scs8hd_fill_2
XFILLER_9_82 vpwr vgnd scs8hd_fill_2
XFILLER_56_144 vpwr vgnd scs8hd_fill_2
XFILLER_44_46 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_69 vpwr vgnd scs8hd_fill_2
XFILLER_60_67 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_62_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_100 vgnd vpwr scs8hd_decap_8
XANTENNA__082__C _067_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_59 vgnd vpwr scs8hd_decap_3
XFILLER_39_57 vpwr vgnd scs8hd_fill_2
XFILLER_44_136 vgnd vpwr scs8hd_decap_8
XFILLER_44_125 vpwr vgnd scs8hd_fill_2
XANTENNA__167__C _161_/C vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_8
XPHY_59 vgnd vpwr scs8hd_decap_3
Xmux_right_ipin_5.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_36 vgnd vpwr scs8hd_decap_4
XANTENNA__093__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_103 vpwr vgnd scs8hd_fill_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_32_139 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_6.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__088__B _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_36 vgnd vpwr scs8hd_fill_1
XFILLER_36_69 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_170_ _170_/HI _170_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_143 vgnd vpwr scs8hd_decap_3
XFILLER_9_110 vpwr vgnd scs8hd_fill_2
XFILLER_47_3 vgnd vpwr scs8hd_decap_12
XANTENNA__189__A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_3
XFILLER_22_16 vgnd vpwr scs8hd_decap_12
XANTENNA__099__A _090_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _172_/HI vgnd vpwr
+ scs8hd_diode_2
X_153_ address[4] address[3] _066_/C _154_/C vgnd vpwr scs8hd_or3_4
X_084_ _156_/A _083_/X _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_93 vgnd vpwr scs8hd_decap_12
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_15 vgnd vpwr scs8hd_decap_8
XFILLER_33_48 vgnd vpwr scs8hd_decap_6
Xmem_right_ipin_7.LATCH_2_.latch data_in mem_right_ipin_7.LATCH_2_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_105 vpwr vgnd scs8hd_fill_2
XFILLER_59_131 vpwr vgnd scs8hd_fill_2
XFILLER_59_120 vpwr vgnd scs8hd_fill_2
XFILLER_58_89 vgnd vpwr scs8hd_decap_3
X_136_ _135_/X _140_/B vgnd vpwr scs8hd_buf_1
XFILLER_23_92 vgnd vpwr scs8hd_decap_3
X_067_ _066_/X _067_/X vgnd vpwr scs8hd_buf_1
Xmux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_3.LATCH_2_.latch/Q mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_50 vgnd vpwr scs8hd_decap_8
XFILLER_0_108 vgnd vpwr scs8hd_decap_4
XANTENNA__096__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_62_137 vgnd vpwr scs8hd_decap_8
XFILLER_47_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_119_ _119_/A _120_/B vgnd vpwr scs8hd_buf_1
XANTENNA__197__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _172_/HI mem_right_ipin_0.LATCH_5_.latch/Q
+ mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_16 vgnd vpwr scs8hd_fill_1
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XFILLER_39_36 vpwr vgnd scs8hd_fill_2
XFILLER_55_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_45_90 vpwr vgnd scs8hd_fill_2
XFILLER_35_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_118 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_25_49 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_40_140 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_48 vgnd vpwr scs8hd_decap_8
XFILLER_7_3 vgnd vpwr scs8hd_decap_8
Xmux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_3.INVTX1_1_.scs8hd_inv_1 chany_top_in[0] mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_91 vgnd vpwr scs8hd_fill_1
XFILLER_3_41 vgnd vpwr scs8hd_decap_3
XFILLER_22_28 vgnd vpwr scs8hd_decap_3
XANTENNA__099__B address[6] vgnd vpwr scs8hd_diode_2
X_083_ _082_/X _083_/X vgnd vpwr scs8hd_buf_1
XFILLER_12_72 vgnd vpwr scs8hd_decap_4
X_152_ enable _066_/C vgnd vpwr scs8hd_inv_8
Xmux_right_ipin_4.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_39 vpwr vgnd scs8hd_fill_2
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_59_143 vgnd vpwr scs8hd_decap_3
XFILLER_58_68 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_71 vpwr vgnd scs8hd_fill_2
X_135_ address[5] _127_/B _066_/C _101_/X _135_/X vgnd vpwr scs8hd_or4_4
X_066_ address[5] address[6] _066_/C _066_/X vgnd vpwr scs8hd_or3_4
XFILLER_9_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_16 vgnd vpwr scs8hd_decap_4
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XFILLER_44_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XFILLER_47_113 vpwr vgnd scs8hd_fill_2
XFILLER_47_102 vgnd vpwr scs8hd_decap_4
XFILLER_47_135 vgnd vpwr scs8hd_decap_8
X_118_ _065_/Y _100_/B _099_/X _119_/A vgnd vpwr scs8hd_or3_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_8
XFILLER_53_116 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_0.LATCH_3_.latch data_in mem_right_ipin_0.LATCH_3_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_102 vpwr vgnd scs8hd_fill_2
XFILLER_55_47 vgnd vpwr scs8hd_decap_3
XFILLER_29_113 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_81 vpwr vgnd scs8hd_fill_2
XFILLER_50_108 vgnd vpwr scs8hd_decap_8
XFILLER_35_105 vpwr vgnd scs8hd_fill_2
XFILLER_61_90 vgnd vpwr scs8hd_decap_3
XFILLER_6_41 vgnd vpwr scs8hd_decap_4
XFILLER_6_96 vgnd vpwr scs8hd_decap_12
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_26_138 vgnd vpwr scs8hd_decap_8
XFILLER_41_16 vpwr vgnd scs8hd_fill_2
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_52_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_108 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_2.LATCH_2_.latch/Q mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
Xmux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_ipin_0.LATCH_0_.latch/Q mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_47_15 vgnd vpwr scs8hd_decap_12
XANTENNA__099__C _066_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_51 vpwr vgnd scs8hd_fill_2
X_082_ _065_/Y _100_/B _067_/X _082_/X vgnd vpwr scs8hd_or3_4
X_151_ _129_/A _156_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _173_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_92 vpwr vgnd scs8hd_fill_2
XFILLER_53_91 vpwr vgnd scs8hd_fill_2
XFILLER_52_3 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[2] mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_58_47 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_134_ _134_/A _133_/B _134_/Y vgnd vpwr scs8hd_nor2_4
X_065_ address[4] _065_/Y vgnd vpwr scs8hd_inv_8
XFILLER_0_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_2.INVTX1_5_.scs8hd_inv_1 chany_top_in[8] mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_56_125 vgnd vpwr scs8hd_decap_4
XFILLER_28_39 vpwr vgnd scs8hd_fill_2
XFILLER_60_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_27 vgnd vpwr scs8hd_decap_4
Xmem_right_ipin_3.LATCH_2_.latch data_in mem_right_ipin_3.LATCH_2_.latch/Q _107_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_50 vpwr vgnd scs8hd_fill_2
X_117_ _117_/A _115_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_8
XFILLER_14_19 vgnd vpwr scs8hd_fill_1
XFILLER_55_15 vgnd vpwr scs8hd_decap_12
XFILLER_44_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_right_ipin_5.LATCH_5_.latch data_in mem_right_ipin_5.LATCH_5_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_73 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_75 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_26_106 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_4
XFILLER_15_62 vgnd vpwr scs8hd_decap_4
XFILLER_15_84 vpwr vgnd scs8hd_fill_2
XFILLER_31_50 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A _099_/X vgnd vpwr scs8hd_diode_2
XFILLER_56_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_52_27 vgnd vpwr scs8hd_decap_4
Xmem_left_ipin_0.LATCH_3_.latch data_in mem_left_ipin_0.LATCH_3_.latch/Q _163_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_135 vgnd vpwr scs8hd_decap_8
XFILLER_42_93 vpwr vgnd scs8hd_fill_2
XFILLER_3_76 vgnd vpwr scs8hd_decap_6
XFILLER_63_15 vgnd vpwr scs8hd_decap_12
XFILLER_47_38 vpwr vgnd scs8hd_fill_2
XFILLER_47_27 vgnd vpwr scs8hd_decap_4
XFILLER_63_59 vpwr vgnd scs8hd_fill_2
X_150_ _149_/X _129_/A vgnd vpwr scs8hd_buf_1
X_081_ address[3] _100_/B vgnd vpwr scs8hd_inv_8
XFILLER_37_71 vgnd vpwr scs8hd_decap_4
XFILLER_45_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_59_112 vgnd vpwr scs8hd_decap_6
XFILLER_58_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_133_ _133_/A _133_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_064_ _166_/A _134_/A _064_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__110__A _065_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_31 vpwr vgnd scs8hd_fill_2
XFILLER_0_77 vgnd vpwr scs8hd_decap_3
XFILLER_0_88 vgnd vpwr scs8hd_decap_4
XFILLER_9_86 vpwr vgnd scs8hd_fill_2
XFILLER_56_104 vgnd vpwr scs8hd_decap_6
Xmem_right_ipin_6.LATCH_1_.latch data_in mem_right_ipin_6.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_60_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_18_73 vpwr vgnd scs8hd_fill_2
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
XFILLER_34_72 vgnd vpwr scs8hd_decap_4
XFILLER_50_93 vpwr vgnd scs8hd_fill_2
XFILLER_50_71 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _071_/X vgnd vpwr scs8hd_diode_2
XFILLER_34_83 vgnd vpwr scs8hd_decap_6
X_116_ _116_/A _115_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_59_91 vpwr vgnd scs8hd_fill_2
XFILLER_30_19 vgnd vpwr scs8hd_fill_1
Xmux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_ipin_1.LATCH_2_.latch/Q mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_126 vpwr vgnd scs8hd_fill_2
XFILLER_55_27 vgnd vpwr scs8hd_decap_12
Xmux_right_ipin_0.INVTX1_5_.scs8hd_inv_1 chany_top_in[6] mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_118 vpwr vgnd scs8hd_fill_2
XFILLER_61_70 vpwr vgnd scs8hd_fill_2
XFILLER_45_82 vpwr vgnd scs8hd_fill_2
XFILLER_45_71 vpwr vgnd scs8hd_fill_2
XFILLER_6_87 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vgnd vpwr scs8hd_decap_4
XFILLER_40_121 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__102__B _101_/X vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_121 vgnd vpwr scs8hd_fill_1
XFILLER_31_143 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_ipin_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[8] mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_42_83 vpwr vgnd scs8hd_fill_2
XFILLER_42_72 vpwr vgnd scs8hd_fill_2
XFILLER_9_114 vgnd vpwr scs8hd_decap_8
XFILLER_9_103 vgnd vpwr scs8hd_decap_4
XFILLER_13_143 vgnd vpwr scs8hd_decap_3
XANTENNA__113__A _071_/X vgnd vpwr scs8hd_diode_2
XFILLER_63_27 vgnd vpwr scs8hd_decap_12
X_080_ _117_/A _076_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_102 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _174_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_53_71 vpwr vgnd scs8hd_fill_2
XANTENNA__108__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_109 vgnd vpwr scs8hd_decap_12
XFILLER_59_135 vgnd vpwr scs8hd_decap_8
XFILLER_58_27 vgnd vpwr scs8hd_decap_4
X_132_ _132_/A _133_/B _132_/Y vgnd vpwr scs8hd_nor2_4
X_063_ _062_/X _134_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_120 vgnd vpwr scs8hd_decap_12
XFILLER_48_82 vpwr vgnd scs8hd_fill_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__105__B _106_/B vgnd vpwr scs8hd_diode_2
X_115_ _115_/A _115_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__A _071_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_55_39 vgnd vpwr scs8hd_decap_8
XFILLER_44_119 vgnd vpwr scs8hd_decap_4
XFILLER_29_51 vpwr vgnd scs8hd_fill_2
XFILLER_29_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_11 vgnd vpwr scs8hd_decap_3
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_26_119 vgnd vpwr scs8hd_decap_12
XFILLER_40_100 vpwr vgnd scs8hd_fill_2
XFILLER_15_20 vgnd vpwr scs8hd_decap_4
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XFILLER_31_30 vpwr vgnd scs8hd_fill_2
Xmem_right_ipin_1.LATCH_5_.latch data_in mem_right_ipin_1.LATCH_5_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_111 vpwr vgnd scs8hd_fill_2
Xmux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ left_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

