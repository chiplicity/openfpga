magic
tech sky130A
magscale 1 2
timestamp 1606475702
<< locali >>
rect 12449 17595 12483 17833
rect 4721 17187 4755 17289
rect 10241 17051 10275 17221
rect 3801 15351 3835 15521
rect 3893 15487 3927 15657
rect 5917 15487 5951 15657
rect 3985 13719 4019 13889
rect 7205 13243 7239 13345
rect 11437 13175 11471 13277
rect 3617 12631 3651 12733
rect 12817 12699 12851 12801
rect 15393 12631 15427 12733
rect 10793 11543 10827 11713
rect 2145 10115 2179 10217
rect 4905 9979 4939 10217
rect 4997 9911 5031 10149
rect 14289 9503 14323 9605
rect 10517 9367 10551 9469
rect 9229 8823 9263 9129
rect 12265 8347 12299 8517
rect 7205 7871 7239 8041
rect 7389 6647 7423 6817
rect 16773 5627 16807 5797
rect 14289 5151 14323 5321
rect 10793 3995 10827 4165
rect 13369 2907 13403 3145
<< viali >>
rect 4445 20009 4479 20043
rect 4537 20009 4571 20043
rect 10701 20009 10735 20043
rect 12817 20009 12851 20043
rect 13369 20009 13403 20043
rect 14381 20009 14415 20043
rect 14933 20009 14967 20043
rect 15669 20009 15703 20043
rect 16221 20009 16255 20043
rect 17325 20009 17359 20043
rect 3341 19941 3375 19975
rect 9137 19941 9171 19975
rect 11529 19941 11563 19975
rect 1685 19873 1719 19907
rect 2237 19873 2271 19907
rect 3065 19873 3099 19907
rect 5448 19873 5482 19907
rect 7113 19873 7147 19907
rect 8217 19873 8251 19907
rect 8861 19873 8895 19907
rect 10609 19873 10643 19907
rect 11253 19873 11287 19907
rect 11989 19873 12023 19907
rect 12639 19873 12673 19907
rect 13185 19873 13219 19907
rect 14197 19873 14231 19907
rect 14749 19873 14783 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 17141 19873 17175 19907
rect 2421 19805 2455 19839
rect 4721 19805 4755 19839
rect 5181 19805 5215 19839
rect 7297 19805 7331 19839
rect 8309 19805 8343 19839
rect 8401 19805 8435 19839
rect 9781 19805 9815 19839
rect 10885 19805 10919 19839
rect 7849 19737 7883 19771
rect 12173 19737 12207 19771
rect 1869 19669 1903 19703
rect 4077 19669 4111 19703
rect 6561 19669 6595 19703
rect 10241 19669 10275 19703
rect 7021 19465 7055 19499
rect 11989 19329 12023 19363
rect 1593 19261 1627 19295
rect 2145 19261 2179 19295
rect 2973 19261 3007 19295
rect 3240 19261 3274 19295
rect 5089 19261 5123 19295
rect 6837 19261 6871 19295
rect 7389 19261 7423 19295
rect 9045 19261 9079 19295
rect 9505 19261 9539 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 14933 19261 14967 19295
rect 16037 19261 16071 19295
rect 16589 19261 16623 19295
rect 17141 19261 17175 19295
rect 18061 19261 18095 19295
rect 18613 19261 18647 19295
rect 19349 19261 19383 19295
rect 2421 19193 2455 19227
rect 4629 19193 4663 19227
rect 5356 19193 5390 19227
rect 7656 19193 7690 19227
rect 9772 19193 9806 19227
rect 12716 19193 12750 19227
rect 15577 19193 15611 19227
rect 1777 19125 1811 19159
rect 4353 19125 4387 19159
rect 6469 19125 6503 19159
rect 8769 19125 8803 19159
rect 10885 19125 10919 19159
rect 11345 19125 11379 19159
rect 11713 19125 11747 19159
rect 11805 19125 11839 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 16221 19125 16255 19159
rect 16773 19125 16807 19159
rect 17325 19125 17359 19159
rect 18245 19125 18279 19159
rect 18797 19125 18831 19159
rect 19533 19125 19567 19159
rect 2973 18921 3007 18955
rect 3341 18921 3375 18955
rect 3433 18921 3467 18955
rect 6561 18921 6595 18955
rect 8677 18921 8711 18955
rect 8953 18921 8987 18955
rect 13277 18921 13311 18955
rect 4445 18853 4479 18887
rect 6837 18853 6871 18887
rect 7564 18853 7598 18887
rect 9956 18853 9990 18887
rect 13829 18853 13863 18887
rect 14565 18853 14599 18887
rect 15577 18853 15611 18887
rect 18705 18853 18739 18887
rect 1409 18785 1443 18819
rect 2329 18785 2363 18819
rect 5181 18785 5215 18819
rect 5448 18785 5482 18819
rect 11345 18785 11379 18819
rect 11897 18785 11931 18819
rect 12164 18785 12198 18819
rect 13553 18785 13587 18819
rect 14289 18785 14323 18819
rect 15301 18785 15335 18819
rect 18429 18785 18463 18819
rect 2421 18717 2455 18751
rect 2605 18717 2639 18751
rect 3617 18717 3651 18751
rect 4537 18717 4571 18751
rect 4629 18717 4663 18751
rect 7297 18717 7331 18751
rect 9689 18717 9723 18751
rect 1593 18649 1627 18683
rect 4077 18649 4111 18683
rect 1961 18581 1995 18615
rect 11069 18581 11103 18615
rect 11529 18581 11563 18615
rect 4905 18377 4939 18411
rect 6837 18377 6871 18411
rect 8217 18377 8251 18411
rect 10885 18377 10919 18411
rect 14657 18377 14691 18411
rect 1685 18309 1719 18343
rect 5181 18309 5215 18343
rect 6377 18309 6411 18343
rect 9229 18309 9263 18343
rect 13461 18309 13495 18343
rect 2237 18241 2271 18275
rect 3525 18241 3559 18275
rect 5733 18241 5767 18275
rect 7297 18241 7331 18275
rect 7389 18241 7423 18275
rect 8861 18241 8895 18275
rect 9781 18241 9815 18275
rect 11529 18241 11563 18275
rect 13001 18241 13035 18275
rect 14013 18241 14047 18275
rect 1501 18173 1535 18207
rect 2053 18173 2087 18207
rect 2789 18173 2823 18207
rect 3792 18173 3826 18207
rect 5641 18173 5675 18207
rect 6193 18173 6227 18207
rect 8585 18173 8619 18207
rect 9689 18173 9723 18207
rect 11897 18173 11931 18207
rect 12817 18173 12851 18207
rect 14473 18173 14507 18207
rect 3065 18105 3099 18139
rect 5549 18105 5583 18139
rect 8677 18105 8711 18139
rect 11345 18105 11379 18139
rect 13829 18105 13863 18139
rect 7205 18037 7239 18071
rect 9597 18037 9631 18071
rect 11253 18037 11287 18071
rect 12449 18037 12483 18071
rect 12909 18037 12943 18071
rect 13921 18037 13955 18071
rect 3157 17833 3191 17867
rect 5917 17833 5951 17867
rect 6929 17833 6963 17867
rect 12449 17833 12483 17867
rect 13921 17833 13955 17867
rect 14473 17833 14507 17867
rect 1501 17697 1535 17731
rect 2237 17697 2271 17731
rect 2973 17697 3007 17731
rect 4077 17697 4111 17731
rect 4344 17697 4378 17731
rect 5733 17697 5767 17731
rect 6837 17697 6871 17731
rect 7748 17697 7782 17731
rect 9137 17697 9171 17731
rect 10057 17697 10091 17731
rect 10885 17697 10919 17731
rect 11152 17697 11186 17731
rect 1685 17629 1719 17663
rect 2513 17629 2547 17663
rect 3525 17629 3559 17663
rect 7113 17629 7147 17663
rect 7481 17629 7515 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 12808 17765 12842 17799
rect 14289 17697 14323 17731
rect 12541 17629 12575 17663
rect 8861 17561 8895 17595
rect 12265 17561 12299 17595
rect 12449 17561 12483 17595
rect 5457 17493 5491 17527
rect 6469 17493 6503 17527
rect 9689 17493 9723 17527
rect 1777 17289 1811 17323
rect 4629 17289 4663 17323
rect 4721 17289 4755 17323
rect 11713 17289 11747 17323
rect 11989 17289 12023 17323
rect 12449 17289 12483 17323
rect 13645 17289 13679 17323
rect 14197 17289 14231 17323
rect 10057 17221 10091 17255
rect 10241 17221 10275 17255
rect 2421 17153 2455 17187
rect 4721 17153 4755 17187
rect 5457 17153 5491 17187
rect 1593 17085 1627 17119
rect 2145 17085 2179 17119
rect 3249 17085 3283 17119
rect 5365 17085 5399 17119
rect 5917 17085 5951 17119
rect 6653 17085 6687 17119
rect 6837 17085 6871 17119
rect 8677 17085 8711 17119
rect 8944 17085 8978 17119
rect 10333 17153 10367 17187
rect 13001 17153 13035 17187
rect 12173 17085 12207 17119
rect 13461 17085 13495 17119
rect 14013 17085 14047 17119
rect 3516 17017 3550 17051
rect 7104 17017 7138 17051
rect 10241 17017 10275 17051
rect 10578 17017 10612 17051
rect 4905 16949 4939 16983
rect 5273 16949 5307 16983
rect 6101 16949 6135 16983
rect 6469 16949 6503 16983
rect 8217 16949 8251 16983
rect 12817 16949 12851 16983
rect 12909 16949 12943 16983
rect 1869 16745 1903 16779
rect 2973 16745 3007 16779
rect 3341 16745 3375 16779
rect 3433 16745 3467 16779
rect 6009 16745 6043 16779
rect 9137 16745 9171 16779
rect 9965 16745 9999 16779
rect 10425 16745 10459 16779
rect 10977 16745 11011 16779
rect 11437 16745 11471 16779
rect 2513 16677 2547 16711
rect 6530 16677 6564 16711
rect 8493 16677 8527 16711
rect 8585 16677 8619 16711
rect 10333 16677 10367 16711
rect 14565 16677 14599 16711
rect 1685 16609 1719 16643
rect 2237 16609 2271 16643
rect 4077 16609 4111 16643
rect 4629 16609 4663 16643
rect 4896 16609 4930 16643
rect 11345 16609 11379 16643
rect 11989 16609 12023 16643
rect 12889 16609 12923 16643
rect 14289 16609 14323 16643
rect 3617 16541 3651 16575
rect 6285 16541 6319 16575
rect 8677 16541 8711 16575
rect 10517 16541 10551 16575
rect 11621 16541 11655 16575
rect 12633 16541 12667 16575
rect 4261 16473 4295 16507
rect 7665 16473 7699 16507
rect 14013 16473 14047 16507
rect 8125 16405 8159 16439
rect 1593 16201 1627 16235
rect 2973 16201 3007 16235
rect 9045 16201 9079 16235
rect 10057 16201 10091 16235
rect 3985 16133 4019 16167
rect 6377 16133 6411 16167
rect 11069 16133 11103 16167
rect 2605 16065 2639 16099
rect 3617 16065 3651 16099
rect 4629 16065 4663 16099
rect 5825 16065 5859 16099
rect 7481 16065 7515 16099
rect 8401 16065 8435 16099
rect 8585 16065 8619 16099
rect 9689 16065 9723 16099
rect 10701 16065 10735 16099
rect 11621 16065 11655 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 1409 15997 1443 16031
rect 2329 15997 2363 16031
rect 5549 15997 5583 16031
rect 6193 15997 6227 16031
rect 7205 15997 7239 16031
rect 7297 15997 7331 16031
rect 9505 15997 9539 16031
rect 11437 15997 11471 16031
rect 13553 15997 13587 16031
rect 2421 15929 2455 15963
rect 3433 15929 3467 15963
rect 9413 15929 9447 15963
rect 10517 15929 10551 15963
rect 13829 15929 13863 15963
rect 1961 15861 1995 15895
rect 3341 15861 3375 15895
rect 4353 15861 4387 15895
rect 4445 15861 4479 15895
rect 5181 15861 5215 15895
rect 5641 15861 5675 15895
rect 6837 15861 6871 15895
rect 7941 15861 7975 15895
rect 8309 15861 8343 15895
rect 10425 15861 10459 15895
rect 11529 15861 11563 15895
rect 12541 15861 12575 15895
rect 12909 15861 12943 15895
rect 1593 15657 1627 15691
rect 2329 15657 2363 15691
rect 3893 15657 3927 15691
rect 4077 15657 4111 15691
rect 4537 15657 4571 15691
rect 5089 15657 5123 15691
rect 5457 15657 5491 15691
rect 5549 15657 5583 15691
rect 5917 15657 5951 15691
rect 6101 15657 6135 15691
rect 6745 15657 6779 15691
rect 7113 15657 7147 15691
rect 7205 15657 7239 15691
rect 9321 15657 9355 15691
rect 11069 15657 11103 15691
rect 11621 15657 11655 15691
rect 11989 15657 12023 15691
rect 14289 15657 14323 15691
rect 1409 15521 1443 15555
rect 2421 15521 2455 15555
rect 3341 15521 3375 15555
rect 3801 15521 3835 15555
rect 2605 15453 2639 15487
rect 3433 15453 3467 15487
rect 3617 15453 3651 15487
rect 2973 15385 3007 15419
rect 4445 15521 4479 15555
rect 9934 15589 9968 15623
rect 8197 15521 8231 15555
rect 9689 15521 9723 15555
rect 12081 15521 12115 15555
rect 12900 15521 12934 15555
rect 3893 15453 3927 15487
rect 4721 15453 4755 15487
rect 5641 15453 5675 15487
rect 5917 15453 5951 15487
rect 7389 15453 7423 15487
rect 7941 15453 7975 15487
rect 12265 15453 12299 15487
rect 12633 15453 12667 15487
rect 1961 15317 1995 15351
rect 3801 15317 3835 15351
rect 14013 15317 14047 15351
rect 3433 15113 3467 15147
rect 5733 15113 5767 15147
rect 8493 15113 8527 15147
rect 9137 15113 9171 15147
rect 14013 15113 14047 15147
rect 15025 15113 15059 15147
rect 5457 15045 5491 15079
rect 8217 15045 8251 15079
rect 1685 14977 1719 15011
rect 2881 14977 2915 15011
rect 6377 14977 6411 15011
rect 9689 14977 9723 15011
rect 10333 14977 10367 15011
rect 13277 14977 13311 15011
rect 13461 14977 13495 15011
rect 14565 14977 14599 15011
rect 15485 14977 15519 15011
rect 15669 14977 15703 15011
rect 1501 14909 1535 14943
rect 2605 14909 2639 14943
rect 3249 14909 3283 14943
rect 4077 14909 4111 14943
rect 6101 14909 6135 14943
rect 6837 14909 6871 14943
rect 8677 14909 8711 14943
rect 13921 14909 13955 14943
rect 14381 14909 14415 14943
rect 4344 14841 4378 14875
rect 7104 14841 7138 14875
rect 10600 14841 10634 14875
rect 14473 14841 14507 14875
rect 15393 14841 15427 14875
rect 2237 14773 2271 14807
rect 2697 14773 2731 14807
rect 6193 14773 6227 14807
rect 9505 14773 9539 14807
rect 9597 14773 9631 14807
rect 11713 14773 11747 14807
rect 12817 14773 12851 14807
rect 13185 14773 13219 14807
rect 1685 14569 1719 14603
rect 4445 14569 4479 14603
rect 5089 14569 5123 14603
rect 5549 14569 5583 14603
rect 8217 14569 8251 14603
rect 9689 14569 9723 14603
rect 10057 14569 10091 14603
rect 10149 14569 10183 14603
rect 15301 14569 15335 14603
rect 15669 14569 15703 14603
rect 15761 14569 15795 14603
rect 4537 14501 4571 14535
rect 5457 14501 5491 14535
rect 6469 14501 6503 14535
rect 8677 14501 8711 14535
rect 11428 14501 11462 14535
rect 1501 14433 1535 14467
rect 2309 14433 2343 14467
rect 6561 14433 6595 14467
rect 7573 14433 7607 14467
rect 8585 14433 8619 14467
rect 10885 14433 10919 14467
rect 11161 14433 11195 14467
rect 12817 14433 12851 14467
rect 13084 14433 13118 14467
rect 2053 14365 2087 14399
rect 4629 14365 4663 14399
rect 5641 14365 5675 14399
rect 6653 14365 6687 14399
rect 7665 14365 7699 14399
rect 7757 14365 7791 14399
rect 8861 14365 8895 14399
rect 10241 14365 10275 14399
rect 15945 14365 15979 14399
rect 3433 14297 3467 14331
rect 7205 14297 7239 14331
rect 14197 14297 14231 14331
rect 4077 14229 4111 14263
rect 6101 14229 6135 14263
rect 10701 14229 10735 14263
rect 12541 14229 12575 14263
rect 1501 14025 1535 14059
rect 4169 14025 4203 14059
rect 6837 14025 6871 14059
rect 7849 14025 7883 14059
rect 9321 14025 9355 14059
rect 13829 14025 13863 14059
rect 16037 14025 16071 14059
rect 3893 13957 3927 13991
rect 5181 13957 5215 13991
rect 8861 13957 8895 13991
rect 10977 13957 11011 13991
rect 2145 13889 2179 13923
rect 2513 13889 2547 13923
rect 3985 13889 4019 13923
rect 4629 13889 4663 13923
rect 4721 13889 4755 13923
rect 5733 13889 5767 13923
rect 7481 13889 7515 13923
rect 8401 13889 8435 13923
rect 9965 13889 9999 13923
rect 11437 13889 11471 13923
rect 11621 13889 11655 13923
rect 1961 13821 1995 13855
rect 2780 13821 2814 13855
rect 1869 13753 1903 13787
rect 4537 13821 4571 13855
rect 5641 13821 5675 13855
rect 6377 13821 6411 13855
rect 8309 13821 8343 13855
rect 9045 13821 9079 13855
rect 12173 13821 12207 13855
rect 12449 13821 12483 13855
rect 12705 13821 12739 13855
rect 14657 13821 14691 13855
rect 14924 13821 14958 13855
rect 9689 13753 9723 13787
rect 10333 13753 10367 13787
rect 3985 13685 4019 13719
rect 5549 13685 5583 13719
rect 6193 13685 6227 13719
rect 7205 13685 7239 13719
rect 7297 13685 7331 13719
rect 8217 13685 8251 13719
rect 9781 13685 9815 13719
rect 11345 13685 11379 13719
rect 11989 13685 12023 13719
rect 2145 13481 2179 13515
rect 3341 13481 3375 13515
rect 5457 13481 5491 13515
rect 8769 13481 8803 13515
rect 11069 13481 11103 13515
rect 13369 13481 13403 13515
rect 14381 13481 14415 13515
rect 15301 13481 15335 13515
rect 16313 13481 16347 13515
rect 16681 13481 16715 13515
rect 1685 13413 1719 13447
rect 4344 13413 4378 13447
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 2605 13345 2639 13379
rect 3157 13345 3191 13379
rect 5733 13345 5767 13379
rect 6000 13345 6034 13379
rect 7205 13345 7239 13379
rect 7656 13345 7690 13379
rect 9873 13345 9907 13379
rect 10977 13345 11011 13379
rect 11989 13345 12023 13379
rect 13277 13345 13311 13379
rect 14289 13345 14323 13379
rect 15669 13345 15703 13379
rect 2697 13277 2731 13311
rect 4077 13277 4111 13311
rect 7389 13277 7423 13311
rect 10057 13277 10091 13311
rect 11253 13277 11287 13311
rect 11437 13277 11471 13311
rect 12081 13277 12115 13311
rect 12265 13277 12299 13311
rect 13461 13277 13495 13311
rect 14473 13277 14507 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16773 13277 16807 13311
rect 16865 13277 16899 13311
rect 7113 13209 7147 13243
rect 7205 13209 7239 13243
rect 12909 13209 12943 13243
rect 10609 13141 10643 13175
rect 11437 13141 11471 13175
rect 11621 13141 11655 13175
rect 13921 13141 13955 13175
rect 3985 12937 4019 12971
rect 6009 12937 6043 12971
rect 6837 12937 6871 12971
rect 9689 12937 9723 12971
rect 12081 12937 12115 12971
rect 9229 12869 9263 12903
rect 14289 12869 14323 12903
rect 2421 12801 2455 12835
rect 3249 12801 3283 12835
rect 3433 12801 3467 12835
rect 4629 12801 4663 12835
rect 7297 12801 7331 12835
rect 7389 12801 7423 12835
rect 10333 12801 10367 12835
rect 12449 12801 12483 12835
rect 12817 12801 12851 12835
rect 12909 12801 12943 12835
rect 15117 12801 15151 12835
rect 16129 12801 16163 12835
rect 3157 12733 3191 12767
rect 3617 12733 3651 12767
rect 3801 12733 3835 12767
rect 4896 12733 4930 12767
rect 7849 12733 7883 12767
rect 8105 12733 8139 12767
rect 10057 12733 10091 12767
rect 10701 12733 10735 12767
rect 2237 12665 2271 12699
rect 14933 12733 14967 12767
rect 15025 12733 15059 12767
rect 15393 12733 15427 12767
rect 15945 12733 15979 12767
rect 7205 12665 7239 12699
rect 10968 12665 11002 12699
rect 12817 12665 12851 12699
rect 13176 12665 13210 12699
rect 16037 12665 16071 12699
rect 1777 12597 1811 12631
rect 2145 12597 2179 12631
rect 2789 12597 2823 12631
rect 3617 12597 3651 12631
rect 10149 12597 10183 12631
rect 14565 12597 14599 12631
rect 15393 12597 15427 12631
rect 15577 12597 15611 12631
rect 1777 12393 1811 12427
rect 2237 12393 2271 12427
rect 2789 12393 2823 12427
rect 3157 12393 3191 12427
rect 4445 12393 4479 12427
rect 4537 12393 4571 12427
rect 5273 12393 5307 12427
rect 7573 12393 7607 12427
rect 8953 12393 8987 12427
rect 11897 12393 11931 12427
rect 12357 12393 12391 12427
rect 8033 12325 8067 12359
rect 13820 12325 13854 12359
rect 2145 12257 2179 12291
rect 3249 12257 3283 12291
rect 5095 12257 5129 12291
rect 5917 12257 5951 12291
rect 6184 12257 6218 12291
rect 7941 12257 7975 12291
rect 10508 12257 10542 12291
rect 12265 12257 12299 12291
rect 13553 12257 13587 12291
rect 2421 12189 2455 12223
rect 3433 12189 3467 12223
rect 4629 12189 4663 12223
rect 8125 12189 8159 12223
rect 9045 12189 9079 12223
rect 9229 12189 9263 12223
rect 9689 12189 9723 12223
rect 10241 12189 10275 12223
rect 12449 12189 12483 12223
rect 13093 12189 13127 12223
rect 4077 12053 4111 12087
rect 7297 12053 7331 12087
rect 8585 12053 8619 12087
rect 11621 12053 11655 12087
rect 14933 12053 14967 12087
rect 4997 11849 5031 11883
rect 7389 11849 7423 11883
rect 10885 11849 10919 11883
rect 3709 11781 3743 11815
rect 1869 11713 1903 11747
rect 4537 11713 4571 11747
rect 5457 11713 5491 11747
rect 5549 11713 5583 11747
rect 6009 11713 6043 11747
rect 8033 11713 8067 11747
rect 10793 11713 10827 11747
rect 11529 11713 11563 11747
rect 12449 11713 12483 11747
rect 14657 11713 14691 11747
rect 16957 11713 16991 11747
rect 1593 11645 1627 11679
rect 2329 11645 2363 11679
rect 2596 11645 2630 11679
rect 8401 11645 8435 11679
rect 5365 11577 5399 11611
rect 7757 11577 7791 11611
rect 14473 11645 14507 11679
rect 16681 11645 16715 11679
rect 11253 11577 11287 11611
rect 12716 11577 12750 11611
rect 14565 11577 14599 11611
rect 3985 11509 4019 11543
rect 4353 11509 4387 11543
rect 4445 11509 4479 11543
rect 7849 11509 7883 11543
rect 9689 11509 9723 11543
rect 10793 11509 10827 11543
rect 11345 11509 11379 11543
rect 13829 11509 13863 11543
rect 14105 11509 14139 11543
rect 2789 11305 2823 11339
rect 4077 11305 4111 11339
rect 6193 11305 6227 11339
rect 7297 11305 7331 11339
rect 11069 11305 11103 11339
rect 11529 11305 11563 11339
rect 14105 11305 14139 11339
rect 1676 11237 1710 11271
rect 3341 11237 3375 11271
rect 9934 11237 9968 11271
rect 11621 11237 11655 11271
rect 12357 11237 12391 11271
rect 1409 11169 1443 11203
rect 3065 11169 3099 11203
rect 5080 11169 5114 11203
rect 7205 11169 7239 11203
rect 7941 11169 7975 11203
rect 8208 11169 8242 11203
rect 9689 11169 9723 11203
rect 13185 11169 13219 11203
rect 13277 11169 13311 11203
rect 14473 11169 14507 11203
rect 4813 11101 4847 11135
rect 7389 11101 7423 11135
rect 11713 11101 11747 11135
rect 12449 11101 12483 11135
rect 12541 11101 12575 11135
rect 13369 11101 13403 11135
rect 14565 11101 14599 11135
rect 14657 11101 14691 11135
rect 6837 11033 6871 11067
rect 9321 11033 9355 11067
rect 11161 11033 11195 11067
rect 12817 11033 12851 11067
rect 11989 10965 12023 10999
rect 3433 10761 3467 10795
rect 5917 10761 5951 10795
rect 9229 10761 9263 10795
rect 11989 10761 12023 10795
rect 12449 10761 12483 10795
rect 13461 10761 13495 10795
rect 5825 10693 5859 10727
rect 8953 10693 8987 10727
rect 10241 10693 10275 10727
rect 14289 10693 14323 10727
rect 6561 10625 6595 10659
rect 9781 10625 9815 10659
rect 10609 10625 10643 10659
rect 13093 10625 13127 10659
rect 14013 10625 14047 10659
rect 14841 10625 14875 10659
rect 2053 10557 2087 10591
rect 4445 10557 4479 10591
rect 6285 10557 6319 10591
rect 7573 10557 7607 10591
rect 7840 10557 7874 10591
rect 9689 10557 9723 10591
rect 10425 10557 10459 10591
rect 13829 10557 13863 10591
rect 14657 10557 14691 10591
rect 2320 10489 2354 10523
rect 4690 10489 4724 10523
rect 9597 10489 9631 10523
rect 10876 10489 10910 10523
rect 3985 10421 4019 10455
rect 6377 10421 6411 10455
rect 7113 10421 7147 10455
rect 12817 10421 12851 10455
rect 12909 10421 12943 10455
rect 13921 10421 13955 10455
rect 14749 10421 14783 10455
rect 2145 10217 2179 10251
rect 3709 10217 3743 10251
rect 4445 10217 4479 10251
rect 4905 10217 4939 10251
rect 5089 10217 5123 10251
rect 8217 10217 8251 10251
rect 12817 10217 12851 10251
rect 13093 10217 13127 10251
rect 1593 10081 1627 10115
rect 1869 10081 1903 10115
rect 2145 10081 2179 10115
rect 2596 10081 2630 10115
rect 4537 10081 4571 10115
rect 2329 10013 2363 10047
rect 4721 10013 4755 10047
rect 4905 9945 4939 9979
rect 4997 10149 5031 10183
rect 8585 10149 8619 10183
rect 9956 10149 9990 10183
rect 11704 10149 11738 10183
rect 5457 10081 5491 10115
rect 6377 10081 6411 10115
rect 6644 10081 6678 10115
rect 9689 10081 9723 10115
rect 11437 10081 11471 10115
rect 13461 10081 13495 10115
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 8677 10013 8711 10047
rect 8861 10013 8895 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 4077 9877 4111 9911
rect 4997 9877 5031 9911
rect 7757 9877 7791 9911
rect 11069 9877 11103 9911
rect 1961 9605 1995 9639
rect 4997 9605 5031 9639
rect 8125 9605 8159 9639
rect 9597 9605 9631 9639
rect 10609 9605 10643 9639
rect 12449 9605 12483 9639
rect 14289 9605 14323 9639
rect 14473 9605 14507 9639
rect 2605 9537 2639 9571
rect 3525 9537 3559 9571
rect 4445 9537 4479 9571
rect 4629 9537 4663 9571
rect 5641 9537 5675 9571
rect 7389 9537 7423 9571
rect 8677 9537 8711 9571
rect 10149 9537 10183 9571
rect 11161 9537 11195 9571
rect 12909 9537 12943 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 15025 9537 15059 9571
rect 5457 9469 5491 9503
rect 6653 9469 6687 9503
rect 8033 9469 8067 9503
rect 10517 9469 10551 9503
rect 12817 9469 12851 9503
rect 13829 9469 13863 9503
rect 14289 9469 14323 9503
rect 3341 9401 3375 9435
rect 6009 9401 6043 9435
rect 7205 9401 7239 9435
rect 7297 9401 7331 9435
rect 10977 9401 11011 9435
rect 11621 9401 11655 9435
rect 14841 9401 14875 9435
rect 2329 9333 2363 9367
rect 2421 9333 2455 9367
rect 2973 9333 3007 9367
rect 3433 9333 3467 9367
rect 3985 9333 4019 9367
rect 4353 9333 4387 9367
rect 5365 9333 5399 9367
rect 6469 9333 6503 9367
rect 6837 9333 6871 9367
rect 7849 9333 7883 9367
rect 8493 9333 8527 9367
rect 8585 9333 8619 9367
rect 9965 9333 9999 9367
rect 10057 9333 10091 9367
rect 10517 9333 10551 9367
rect 11069 9333 11103 9367
rect 13461 9333 13495 9367
rect 13921 9333 13955 9367
rect 14933 9333 14967 9367
rect 4077 9129 4111 9163
rect 4537 9129 4571 9163
rect 6837 9129 6871 9163
rect 8309 9129 8343 9163
rect 9229 9129 9263 9163
rect 10149 9129 10183 9163
rect 11069 9129 11103 9163
rect 13185 9129 13219 9163
rect 13737 9129 13771 9163
rect 14105 9129 14139 9163
rect 2320 9061 2354 9095
rect 8217 9061 8251 9095
rect 8861 9061 8895 9095
rect 3893 8993 3927 9027
rect 4445 8993 4479 9027
rect 5181 8993 5215 9027
rect 5448 8993 5482 9027
rect 7205 8993 7239 9027
rect 1593 8925 1627 8959
rect 2053 8925 2087 8959
rect 4629 8925 4663 8959
rect 7297 8925 7331 8959
rect 7389 8925 7423 8959
rect 8401 8925 8435 8959
rect 12081 9061 12115 9095
rect 13093 9061 13127 9095
rect 9505 8993 9539 9027
rect 10057 8993 10091 9027
rect 10241 8925 10275 8959
rect 11161 8925 11195 8959
rect 11253 8925 11287 8959
rect 12173 8925 12207 8959
rect 12357 8925 12391 8959
rect 13277 8925 13311 8959
rect 14197 8925 14231 8959
rect 14289 8925 14323 8959
rect 9321 8857 9355 8891
rect 10701 8857 10735 8891
rect 11713 8857 11747 8891
rect 3433 8789 3467 8823
rect 3709 8789 3743 8823
rect 6561 8789 6595 8823
rect 7849 8789 7883 8823
rect 9229 8789 9263 8823
rect 9689 8789 9723 8823
rect 12725 8789 12759 8823
rect 3065 8585 3099 8619
rect 6469 8585 6503 8619
rect 10149 8585 10183 8619
rect 14473 8585 14507 8619
rect 2789 8517 2823 8551
rect 12081 8517 12115 8551
rect 12265 8517 12299 8551
rect 13461 8517 13495 8551
rect 1409 8449 1443 8483
rect 3617 8449 3651 8483
rect 4537 8449 4571 8483
rect 4721 8449 4755 8483
rect 5089 8449 5123 8483
rect 1676 8381 1710 8415
rect 3525 8381 3559 8415
rect 7113 8381 7147 8415
rect 8769 8381 8803 8415
rect 10701 8381 10735 8415
rect 13093 8449 13127 8483
rect 13921 8449 13955 8483
rect 14105 8449 14139 8483
rect 15025 8449 15059 8483
rect 14841 8381 14875 8415
rect 5356 8313 5390 8347
rect 7380 8313 7414 8347
rect 9036 8313 9070 8347
rect 10946 8313 10980 8347
rect 12265 8313 12299 8347
rect 12817 8313 12851 8347
rect 3433 8245 3467 8279
rect 4077 8245 4111 8279
rect 4445 8245 4479 8279
rect 8493 8245 8527 8279
rect 12449 8245 12483 8279
rect 12909 8245 12943 8279
rect 13829 8245 13863 8279
rect 14933 8245 14967 8279
rect 2329 8041 2363 8075
rect 3433 8041 3467 8075
rect 4261 8041 4295 8075
rect 7205 8041 7239 8075
rect 7481 8041 7515 8075
rect 7849 8041 7883 8075
rect 8493 8041 8527 8075
rect 11345 8041 11379 8075
rect 3341 7973 3375 8007
rect 4721 7973 4755 8007
rect 6745 7973 6779 8007
rect 2421 7905 2455 7939
rect 4629 7905 4663 7939
rect 5825 7905 5859 7939
rect 5917 7905 5951 7939
rect 6653 7905 6687 7939
rect 8953 7973 8987 8007
rect 9956 7973 9990 8007
rect 8861 7905 8895 7939
rect 9689 7905 9723 7939
rect 11805 7905 11839 7939
rect 12072 7905 12106 7939
rect 13728 7905 13762 7939
rect 2513 7837 2547 7871
rect 3617 7837 3651 7871
rect 4905 7837 4939 7871
rect 6101 7837 6135 7871
rect 6837 7837 6871 7871
rect 7205 7837 7239 7871
rect 7941 7837 7975 7871
rect 8033 7837 8067 7871
rect 9137 7837 9171 7871
rect 13461 7837 13495 7871
rect 1961 7769 1995 7803
rect 2973 7701 3007 7735
rect 5457 7701 5491 7735
rect 6285 7701 6319 7735
rect 7389 7701 7423 7735
rect 11069 7701 11103 7735
rect 13185 7701 13219 7735
rect 14841 7701 14875 7735
rect 7849 7497 7883 7531
rect 12449 7497 12483 7531
rect 10609 7429 10643 7463
rect 13461 7429 13495 7463
rect 2513 7361 2547 7395
rect 3525 7361 3559 7395
rect 4169 7361 4203 7395
rect 7389 7361 7423 7395
rect 8401 7361 8435 7395
rect 8861 7361 8895 7395
rect 10057 7361 10091 7395
rect 10241 7361 10275 7395
rect 11805 7361 11839 7395
rect 11989 7361 12023 7395
rect 13093 7361 13127 7395
rect 14105 7361 14139 7395
rect 15117 7361 15151 7395
rect 2329 7293 2363 7327
rect 2421 7293 2455 7327
rect 4629 7293 4663 7327
rect 4885 7293 4919 7327
rect 7205 7293 7239 7327
rect 8217 7293 8251 7327
rect 10793 7293 10827 7327
rect 11713 7293 11747 7327
rect 14841 7293 14875 7327
rect 9965 7225 9999 7259
rect 12817 7225 12851 7259
rect 13829 7225 13863 7259
rect 14933 7225 14967 7259
rect 1961 7157 1995 7191
rect 2973 7157 3007 7191
rect 3341 7157 3375 7191
rect 3433 7157 3467 7191
rect 6009 7157 6043 7191
rect 6837 7157 6871 7191
rect 7297 7157 7331 7191
rect 8309 7157 8343 7191
rect 9597 7157 9631 7191
rect 11345 7157 11379 7191
rect 12909 7157 12943 7191
rect 13921 7157 13955 7191
rect 14473 7157 14507 7191
rect 7941 6953 7975 6987
rect 9045 6953 9079 6987
rect 13093 6953 13127 6987
rect 13737 6953 13771 6987
rect 15669 6953 15703 6987
rect 1952 6885 1986 6919
rect 4344 6885 4378 6919
rect 8953 6885 8987 6919
rect 1685 6817 1719 6851
rect 4077 6817 4111 6851
rect 6184 6817 6218 6851
rect 7389 6817 7423 6851
rect 9689 6817 9723 6851
rect 9956 6817 9990 6851
rect 11980 6817 12014 6851
rect 13829 6817 13863 6851
rect 15761 6817 15795 6851
rect 3341 6749 3375 6783
rect 5917 6749 5951 6783
rect 3065 6681 3099 6715
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 9229 6749 9263 6783
rect 11713 6749 11747 6783
rect 13921 6749 13955 6783
rect 14749 6749 14783 6783
rect 15853 6749 15887 6783
rect 11069 6681 11103 6715
rect 13369 6681 13403 6715
rect 5457 6613 5491 6647
rect 7297 6613 7331 6647
rect 7389 6613 7423 6647
rect 7573 6613 7607 6647
rect 8585 6613 8619 6647
rect 15301 6613 15335 6647
rect 2973 6409 3007 6443
rect 3249 6409 3283 6443
rect 5733 6409 5767 6443
rect 9321 6341 9355 6375
rect 3801 6273 3835 6307
rect 4905 6273 4939 6307
rect 6285 6273 6319 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 10977 6273 11011 6307
rect 11989 6273 12023 6307
rect 13001 6273 13035 6307
rect 16405 6273 16439 6307
rect 1593 6205 1627 6239
rect 1860 6205 1894 6239
rect 4629 6205 4663 6239
rect 5457 6205 5491 6239
rect 7941 6205 7975 6239
rect 8208 6205 8242 6239
rect 14197 6205 14231 6239
rect 10793 6137 10827 6171
rect 11713 6137 11747 6171
rect 13461 6137 13495 6171
rect 14464 6137 14498 6171
rect 3617 6069 3651 6103
rect 3709 6069 3743 6103
rect 4261 6069 4295 6103
rect 4721 6069 4755 6103
rect 5273 6069 5307 6103
rect 6101 6069 6135 6103
rect 6193 6069 6227 6103
rect 6837 6069 6871 6103
rect 7205 6069 7239 6103
rect 10333 6069 10367 6103
rect 10701 6069 10735 6103
rect 11345 6069 11379 6103
rect 11805 6069 11839 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 12909 6069 12943 6103
rect 15577 6069 15611 6103
rect 15853 6069 15887 6103
rect 16221 6069 16255 6103
rect 16313 6069 16347 6103
rect 2053 5865 2087 5899
rect 2605 5865 2639 5899
rect 6193 5865 6227 5899
rect 10517 5865 10551 5899
rect 10885 5865 10919 5899
rect 10977 5865 11011 5899
rect 17417 5865 17451 5899
rect 5080 5797 5114 5831
rect 7656 5797 7690 5831
rect 15568 5797 15602 5831
rect 16773 5797 16807 5831
rect 17325 5797 17359 5831
rect 1961 5729 1995 5763
rect 2973 5729 3007 5763
rect 4813 5729 4847 5763
rect 7389 5729 7423 5763
rect 11796 5729 11830 5763
rect 13553 5729 13587 5763
rect 13820 5729 13854 5763
rect 2145 5661 2179 5695
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 11161 5661 11195 5695
rect 11529 5661 11563 5695
rect 15301 5661 15335 5695
rect 18889 5729 18923 5763
rect 17509 5661 17543 5695
rect 19165 5661 19199 5695
rect 1593 5593 1627 5627
rect 12909 5593 12943 5627
rect 16681 5593 16715 5627
rect 16773 5593 16807 5627
rect 8769 5525 8803 5559
rect 14933 5525 14967 5559
rect 16957 5525 16991 5559
rect 6009 5321 6043 5355
rect 8493 5321 8527 5355
rect 11345 5321 11379 5355
rect 14289 5321 14323 5355
rect 14381 5321 14415 5355
rect 16405 5321 16439 5355
rect 13369 5253 13403 5287
rect 3893 5185 3927 5219
rect 8953 5185 8987 5219
rect 9045 5185 9079 5219
rect 10517 5185 10551 5219
rect 11989 5185 12023 5219
rect 14013 5185 14047 5219
rect 14933 5185 14967 5219
rect 15945 5185 15979 5219
rect 16957 5185 16991 5219
rect 2053 5117 2087 5151
rect 2320 5117 2354 5151
rect 3709 5117 3743 5151
rect 4629 5117 4663 5151
rect 6837 5117 6871 5151
rect 7104 5117 7138 5151
rect 12817 5117 12851 5151
rect 14289 5117 14323 5151
rect 14749 5117 14783 5151
rect 14841 5117 14875 5151
rect 15853 5117 15887 5151
rect 19809 5117 19843 5151
rect 4896 5049 4930 5083
rect 8861 5049 8895 5083
rect 13737 5049 13771 5083
rect 15761 5049 15795 5083
rect 16865 5049 16899 5083
rect 3433 4981 3467 5015
rect 8217 4981 8251 5015
rect 9873 4981 9907 5015
rect 10241 4981 10275 5015
rect 10333 4981 10367 5015
rect 11713 4981 11747 5015
rect 11805 4981 11839 5015
rect 13001 4981 13035 5015
rect 13829 4981 13863 5015
rect 15393 4981 15427 5015
rect 16773 4981 16807 5015
rect 19993 4981 20027 5015
rect 1869 4777 1903 4811
rect 6285 4777 6319 4811
rect 7389 4777 7423 4811
rect 10149 4777 10183 4811
rect 12633 4777 12667 4811
rect 12909 4777 12943 4811
rect 14197 4777 14231 4811
rect 15301 4777 15335 4811
rect 4436 4709 4470 4743
rect 7757 4709 7791 4743
rect 14565 4709 14599 4743
rect 2237 4641 2271 4675
rect 2329 4641 2363 4675
rect 3249 4641 3283 4675
rect 4169 4641 4203 4675
rect 6653 4641 6687 4675
rect 8769 4641 8803 4675
rect 8861 4641 8895 4675
rect 10057 4641 10091 4675
rect 11520 4641 11554 4675
rect 13277 4641 13311 4675
rect 14657 4641 14691 4675
rect 15669 4641 15703 4675
rect 15761 4641 15795 4675
rect 17049 4641 17083 4675
rect 17325 4641 17359 4675
rect 17877 4641 17911 4675
rect 2421 4573 2455 4607
rect 3341 4573 3375 4607
rect 3433 4573 3467 4607
rect 6745 4573 6779 4607
rect 6929 4573 6963 4607
rect 7849 4573 7883 4607
rect 8033 4573 8067 4607
rect 8953 4573 8987 4607
rect 10241 4573 10275 4607
rect 10701 4573 10735 4607
rect 11253 4573 11287 4607
rect 13369 4573 13403 4607
rect 13553 4573 13587 4607
rect 14749 4573 14783 4607
rect 15945 4573 15979 4607
rect 5549 4505 5583 4539
rect 8401 4505 8435 4539
rect 2881 4437 2915 4471
rect 9689 4437 9723 4471
rect 18061 4437 18095 4471
rect 3157 4233 3191 4267
rect 5641 4233 5675 4267
rect 7113 4233 7147 4267
rect 8125 4233 8159 4267
rect 9321 4233 9355 4267
rect 13829 4233 13863 4267
rect 4813 4165 4847 4199
rect 10609 4165 10643 4199
rect 10793 4165 10827 4199
rect 10977 4165 11011 4199
rect 14105 4165 14139 4199
rect 6193 4097 6227 4131
rect 7665 4097 7699 4131
rect 8677 4097 8711 4131
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 1777 4029 1811 4063
rect 3433 4029 3467 4063
rect 6101 4029 6135 4063
rect 8493 4029 8527 4063
rect 9689 4029 9723 4063
rect 10425 4029 10459 4063
rect 11437 4097 11471 4131
rect 11529 4097 11563 4131
rect 14657 4097 14691 4131
rect 12449 4029 12483 4063
rect 14473 4029 14507 4063
rect 15117 4029 15151 4063
rect 2044 3961 2078 3995
rect 3700 3961 3734 3995
rect 10793 3961 10827 3995
rect 12716 3961 12750 3995
rect 14565 3961 14599 3995
rect 5181 3893 5215 3927
rect 6009 3893 6043 3927
rect 7481 3893 7515 3927
rect 7573 3893 7607 3927
rect 8585 3893 8619 3927
rect 11345 3893 11379 3927
rect 15301 3893 15335 3927
rect 6193 3689 6227 3723
rect 11161 3689 11195 3723
rect 13093 3689 13127 3723
rect 2044 3621 2078 3655
rect 8953 3621 8987 3655
rect 10048 3621 10082 3655
rect 11682 3621 11716 3655
rect 4169 3553 4203 3587
rect 4436 3553 4470 3587
rect 7021 3553 7055 3587
rect 7288 3553 7322 3587
rect 8677 3553 8711 3587
rect 13461 3553 13495 3587
rect 14105 3553 14139 3587
rect 15301 3553 15335 3587
rect 16037 3553 16071 3587
rect 1777 3485 1811 3519
rect 3433 3485 3467 3519
rect 6285 3485 6319 3519
rect 6377 3485 6411 3519
rect 9781 3485 9815 3519
rect 11437 3485 11471 3519
rect 13553 3485 13587 3519
rect 13645 3485 13679 3519
rect 14289 3485 14323 3519
rect 15577 3485 15611 3519
rect 5825 3417 5859 3451
rect 12817 3417 12851 3451
rect 3157 3349 3191 3383
rect 5549 3349 5583 3383
rect 8401 3349 8435 3383
rect 16221 3349 16255 3383
rect 2329 3145 2363 3179
rect 3709 3145 3743 3179
rect 4721 3145 4755 3179
rect 5733 3145 5767 3179
rect 9597 3145 9631 3179
rect 12449 3145 12483 3179
rect 13369 3145 13403 3179
rect 14381 3145 14415 3179
rect 2973 3009 3007 3043
rect 4261 3009 4295 3043
rect 5273 3009 5307 3043
rect 6377 3009 6411 3043
rect 7481 3009 7515 3043
rect 7573 3009 7607 3043
rect 10425 3009 10459 3043
rect 11437 3009 11471 3043
rect 13093 3009 13127 3043
rect 2697 2941 2731 2975
rect 5181 2941 5215 2975
rect 8217 2941 8251 2975
rect 10241 2941 10275 2975
rect 12817 2941 12851 2975
rect 14933 3077 14967 3111
rect 18521 3077 18555 3111
rect 13737 3009 13771 3043
rect 13461 2941 13495 2975
rect 14197 2941 14231 2975
rect 14749 2941 14783 2975
rect 15301 2941 15335 2975
rect 16129 2941 16163 2975
rect 17049 2941 17083 2975
rect 18337 2941 18371 2975
rect 18889 2941 18923 2975
rect 4077 2873 4111 2907
rect 5089 2873 5123 2907
rect 6101 2873 6135 2907
rect 8462 2873 8496 2907
rect 11345 2873 11379 2907
rect 13369 2873 13403 2907
rect 2789 2805 2823 2839
rect 4169 2805 4203 2839
rect 6193 2805 6227 2839
rect 7021 2805 7055 2839
rect 7389 2805 7423 2839
rect 9873 2805 9907 2839
rect 10333 2805 10367 2839
rect 10885 2805 10919 2839
rect 11253 2805 11287 2839
rect 12909 2805 12943 2839
rect 15485 2805 15519 2839
rect 16313 2805 16347 2839
rect 17233 2805 17267 2839
rect 19073 2805 19107 2839
rect 2237 2601 2271 2635
rect 2605 2601 2639 2635
rect 4077 2601 4111 2635
rect 5365 2601 5399 2635
rect 7573 2601 7607 2635
rect 9045 2601 9079 2635
rect 9137 2601 9171 2635
rect 11161 2601 11195 2635
rect 11989 2601 12023 2635
rect 13553 2601 13587 2635
rect 2697 2533 2731 2567
rect 10149 2533 10183 2567
rect 4445 2465 4479 2499
rect 5733 2465 5767 2499
rect 7941 2465 7975 2499
rect 10241 2465 10275 2499
rect 11805 2465 11839 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 14013 2465 14047 2499
rect 14749 2465 14783 2499
rect 15669 2465 15703 2499
rect 16589 2465 16623 2499
rect 17509 2465 17543 2499
rect 2881 2397 2915 2431
rect 4537 2397 4571 2431
rect 4629 2397 4663 2431
rect 5825 2397 5859 2431
rect 6009 2397 6043 2431
rect 8033 2397 8067 2431
rect 8217 2397 8251 2431
rect 9321 2397 9355 2431
rect 10333 2397 10367 2431
rect 11253 2397 11287 2431
rect 11437 2397 11471 2431
rect 12817 2397 12851 2431
rect 8677 2329 8711 2363
rect 10793 2329 10827 2363
rect 14197 2329 14231 2363
rect 9781 2261 9815 2295
rect 14933 2261 14967 2295
rect 15853 2261 15887 2295
rect 16773 2261 16807 2295
rect 17693 2261 17727 2295
<< metal1 >>
rect 3878 20544 3884 20596
rect 3936 20584 3942 20596
rect 6362 20584 6368 20596
rect 3936 20556 6368 20584
rect 3936 20544 3942 20556
rect 6362 20544 6368 20556
rect 6420 20544 6426 20596
rect 4430 20204 4436 20256
rect 4488 20244 4494 20256
rect 8938 20244 8944 20256
rect 4488 20216 8944 20244
rect 4488 20204 4494 20216
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4430 20040 4436 20052
rect 4212 20012 4436 20040
rect 4212 20000 4218 20012
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 5166 20040 5172 20052
rect 4571 20012 5172 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 10689 20043 10747 20049
rect 10689 20009 10701 20043
rect 10735 20040 10747 20043
rect 12434 20040 12440 20052
rect 10735 20012 12440 20040
rect 10735 20009 10747 20012
rect 10689 20003 10747 20009
rect 12434 20000 12440 20012
rect 12492 20000 12498 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 12894 20040 12900 20052
rect 12851 20012 12900 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13354 20040 13360 20052
rect 13315 20012 13360 20040
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 14369 20043 14427 20049
rect 14369 20009 14381 20043
rect 14415 20040 14427 20043
rect 14550 20040 14556 20052
rect 14415 20012 14556 20040
rect 14415 20009 14427 20012
rect 14369 20003 14427 20009
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20040 14979 20043
rect 15194 20040 15200 20052
rect 14967 20012 15200 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15654 20040 15660 20052
rect 15615 20012 15660 20040
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 16209 20043 16267 20049
rect 16209 20009 16221 20043
rect 16255 20040 16267 20043
rect 16574 20040 16580 20052
rect 16255 20012 16580 20040
rect 16255 20009 16267 20012
rect 16209 20003 16267 20009
rect 16574 20000 16580 20012
rect 16632 20000 16638 20052
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 17954 20040 17960 20052
rect 17359 20012 17960 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 3329 19975 3387 19981
rect 1688 19944 3280 19972
rect 1688 19913 1716 19944
rect 1673 19907 1731 19913
rect 1673 19873 1685 19907
rect 1719 19873 1731 19907
rect 1673 19867 1731 19873
rect 2225 19907 2283 19913
rect 2225 19873 2237 19907
rect 2271 19904 2283 19907
rect 2866 19904 2872 19916
rect 2271 19876 2872 19904
rect 2271 19873 2283 19876
rect 2225 19867 2283 19873
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 3050 19904 3056 19916
rect 3011 19876 3056 19904
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 3252 19904 3280 19944
rect 3329 19941 3341 19975
rect 3375 19972 3387 19975
rect 5810 19972 5816 19984
rect 3375 19944 5816 19972
rect 3375 19941 3387 19944
rect 3329 19935 3387 19941
rect 5810 19932 5816 19944
rect 5868 19932 5874 19984
rect 6914 19932 6920 19984
rect 6972 19972 6978 19984
rect 9125 19975 9183 19981
rect 9125 19972 9137 19975
rect 6972 19944 9137 19972
rect 6972 19932 6978 19944
rect 9125 19941 9137 19944
rect 9171 19941 9183 19975
rect 9125 19935 9183 19941
rect 11517 19975 11575 19981
rect 11517 19941 11529 19975
rect 11563 19972 11575 19975
rect 11563 19944 12664 19972
rect 11563 19941 11575 19944
rect 11517 19935 11575 19941
rect 5258 19904 5264 19916
rect 3252 19876 5264 19904
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5436 19907 5494 19913
rect 5436 19873 5448 19907
rect 5482 19904 5494 19907
rect 6454 19904 6460 19916
rect 5482 19876 6460 19904
rect 5482 19873 5494 19876
rect 5436 19867 5494 19873
rect 6454 19864 6460 19876
rect 6512 19864 6518 19916
rect 7101 19907 7159 19913
rect 7101 19873 7113 19907
rect 7147 19873 7159 19907
rect 7101 19867 7159 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 8754 19904 8760 19916
rect 8251 19876 8760 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19805 2467 19839
rect 4706 19836 4712 19848
rect 4667 19808 4712 19836
rect 2409 19799 2467 19805
rect 2424 19768 2452 19799
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 4982 19796 4988 19848
rect 5040 19836 5046 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 5040 19808 5181 19836
rect 5040 19796 5046 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 7116 19768 7144 19867
rect 8754 19864 8760 19876
rect 8812 19864 8818 19916
rect 8849 19907 8907 19913
rect 8849 19873 8861 19907
rect 8895 19873 8907 19907
rect 10594 19904 10600 19916
rect 10555 19876 10600 19904
rect 8849 19867 8907 19873
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 7285 19839 7343 19845
rect 7285 19836 7297 19839
rect 7248 19808 7297 19836
rect 7248 19796 7254 19808
rect 7285 19805 7297 19808
rect 7331 19805 7343 19839
rect 8294 19836 8300 19848
rect 8255 19808 8300 19836
rect 7285 19799 7343 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 8389 19839 8447 19845
rect 8389 19805 8401 19839
rect 8435 19805 8447 19839
rect 8389 19799 8447 19805
rect 7837 19771 7895 19777
rect 7837 19768 7849 19771
rect 2424 19740 4384 19768
rect 7116 19740 7849 19768
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 4062 19700 4068 19712
rect 4023 19672 4068 19700
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 4356 19700 4384 19740
rect 7837 19737 7849 19740
rect 7883 19737 7895 19771
rect 7837 19731 7895 19737
rect 8202 19728 8208 19780
rect 8260 19768 8266 19780
rect 8404 19768 8432 19799
rect 8478 19796 8484 19848
rect 8536 19836 8542 19848
rect 8864 19836 8892 19867
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11241 19907 11299 19913
rect 11241 19904 11253 19907
rect 11112 19876 11253 19904
rect 11112 19864 11118 19876
rect 11241 19873 11253 19876
rect 11287 19873 11299 19907
rect 11241 19867 11299 19873
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 12250 19904 12256 19916
rect 12023 19876 12256 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 12636 19913 12664 19944
rect 12627 19907 12685 19913
rect 12627 19873 12639 19907
rect 12673 19873 12685 19907
rect 12627 19867 12685 19873
rect 13173 19907 13231 19913
rect 13173 19873 13185 19907
rect 13219 19904 13231 19907
rect 13814 19904 13820 19916
rect 13219 19876 13820 19904
rect 13219 19873 13231 19876
rect 13173 19867 13231 19873
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 14182 19904 14188 19916
rect 14143 19876 14188 19904
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14516 19876 14749 19904
rect 14516 19864 14522 19876
rect 14737 19873 14749 19876
rect 14783 19873 14795 19907
rect 15470 19904 15476 19916
rect 15431 19876 15476 19904
rect 14737 19867 14795 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 16025 19907 16083 19913
rect 16025 19904 16037 19907
rect 15620 19876 16037 19904
rect 15620 19864 15626 19876
rect 16025 19873 16037 19876
rect 16071 19873 16083 19907
rect 17126 19904 17132 19916
rect 17087 19876 17132 19904
rect 16025 19867 16083 19873
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 8536 19808 8892 19836
rect 8536 19796 8542 19808
rect 9674 19796 9680 19848
rect 9732 19836 9738 19848
rect 9769 19839 9827 19845
rect 9769 19836 9781 19839
rect 9732 19808 9781 19836
rect 9732 19796 9738 19808
rect 9769 19805 9781 19808
rect 9815 19805 9827 19839
rect 9769 19799 9827 19805
rect 10873 19839 10931 19845
rect 10873 19805 10885 19839
rect 10919 19836 10931 19839
rect 10962 19836 10968 19848
rect 10919 19808 10968 19836
rect 10919 19805 10931 19808
rect 10873 19799 10931 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 8260 19740 8432 19768
rect 12161 19771 12219 19777
rect 8260 19728 8266 19740
rect 12161 19737 12173 19771
rect 12207 19768 12219 19771
rect 19334 19768 19340 19780
rect 12207 19740 19340 19768
rect 12207 19737 12219 19740
rect 12161 19731 12219 19737
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 5350 19700 5356 19712
rect 4356 19672 5356 19700
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6549 19703 6607 19709
rect 6549 19700 6561 19703
rect 5592 19672 6561 19700
rect 5592 19660 5598 19672
rect 6549 19669 6561 19672
rect 6595 19669 6607 19703
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 6549 19663 6607 19669
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 2774 19496 2780 19508
rect 2608 19468 2780 19496
rect 1581 19295 1639 19301
rect 1581 19261 1593 19295
rect 1627 19261 1639 19295
rect 1581 19255 1639 19261
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 2608 19292 2636 19468
rect 2774 19456 2780 19468
rect 2832 19456 2838 19508
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 4028 19468 7021 19496
rect 4028 19456 4034 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 6187 19332 7052 19360
rect 2179 19264 2636 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 1596 19224 1624 19255
rect 2682 19252 2688 19304
rect 2740 19292 2746 19304
rect 2961 19295 3019 19301
rect 2961 19292 2973 19295
rect 2740 19264 2973 19292
rect 2740 19252 2746 19264
rect 2961 19261 2973 19264
rect 3007 19261 3019 19295
rect 2961 19255 3019 19261
rect 3228 19295 3286 19301
rect 3228 19261 3240 19295
rect 3274 19292 3286 19295
rect 4706 19292 4712 19304
rect 3274 19264 4712 19292
rect 3274 19261 3286 19264
rect 3228 19255 3286 19261
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 4982 19252 4988 19304
rect 5040 19292 5046 19304
rect 5077 19295 5135 19301
rect 5077 19292 5089 19295
rect 5040 19264 5089 19292
rect 5040 19252 5046 19264
rect 5077 19261 5089 19264
rect 5123 19292 5135 19295
rect 6187 19292 6215 19332
rect 5123 19264 6215 19292
rect 6825 19295 6883 19301
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 6914 19292 6920 19304
rect 6871 19264 6920 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7024 19292 7052 19332
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11238 19360 11244 19372
rect 11112 19332 11244 19360
rect 11112 19320 11118 19332
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12023 19332 12572 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 7282 19292 7288 19304
rect 7024 19264 7288 19292
rect 7282 19252 7288 19264
rect 7340 19292 7346 19304
rect 7377 19295 7435 19301
rect 7377 19292 7389 19295
rect 7340 19264 7389 19292
rect 7340 19252 7346 19264
rect 7377 19261 7389 19264
rect 7423 19261 7435 19295
rect 9033 19295 9091 19301
rect 9033 19292 9045 19295
rect 7377 19255 7435 19261
rect 7484 19264 9045 19292
rect 2222 19224 2228 19236
rect 1596 19196 2228 19224
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 2409 19227 2467 19233
rect 2409 19193 2421 19227
rect 2455 19224 2467 19227
rect 2455 19196 3280 19224
rect 2455 19193 2467 19196
rect 2409 19187 2467 19193
rect 1762 19156 1768 19168
rect 1723 19128 1768 19156
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 3252 19156 3280 19196
rect 3326 19184 3332 19236
rect 3384 19224 3390 19236
rect 4617 19227 4675 19233
rect 4617 19224 4629 19227
rect 3384 19196 4629 19224
rect 3384 19184 3390 19196
rect 4617 19193 4629 19196
rect 4663 19193 4675 19227
rect 4617 19187 4675 19193
rect 5344 19227 5402 19233
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 5718 19224 5724 19236
rect 5390 19196 5724 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 6638 19184 6644 19236
rect 6696 19224 6702 19236
rect 7484 19224 7512 19264
rect 9033 19261 9045 19264
rect 9079 19261 9091 19295
rect 9033 19255 9091 19261
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9582 19292 9588 19304
rect 9539 19264 9588 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9582 19252 9588 19264
rect 9640 19292 9646 19304
rect 11882 19292 11888 19304
rect 9640 19264 11888 19292
rect 9640 19252 9646 19264
rect 11882 19252 11888 19264
rect 11940 19292 11946 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11940 19264 12449 19292
rect 11940 19252 11946 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12544 19292 12572 19332
rect 12544 19264 12756 19292
rect 12437 19255 12495 19261
rect 6696 19196 7512 19224
rect 7644 19227 7702 19233
rect 6696 19184 6702 19196
rect 7644 19193 7656 19227
rect 7690 19224 7702 19227
rect 9398 19224 9404 19236
rect 7690 19196 9404 19224
rect 7690 19193 7702 19196
rect 7644 19187 7702 19193
rect 9398 19184 9404 19196
rect 9456 19184 9462 19236
rect 9760 19227 9818 19233
rect 9760 19193 9772 19227
rect 9806 19224 9818 19227
rect 10962 19224 10968 19236
rect 9806 19196 10968 19224
rect 9806 19193 9818 19196
rect 9760 19187 9818 19193
rect 10962 19184 10968 19196
rect 11020 19224 11026 19236
rect 12728 19233 12756 19264
rect 13998 19252 14004 19304
rect 14056 19292 14062 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 14056 19264 14105 19292
rect 14056 19252 14062 19264
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14093 19255 14151 19261
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19292 14979 19295
rect 16022 19292 16028 19304
rect 14967 19264 15516 19292
rect 15983 19264 16028 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 12704 19227 12762 19233
rect 11020 19196 12664 19224
rect 11020 19184 11026 19196
rect 3418 19156 3424 19168
rect 3252 19128 3424 19156
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 3602 19116 3608 19168
rect 3660 19156 3666 19168
rect 4341 19159 4399 19165
rect 4341 19156 4353 19159
rect 3660 19128 4353 19156
rect 3660 19116 3666 19128
rect 4341 19125 4353 19128
rect 4387 19125 4399 19159
rect 6454 19156 6460 19168
rect 6415 19128 6460 19156
rect 4341 19119 4399 19125
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 8757 19159 8815 19165
rect 8757 19156 8769 19159
rect 8260 19128 8769 19156
rect 8260 19116 8266 19128
rect 8757 19125 8769 19128
rect 8803 19125 8815 19159
rect 10870 19156 10876 19168
rect 10831 19128 10876 19156
rect 8757 19119 8815 19125
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11333 19159 11391 19165
rect 11333 19156 11345 19159
rect 11112 19128 11345 19156
rect 11112 19116 11118 19128
rect 11333 19125 11345 19128
rect 11379 19125 11391 19159
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 11333 19119 11391 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11793 19159 11851 19165
rect 11793 19125 11805 19159
rect 11839 19156 11851 19159
rect 12526 19156 12532 19168
rect 11839 19128 12532 19156
rect 11839 19125 11851 19128
rect 11793 19119 11851 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 12636 19156 12664 19196
rect 12704 19193 12716 19227
rect 12750 19224 12762 19227
rect 13262 19224 13268 19236
rect 12750 19196 13268 19224
rect 12750 19193 12762 19196
rect 12704 19187 12762 19193
rect 13262 19184 13268 19196
rect 13320 19184 13326 19236
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 12636 19128 13829 19156
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 14274 19156 14280 19168
rect 14235 19128 14280 19156
rect 13817 19119 13875 19125
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 15488 19156 15516 19264
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16574 19292 16580 19304
rect 16535 19264 16580 19292
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 16850 19252 16856 19304
rect 16908 19292 16914 19304
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 16908 19264 17141 19292
rect 16908 19252 16914 19264
rect 17129 19261 17141 19264
rect 17175 19261 17187 19295
rect 17129 19255 17187 19261
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17276 19264 18061 19292
rect 17276 19252 17282 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18598 19292 18604 19304
rect 18559 19264 18604 19292
rect 18049 19255 18107 19261
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 18748 19264 19349 19292
rect 18748 19252 18754 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19337 19255 19395 19261
rect 15565 19227 15623 19233
rect 15565 19193 15577 19227
rect 15611 19224 15623 19227
rect 15746 19224 15752 19236
rect 15611 19196 15752 19224
rect 15611 19193 15623 19196
rect 15565 19187 15623 19193
rect 15746 19184 15752 19196
rect 15804 19184 15810 19236
rect 22094 19224 22100 19236
rect 15948 19196 22100 19224
rect 15948 19156 15976 19196
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 15488 19128 15976 19156
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16209 19159 16267 19165
rect 16209 19156 16221 19159
rect 16172 19128 16221 19156
rect 16172 19116 16178 19128
rect 16209 19125 16221 19128
rect 16255 19125 16267 19159
rect 16209 19119 16267 19125
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 17034 19156 17040 19168
rect 16807 19128 17040 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17313 19159 17371 19165
rect 17313 19125 17325 19159
rect 17359 19156 17371 19159
rect 17494 19156 17500 19168
rect 17359 19128 17500 19156
rect 17359 19125 17371 19128
rect 17313 19119 17371 19125
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18506 19156 18512 19168
rect 18279 19128 18512 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18785 19159 18843 19165
rect 18785 19125 18797 19159
rect 18831 19156 18843 19159
rect 18874 19156 18880 19168
rect 18831 19128 18880 19156
rect 18831 19125 18843 19128
rect 18785 19119 18843 19125
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 19521 19159 19579 19165
rect 19521 19125 19533 19159
rect 19567 19156 19579 19159
rect 20254 19156 20260 19168
rect 19567 19128 20260 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 2961 18955 3019 18961
rect 2961 18952 2973 18955
rect 2924 18924 2973 18952
rect 2924 18912 2930 18924
rect 2961 18921 2973 18924
rect 3007 18921 3019 18955
rect 3326 18952 3332 18964
rect 3287 18924 3332 18952
rect 2961 18915 3019 18921
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 4062 18952 4068 18964
rect 3467 18924 4068 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 5442 18952 5448 18964
rect 4172 18924 5448 18952
rect 4172 18884 4200 18924
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5718 18912 5724 18964
rect 5776 18952 5782 18964
rect 6549 18955 6607 18961
rect 6549 18952 6561 18955
rect 5776 18924 6561 18952
rect 5776 18912 5782 18924
rect 6549 18921 6561 18924
rect 6595 18921 6607 18955
rect 6549 18915 6607 18921
rect 8665 18955 8723 18961
rect 8665 18921 8677 18955
rect 8711 18921 8723 18955
rect 8665 18915 8723 18921
rect 2608 18856 4200 18884
rect 4433 18887 4491 18893
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 2314 18816 2320 18828
rect 2275 18788 2320 18816
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2608 18757 2636 18856
rect 4433 18853 4445 18887
rect 4479 18884 4491 18887
rect 6825 18887 6883 18893
rect 6825 18884 6837 18887
rect 4479 18856 6837 18884
rect 4479 18853 4491 18856
rect 4433 18847 4491 18853
rect 6825 18853 6837 18856
rect 6871 18853 6883 18887
rect 6825 18847 6883 18853
rect 7552 18887 7610 18893
rect 7552 18853 7564 18887
rect 7598 18884 7610 18887
rect 8202 18884 8208 18896
rect 7598 18856 8208 18884
rect 7598 18853 7610 18856
rect 7552 18847 7610 18853
rect 8202 18844 8208 18856
rect 8260 18844 8266 18896
rect 2792 18788 3740 18816
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18717 2651 18751
rect 2792 18748 2820 18788
rect 3602 18748 3608 18760
rect 2593 18711 2651 18717
rect 2700 18720 2820 18748
rect 3563 18720 3608 18748
rect 1578 18680 1584 18692
rect 1539 18652 1584 18680
rect 1578 18640 1584 18652
rect 1636 18640 1642 18692
rect 2424 18680 2452 18711
rect 2700 18680 2728 18720
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 3712 18748 3740 18788
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 4890 18816 4896 18828
rect 3844 18788 4896 18816
rect 3844 18776 3850 18788
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 4982 18776 4988 18828
rect 5040 18816 5046 18828
rect 5442 18825 5448 18828
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 5040 18788 5181 18816
rect 5040 18776 5046 18788
rect 5169 18785 5181 18788
rect 5215 18785 5227 18819
rect 5436 18816 5448 18825
rect 5355 18788 5448 18816
rect 5169 18779 5227 18785
rect 5436 18779 5448 18788
rect 5500 18816 5506 18828
rect 8680 18816 8708 18915
rect 8754 18912 8760 18964
rect 8812 18952 8818 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8812 18924 8953 18952
rect 8812 18912 8818 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 10410 18952 10416 18964
rect 9364 18924 10416 18952
rect 9364 18912 9370 18924
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 11974 18912 11980 18964
rect 12032 18952 12038 18964
rect 12802 18952 12808 18964
rect 12032 18924 12808 18952
rect 12032 18912 12038 18924
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 13262 18952 13268 18964
rect 13223 18924 13268 18952
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 21174 18952 21180 18964
rect 19392 18924 21180 18952
rect 19392 18912 19398 18924
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 8846 18844 8852 18896
rect 8904 18884 8910 18896
rect 9944 18887 10002 18893
rect 9944 18884 9956 18887
rect 8904 18856 9956 18884
rect 8904 18844 8910 18856
rect 9944 18853 9956 18856
rect 9990 18884 10002 18887
rect 10870 18884 10876 18896
rect 9990 18856 10876 18884
rect 9990 18853 10002 18856
rect 9944 18847 10002 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11606 18844 11612 18896
rect 11664 18884 11670 18896
rect 12894 18884 12900 18896
rect 11664 18856 12900 18884
rect 11664 18844 11670 18856
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 13814 18884 13820 18896
rect 13775 18856 13820 18884
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 14553 18887 14611 18893
rect 14553 18884 14565 18887
rect 14240 18856 14565 18884
rect 14240 18844 14246 18856
rect 14553 18853 14565 18856
rect 14599 18853 14611 18887
rect 15562 18884 15568 18896
rect 15523 18856 15568 18884
rect 14553 18847 14611 18853
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 18690 18884 18696 18896
rect 18651 18856 18696 18884
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 11054 18816 11060 18828
rect 5500 18788 8708 18816
rect 8772 18788 11060 18816
rect 5442 18776 5448 18779
rect 5500 18776 5506 18788
rect 4338 18748 4344 18760
rect 3712 18720 4344 18748
rect 4338 18708 4344 18720
rect 4396 18708 4402 18760
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 2424 18652 2728 18680
rect 3050 18640 3056 18692
rect 3108 18680 3114 18692
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3108 18652 4077 18680
rect 3108 18640 3114 18652
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4065 18643 4123 18649
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 4154 18612 4160 18624
rect 1995 18584 4160 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4540 18612 4568 18711
rect 4614 18708 4620 18760
rect 4672 18748 4678 18760
rect 7282 18748 7288 18760
rect 4672 18720 4717 18748
rect 7243 18720 7288 18748
rect 4672 18708 4678 18720
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 5074 18680 5080 18692
rect 4816 18652 5080 18680
rect 4816 18612 4844 18652
rect 5074 18640 5080 18652
rect 5132 18640 5138 18692
rect 4540 18584 4844 18612
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 8772 18612 8800 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11146 18776 11152 18828
rect 11204 18776 11210 18828
rect 11333 18819 11391 18825
rect 11333 18785 11345 18819
rect 11379 18785 11391 18819
rect 11882 18816 11888 18828
rect 11843 18788 11888 18816
rect 11333 18779 11391 18785
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 9640 18720 9689 18748
rect 9640 18708 9646 18720
rect 9677 18717 9689 18720
rect 9723 18717 9735 18751
rect 9677 18711 9735 18717
rect 11164 18624 11192 18776
rect 11348 18748 11376 18779
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12152 18819 12210 18825
rect 12152 18785 12164 18819
rect 12198 18816 12210 18819
rect 12986 18816 12992 18828
rect 12198 18788 12992 18816
rect 12198 18785 12210 18788
rect 12152 18779 12210 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13078 18776 13084 18828
rect 13136 18816 13142 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 13136 18788 13553 18816
rect 13136 18776 13142 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18785 14335 18819
rect 15286 18816 15292 18828
rect 15247 18788 15292 18816
rect 14277 18779 14335 18785
rect 11790 18748 11796 18760
rect 11348 18720 11796 18748
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 14292 18748 14320 18779
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 18012 18788 18429 18816
rect 18012 18776 18018 18788
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 15562 18748 15568 18760
rect 14292 18720 15568 18748
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 4948 18584 8800 18612
rect 4948 18572 4954 18584
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 11057 18615 11115 18621
rect 11057 18612 11069 18615
rect 9456 18584 11069 18612
rect 9456 18572 9462 18584
rect 11057 18581 11069 18584
rect 11103 18581 11115 18615
rect 11057 18575 11115 18581
rect 11146 18572 11152 18624
rect 11204 18572 11210 18624
rect 11517 18615 11575 18621
rect 11517 18581 11529 18615
rect 11563 18612 11575 18615
rect 19794 18612 19800 18624
rect 11563 18584 19800 18612
rect 11563 18581 11575 18584
rect 11517 18575 11575 18581
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 198 18368 204 18420
rect 256 18408 262 18420
rect 2590 18408 2596 18420
rect 256 18380 2596 18408
rect 256 18368 262 18380
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 2832 18380 4476 18408
rect 2832 18368 2838 18380
rect 1670 18340 1676 18352
rect 1631 18312 1676 18340
rect 1670 18300 1676 18312
rect 1728 18300 1734 18352
rect 2314 18300 2320 18352
rect 2372 18340 2378 18352
rect 3050 18340 3056 18352
rect 2372 18312 3056 18340
rect 2372 18300 2378 18312
rect 3050 18300 3056 18312
rect 3108 18300 3114 18352
rect 4448 18340 4476 18380
rect 4706 18368 4712 18420
rect 4764 18408 4770 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 4764 18380 4905 18408
rect 4764 18368 4770 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 6825 18411 6883 18417
rect 6825 18408 6837 18411
rect 5132 18380 6837 18408
rect 5132 18368 5138 18380
rect 6825 18377 6837 18380
rect 6871 18377 6883 18411
rect 6825 18371 6883 18377
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 8478 18408 8484 18420
rect 8251 18380 8484 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 8628 18380 10885 18408
rect 8628 18368 8634 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 14645 18411 14703 18417
rect 14645 18377 14657 18411
rect 14691 18408 14703 18411
rect 21634 18408 21640 18420
rect 14691 18380 21640 18408
rect 14691 18377 14703 18380
rect 14645 18371 14703 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 5169 18343 5227 18349
rect 5169 18340 5181 18343
rect 4448 18312 5181 18340
rect 5169 18309 5181 18312
rect 5215 18309 5227 18343
rect 6362 18340 6368 18352
rect 6323 18312 6368 18340
rect 5169 18303 5227 18309
rect 6362 18300 6368 18312
rect 6420 18300 6426 18352
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 6512 18312 7420 18340
rect 6512 18300 6518 18312
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 1504 18244 2237 18272
rect 1504 18213 1532 18244
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 2682 18232 2688 18284
rect 2740 18272 2746 18284
rect 3513 18275 3571 18281
rect 3513 18272 3525 18275
rect 2740 18244 3525 18272
rect 2740 18232 2746 18244
rect 3513 18241 3525 18244
rect 3559 18241 3571 18275
rect 5718 18272 5724 18284
rect 5679 18244 5724 18272
rect 3513 18235 3571 18241
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 7006 18232 7012 18284
rect 7064 18272 7070 18284
rect 7392 18281 7420 18312
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 9217 18343 9275 18349
rect 9217 18340 9229 18343
rect 8352 18312 9229 18340
rect 8352 18300 8358 18312
rect 9217 18309 9229 18312
rect 9263 18309 9275 18343
rect 9674 18340 9680 18352
rect 9217 18303 9275 18309
rect 9324 18312 9680 18340
rect 7285 18275 7343 18281
rect 7285 18272 7297 18275
rect 7064 18244 7297 18272
rect 7064 18232 7070 18244
rect 7285 18241 7297 18244
rect 7331 18241 7343 18275
rect 7285 18235 7343 18241
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 8846 18272 8852 18284
rect 8807 18244 8852 18272
rect 7377 18235 7435 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 1489 18207 1547 18213
rect 1489 18173 1501 18207
rect 1535 18173 1547 18207
rect 1489 18167 1547 18173
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 2777 18207 2835 18213
rect 2777 18173 2789 18207
rect 2823 18204 2835 18207
rect 3780 18207 3838 18213
rect 2823 18176 3740 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 2056 18068 2084 18167
rect 2222 18096 2228 18148
rect 2280 18136 2286 18148
rect 3053 18139 3111 18145
rect 3053 18136 3065 18139
rect 2280 18108 3065 18136
rect 2280 18096 2286 18108
rect 3053 18105 3065 18108
rect 3099 18105 3111 18139
rect 3053 18099 3111 18105
rect 3326 18068 3332 18080
rect 2056 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 3712 18068 3740 18176
rect 3780 18173 3792 18207
rect 3826 18204 3838 18207
rect 4062 18204 4068 18216
rect 3826 18176 4068 18204
rect 3826 18173 3838 18176
rect 3780 18167 3838 18173
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 5629 18207 5687 18213
rect 5629 18204 5641 18207
rect 4212 18176 5641 18204
rect 4212 18164 4218 18176
rect 5629 18173 5641 18176
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 7190 18204 7196 18216
rect 6227 18176 7196 18204
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 9324 18204 9352 18312
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 11698 18300 11704 18352
rect 11756 18340 11762 18352
rect 13449 18343 13507 18349
rect 13449 18340 13461 18343
rect 11756 18312 13461 18340
rect 11756 18300 11762 18312
rect 13449 18309 13461 18312
rect 13495 18309 13507 18343
rect 13449 18303 13507 18309
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 9769 18275 9827 18281
rect 9769 18272 9781 18275
rect 9456 18244 9781 18272
rect 9456 18232 9462 18244
rect 9769 18241 9781 18244
rect 9815 18241 9827 18275
rect 11514 18272 11520 18284
rect 11475 18244 11520 18272
rect 9769 18235 9827 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 12986 18232 12992 18244
rect 13044 18272 13050 18284
rect 13814 18272 13820 18284
rect 13044 18244 13820 18272
rect 13044 18232 13050 18244
rect 13814 18232 13820 18244
rect 13872 18272 13878 18284
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13872 18244 14013 18272
rect 13872 18232 13878 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 14001 18235 14059 18241
rect 8619 18176 9352 18204
rect 9677 18207 9735 18213
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 10686 18204 10692 18216
rect 9723 18176 10692 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12805 18207 12863 18213
rect 11931 18176 12296 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 5537 18139 5595 18145
rect 5537 18105 5549 18139
rect 5583 18136 5595 18139
rect 6638 18136 6644 18148
rect 5583 18108 6644 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 8294 18136 8300 18148
rect 6748 18108 8300 18136
rect 4890 18068 4896 18080
rect 3712 18040 4896 18068
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 6748 18068 6776 18108
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 8665 18139 8723 18145
rect 8665 18105 8677 18139
rect 8711 18136 8723 18139
rect 10226 18136 10232 18148
rect 8711 18108 10232 18136
rect 8711 18105 8723 18108
rect 8665 18099 8723 18105
rect 10226 18096 10232 18108
rect 10284 18096 10290 18148
rect 11333 18139 11391 18145
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 12268 18136 12296 18176
rect 12805 18173 12817 18207
rect 12851 18204 12863 18207
rect 13170 18204 13176 18216
rect 12851 18176 13176 18204
rect 12851 18173 12863 18176
rect 12805 18167 12863 18173
rect 13170 18164 13176 18176
rect 13228 18204 13234 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 13228 18176 14473 18204
rect 13228 18164 13234 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 14461 18167 14519 18173
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 11379 18108 12020 18136
rect 12268 18108 12664 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 7190 18068 7196 18080
rect 5132 18040 6776 18068
rect 7151 18040 7196 18068
rect 5132 18028 5138 18040
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7742 18028 7748 18080
rect 7800 18068 7806 18080
rect 8754 18068 8760 18080
rect 7800 18040 8760 18068
rect 7800 18028 7806 18040
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 9585 18071 9643 18077
rect 9585 18068 9597 18071
rect 9272 18040 9597 18068
rect 9272 18028 9278 18040
rect 9585 18037 9597 18040
rect 9631 18037 9643 18071
rect 9585 18031 9643 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 10836 18040 11253 18068
rect 10836 18028 10842 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 11992 18068 12020 18108
rect 12342 18068 12348 18080
rect 11992 18040 12348 18068
rect 11241 18031 11299 18037
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 12437 18071 12495 18077
rect 12437 18037 12449 18071
rect 12483 18068 12495 18071
rect 12526 18068 12532 18080
rect 12483 18040 12532 18068
rect 12483 18037 12495 18040
rect 12437 18031 12495 18037
rect 12526 18028 12532 18040
rect 12584 18028 12590 18080
rect 12636 18068 12664 18108
rect 12789 18108 13829 18136
rect 12789 18068 12817 18108
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 13817 18099 13875 18105
rect 12636 18040 12817 18068
rect 12894 18028 12900 18080
rect 12952 18068 12958 18080
rect 13722 18068 13728 18080
rect 12952 18040 13728 18068
rect 12952 18028 12958 18040
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 14090 18068 14096 18080
rect 13955 18040 14096 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 22554 18068 22560 18080
rect 19484 18040 22560 18068
rect 19484 18028 19490 18040
rect 22554 18028 22560 18040
rect 22612 18028 22618 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 3142 17864 3148 17876
rect 3103 17836 3148 17864
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 5905 17867 5963 17873
rect 5905 17864 5917 17867
rect 3568 17836 5917 17864
rect 3568 17824 3574 17836
rect 5905 17833 5917 17836
rect 5951 17833 5963 17867
rect 5905 17827 5963 17833
rect 6638 17824 6644 17876
rect 6696 17864 6702 17876
rect 6917 17867 6975 17873
rect 6917 17864 6929 17867
rect 6696 17836 6929 17864
rect 6696 17824 6702 17836
rect 6917 17833 6929 17836
rect 6963 17864 6975 17867
rect 7190 17864 7196 17876
rect 6963 17836 7196 17864
rect 6963 17833 6975 17836
rect 6917 17827 6975 17833
rect 7190 17824 7196 17836
rect 7248 17824 7254 17876
rect 7558 17824 7564 17876
rect 7616 17864 7622 17876
rect 11422 17864 11428 17876
rect 7616 17836 11428 17864
rect 7616 17824 7622 17836
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 12483 17836 12848 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 8570 17796 8576 17808
rect 1504 17768 7328 17796
rect 1504 17737 1532 17768
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17697 1547 17731
rect 2222 17728 2228 17740
rect 2183 17700 2228 17728
rect 1489 17691 1547 17697
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 2958 17728 2964 17740
rect 2919 17700 2964 17728
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4154 17728 4160 17740
rect 4111 17700 4160 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 4332 17731 4390 17737
rect 4332 17697 4344 17731
rect 4378 17728 4390 17731
rect 4706 17728 4712 17740
rect 4378 17700 4712 17728
rect 4378 17697 4390 17700
rect 4332 17691 4390 17697
rect 4706 17688 4712 17700
rect 4764 17688 4770 17740
rect 5721 17731 5779 17737
rect 5721 17697 5733 17731
rect 5767 17728 5779 17731
rect 5810 17728 5816 17740
rect 5767 17700 5816 17728
rect 5767 17697 5779 17700
rect 5721 17691 5779 17697
rect 5810 17688 5816 17700
rect 5868 17688 5874 17740
rect 6822 17728 6828 17740
rect 6783 17700 6828 17728
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7300 17728 7328 17768
rect 7576 17768 8576 17796
rect 7576 17728 7604 17768
rect 8570 17756 8576 17768
rect 8628 17756 8634 17808
rect 12820 17805 12848 17836
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 13909 17867 13967 17873
rect 13909 17864 13921 17867
rect 13872 17836 13921 17864
rect 13872 17824 13878 17836
rect 13909 17833 13921 17836
rect 13955 17833 13967 17867
rect 13909 17827 13967 17833
rect 14461 17867 14519 17873
rect 14461 17833 14473 17867
rect 14507 17864 14519 17867
rect 20622 17864 20628 17876
rect 14507 17836 20628 17864
rect 14507 17833 14519 17836
rect 14461 17827 14519 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 12796 17799 12854 17805
rect 8680 17768 11836 17796
rect 7742 17737 7748 17740
rect 7736 17728 7748 17737
rect 7300 17700 7604 17728
rect 7703 17700 7748 17728
rect 7736 17691 7748 17700
rect 7742 17688 7748 17691
rect 7800 17688 7806 17740
rect 1394 17620 1400 17672
rect 1452 17660 1458 17672
rect 1673 17663 1731 17669
rect 1673 17660 1685 17663
rect 1452 17632 1685 17660
rect 1452 17620 1458 17632
rect 1673 17629 1685 17632
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 2501 17663 2559 17669
rect 2501 17629 2513 17663
rect 2547 17660 2559 17663
rect 2547 17632 3280 17660
rect 2547 17629 2559 17632
rect 2501 17623 2559 17629
rect 2590 17484 2596 17536
rect 2648 17524 2654 17536
rect 3142 17524 3148 17536
rect 2648 17496 3148 17524
rect 2648 17484 2654 17496
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 3252 17524 3280 17632
rect 3326 17620 3332 17672
rect 3384 17660 3390 17672
rect 3513 17663 3571 17669
rect 3513 17660 3525 17663
rect 3384 17632 3525 17660
rect 3384 17620 3390 17632
rect 3513 17629 3525 17632
rect 3559 17629 3571 17663
rect 3513 17623 3571 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 7190 17660 7196 17672
rect 7147 17632 7196 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 7282 17620 7288 17672
rect 7340 17660 7346 17672
rect 7469 17663 7527 17669
rect 7469 17660 7481 17663
rect 7340 17632 7481 17660
rect 7340 17620 7346 17632
rect 7469 17629 7481 17632
rect 7515 17629 7527 17663
rect 7469 17623 7527 17629
rect 3694 17552 3700 17604
rect 3752 17592 3758 17604
rect 4062 17592 4068 17604
rect 3752 17564 4068 17592
rect 3752 17552 3758 17564
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 5534 17592 5540 17604
rect 5000 17564 5540 17592
rect 5000 17524 5028 17564
rect 5534 17552 5540 17564
rect 5592 17552 5598 17604
rect 5828 17564 7236 17592
rect 5442 17524 5448 17536
rect 3252 17496 5028 17524
rect 5355 17496 5448 17524
rect 5442 17484 5448 17496
rect 5500 17524 5506 17536
rect 5828 17524 5856 17564
rect 5500 17496 5856 17524
rect 6457 17527 6515 17533
rect 5500 17484 5506 17496
rect 6457 17493 6469 17527
rect 6503 17524 6515 17527
rect 7098 17524 7104 17536
rect 6503 17496 7104 17524
rect 6503 17493 6515 17496
rect 6457 17487 6515 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 7208 17524 7236 17564
rect 8680 17524 8708 17768
rect 9125 17731 9183 17737
rect 9125 17697 9137 17731
rect 9171 17728 9183 17731
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9171 17700 10057 17728
rect 9171 17697 9183 17700
rect 9125 17691 9183 17697
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10873 17731 10931 17737
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 10962 17728 10968 17740
rect 10919 17700 10968 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11140 17731 11198 17737
rect 11140 17697 11152 17731
rect 11186 17728 11198 17731
rect 11698 17728 11704 17740
rect 11186 17700 11704 17728
rect 11186 17697 11198 17700
rect 11140 17691 11198 17697
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11808 17728 11836 17768
rect 12796 17765 12808 17799
rect 12842 17765 12854 17799
rect 12796 17759 12854 17765
rect 11808 17700 14228 17728
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 8996 17632 10149 17660
rect 8996 17620 9002 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10502 17660 10508 17672
rect 10367 17632 10508 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 8849 17595 8907 17601
rect 8849 17561 8861 17595
rect 8895 17592 8907 17595
rect 9766 17592 9772 17604
rect 8895 17564 9772 17592
rect 8895 17561 8907 17564
rect 8849 17555 8907 17561
rect 9766 17552 9772 17564
rect 9824 17592 9830 17604
rect 10336 17592 10364 17623
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 12526 17660 12532 17672
rect 12487 17632 12532 17660
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 14200 17660 14228 17700
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14332 17700 14377 17728
rect 14332 17688 14338 17700
rect 18506 17660 18512 17672
rect 14200 17632 18512 17660
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 9824 17564 10364 17592
rect 9824 17552 9830 17564
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 12253 17595 12311 17601
rect 12253 17592 12265 17595
rect 12216 17564 12265 17592
rect 12216 17552 12222 17564
rect 12253 17561 12265 17564
rect 12299 17592 12311 17595
rect 12437 17595 12495 17601
rect 12437 17592 12449 17595
rect 12299 17564 12449 17592
rect 12299 17561 12311 17564
rect 12253 17555 12311 17561
rect 12437 17561 12449 17564
rect 12483 17561 12495 17595
rect 12437 17555 12495 17561
rect 9674 17524 9680 17536
rect 7208 17496 8708 17524
rect 9635 17496 9680 17524
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 13814 17524 13820 17536
rect 9916 17496 13820 17524
rect 9916 17484 9922 17496
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 4617 17323 4675 17329
rect 2148 17292 4568 17320
rect 1578 17116 1584 17128
rect 1539 17088 1584 17116
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 2148 17125 2176 17292
rect 2682 17212 2688 17264
rect 2740 17252 2746 17264
rect 4540 17252 4568 17292
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 4706 17320 4712 17332
rect 4663 17292 4712 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 6178 17320 6184 17332
rect 5592 17292 6184 17320
rect 5592 17280 5598 17292
rect 6178 17280 6184 17292
rect 6236 17280 6242 17332
rect 9858 17320 9864 17332
rect 6840 17292 9864 17320
rect 6730 17252 6736 17264
rect 2740 17224 3280 17252
rect 4540 17224 6736 17252
rect 2740 17212 2746 17224
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 2958 17184 2964 17196
rect 2455 17156 2964 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 2958 17144 2964 17156
rect 3016 17144 3022 17196
rect 3252 17125 3280 17224
rect 6730 17212 6736 17224
rect 6788 17212 6794 17264
rect 4709 17187 4767 17193
rect 4709 17153 4721 17187
rect 4755 17184 4767 17187
rect 5445 17187 5503 17193
rect 5445 17184 5457 17187
rect 4755 17156 5457 17184
rect 4755 17153 4767 17156
rect 4709 17147 4767 17153
rect 5445 17153 5457 17156
rect 5491 17153 5503 17187
rect 6840 17184 6868 17292
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10962 17320 10968 17332
rect 10336 17292 10968 17320
rect 10042 17252 10048 17264
rect 10003 17224 10048 17252
rect 10042 17212 10048 17224
rect 10100 17252 10106 17264
rect 10229 17255 10287 17261
rect 10229 17252 10241 17255
rect 10100 17224 10241 17252
rect 10100 17212 10106 17224
rect 10229 17221 10241 17224
rect 10275 17221 10287 17255
rect 10229 17215 10287 17221
rect 10336 17193 10364 17292
rect 10962 17280 10968 17292
rect 11020 17320 11026 17332
rect 11698 17320 11704 17332
rect 11020 17292 11284 17320
rect 11659 17292 11704 17320
rect 11020 17280 11026 17292
rect 11256 17252 11284 17292
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 11940 17292 11989 17320
rect 11940 17280 11946 17292
rect 11977 17289 11989 17292
rect 12023 17289 12035 17323
rect 11977 17283 12035 17289
rect 11992 17252 12020 17283
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 13633 17323 13691 17329
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 13633 17289 13645 17323
rect 13679 17320 13691 17323
rect 13906 17320 13912 17332
rect 13679 17292 13912 17320
rect 13679 17289 13691 17292
rect 13633 17283 13691 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 19334 17320 19340 17332
rect 14231 17292 19340 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 19334 17280 19340 17292
rect 19392 17280 19398 17332
rect 12618 17252 12624 17264
rect 11256 17224 12624 17252
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 5445 17147 5503 17153
rect 5552 17156 6868 17184
rect 10321 17187 10379 17193
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17116 3295 17119
rect 3283 17088 4200 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 4172 17060 4200 17088
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 5353 17119 5411 17125
rect 5353 17116 5365 17119
rect 4304 17088 5365 17116
rect 4304 17076 4310 17088
rect 5353 17085 5365 17088
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 3504 17051 3562 17057
rect 3504 17017 3516 17051
rect 3550 17048 3562 17051
rect 3602 17048 3608 17060
rect 3550 17020 3608 17048
rect 3550 17017 3562 17020
rect 3504 17011 3562 17017
rect 3602 17008 3608 17020
rect 3660 17008 3666 17060
rect 4154 17008 4160 17060
rect 4212 17008 4218 17060
rect 5552 17048 5580 17156
rect 10321 17153 10333 17187
rect 10367 17153 10379 17187
rect 10321 17147 10379 17153
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 4724 17020 5580 17048
rect 1670 16940 1676 16992
rect 1728 16980 1734 16992
rect 4724 16980 4752 17020
rect 4890 16980 4896 16992
rect 1728 16952 4752 16980
rect 4851 16952 4896 16980
rect 1728 16940 1734 16952
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 5920 16980 5948 17079
rect 6362 17076 6368 17128
rect 6420 17116 6426 17128
rect 6641 17119 6699 17125
rect 6641 17116 6653 17119
rect 6420 17088 6653 17116
rect 6420 17076 6426 17088
rect 6641 17085 6653 17088
rect 6687 17085 6699 17119
rect 6641 17079 6699 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17085 8723 17119
rect 8665 17079 8723 17085
rect 8932 17119 8990 17125
rect 8932 17085 8944 17119
rect 8978 17116 8990 17119
rect 9766 17116 9772 17128
rect 8978 17088 9772 17116
rect 8978 17085 8990 17088
rect 8932 17079 8990 17085
rect 5408 16952 5948 16980
rect 5408 16940 5414 16952
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6089 16983 6147 16989
rect 6089 16980 6101 16983
rect 6052 16952 6101 16980
rect 6052 16940 6058 16952
rect 6089 16949 6101 16952
rect 6135 16949 6147 16983
rect 6089 16943 6147 16949
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 6328 16952 6469 16980
rect 6328 16940 6334 16952
rect 6457 16949 6469 16952
rect 6503 16980 6515 16983
rect 6840 16980 6868 17079
rect 7092 17051 7150 17057
rect 7092 17017 7104 17051
rect 7138 17048 7150 17051
rect 7190 17048 7196 17060
rect 7138 17020 7196 17048
rect 7138 17017 7150 17020
rect 7092 17011 7150 17017
rect 7190 17008 7196 17020
rect 7248 17048 7254 17060
rect 7650 17048 7656 17060
rect 7248 17020 7656 17048
rect 7248 17008 7254 17020
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 8680 17048 8708 17079
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 10336 17116 10364 17147
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 11756 17156 13001 17184
rect 11756 17144 11762 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 14274 17184 14280 17196
rect 12989 17147 13047 17153
rect 13096 17156 14280 17184
rect 11790 17116 11796 17128
rect 9876 17088 10364 17116
rect 10888 17088 11796 17116
rect 9876 17060 9904 17088
rect 9858 17048 9864 17060
rect 8680 17020 9864 17048
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 10229 17051 10287 17057
rect 10229 17017 10241 17051
rect 10275 17048 10287 17051
rect 10566 17051 10624 17057
rect 10566 17048 10578 17051
rect 10275 17020 10578 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 10566 17017 10578 17020
rect 10612 17017 10624 17051
rect 10566 17011 10624 17017
rect 7282 16980 7288 16992
rect 6503 16952 7288 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7742 16980 7748 16992
rect 7432 16952 7748 16980
rect 7432 16940 7438 16952
rect 7742 16940 7748 16952
rect 7800 16980 7806 16992
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7800 16952 8217 16980
rect 7800 16940 7806 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 8205 16943 8263 16949
rect 8478 16940 8484 16992
rect 8536 16980 8542 16992
rect 10888 16980 10916 17088
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12158 17116 12164 17128
rect 12119 17088 12164 17116
rect 12158 17076 12164 17088
rect 12216 17076 12222 17128
rect 13096 17116 13124 17156
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 13446 17116 13452 17128
rect 12728 17088 13124 17116
rect 13407 17088 13452 17116
rect 11146 17008 11152 17060
rect 11204 17048 11210 17060
rect 12728 17048 12756 17088
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 14016 17048 14044 17079
rect 11204 17020 12756 17048
rect 12820 17020 14044 17048
rect 11204 17008 11210 17020
rect 12820 16992 12848 17020
rect 8536 16952 10916 16980
rect 8536 16940 8542 16952
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11238 16980 11244 16992
rect 11020 16952 11244 16980
rect 11020 16940 11026 16952
rect 11238 16940 11244 16952
rect 11296 16980 11302 16992
rect 11882 16980 11888 16992
rect 11296 16952 11888 16980
rect 11296 16940 11302 16952
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 12986 16980 12992 16992
rect 12943 16952 12992 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2280 16748 2973 16776
rect 2280 16736 2286 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 3326 16776 3332 16788
rect 3287 16748 3332 16776
rect 2961 16739 3019 16745
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 3421 16779 3479 16785
rect 3421 16745 3433 16779
rect 3467 16776 3479 16779
rect 4890 16776 4896 16788
rect 3467 16748 4896 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 5997 16779 6055 16785
rect 5997 16776 6009 16779
rect 5408 16748 6009 16776
rect 5408 16736 5414 16748
rect 5997 16745 6009 16748
rect 6043 16745 6055 16779
rect 5997 16739 6055 16745
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 2501 16711 2559 16717
rect 2501 16708 2513 16711
rect 1636 16680 2513 16708
rect 1636 16668 1642 16680
rect 2501 16677 2513 16680
rect 2547 16677 2559 16711
rect 5074 16708 5080 16720
rect 2501 16671 2559 16677
rect 3344 16680 5080 16708
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 2225 16643 2283 16649
rect 2225 16609 2237 16643
rect 2271 16640 2283 16643
rect 3344 16640 3372 16680
rect 5074 16668 5080 16680
rect 5132 16668 5138 16720
rect 6012 16708 6040 16739
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 6880 16748 9137 16776
rect 6880 16736 6886 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9125 16739 9183 16745
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10134 16736 10140 16788
rect 10192 16736 10198 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10870 16776 10876 16788
rect 10459 16748 10876 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 10965 16779 11023 16785
rect 10965 16745 10977 16779
rect 11011 16776 11023 16779
rect 11238 16776 11244 16788
rect 11011 16748 11244 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 11425 16779 11483 16785
rect 11425 16745 11437 16779
rect 11471 16776 11483 16779
rect 11606 16776 11612 16788
rect 11471 16748 11612 16776
rect 11471 16745 11483 16748
rect 11425 16739 11483 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 6518 16711 6576 16717
rect 6518 16708 6530 16711
rect 6012 16680 6530 16708
rect 6518 16677 6530 16680
rect 6564 16677 6576 16711
rect 8478 16708 8484 16720
rect 8439 16680 8484 16708
rect 6518 16671 6576 16677
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 8573 16711 8631 16717
rect 8573 16677 8585 16711
rect 8619 16708 8631 16711
rect 10152 16708 10180 16736
rect 8619 16680 10180 16708
rect 10321 16711 10379 16717
rect 8619 16677 8631 16680
rect 8573 16671 8631 16677
rect 10321 16677 10333 16711
rect 10367 16708 10379 16711
rect 11146 16708 11152 16720
rect 10367 16680 11152 16708
rect 10367 16677 10379 16680
rect 10321 16671 10379 16677
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 13446 16668 13452 16720
rect 13504 16708 13510 16720
rect 14553 16711 14611 16717
rect 14553 16708 14565 16711
rect 13504 16680 14565 16708
rect 13504 16668 13510 16680
rect 14553 16677 14565 16680
rect 14599 16677 14611 16711
rect 14553 16671 14611 16677
rect 2271 16612 3372 16640
rect 2271 16609 2283 16612
rect 2225 16603 2283 16609
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3476 16612 4077 16640
rect 3476 16600 3482 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4617 16643 4675 16649
rect 4617 16640 4629 16643
rect 4212 16612 4629 16640
rect 4212 16600 4218 16612
rect 4617 16609 4629 16612
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 4884 16643 4942 16649
rect 4884 16609 4896 16643
rect 4930 16640 4942 16643
rect 7558 16640 7564 16652
rect 4930 16612 7564 16640
rect 4930 16609 4942 16612
rect 4884 16603 4942 16609
rect 3602 16572 3608 16584
rect 3563 16544 3608 16572
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 2958 16464 2964 16516
rect 3016 16504 3022 16516
rect 3786 16504 3792 16516
rect 3016 16476 3792 16504
rect 3016 16464 3022 16476
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 4062 16464 4068 16516
rect 4120 16504 4126 16516
rect 4249 16507 4307 16513
rect 4249 16504 4261 16507
rect 4120 16476 4261 16504
rect 4120 16464 4126 16476
rect 4249 16473 4261 16476
rect 4295 16473 4307 16507
rect 4249 16467 4307 16473
rect 566 16396 572 16448
rect 624 16436 630 16448
rect 4154 16436 4160 16448
rect 624 16408 4160 16436
rect 624 16396 630 16408
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 4632 16436 4660 16603
rect 7558 16600 7564 16612
rect 7616 16640 7622 16652
rect 11238 16640 11244 16652
rect 7616 16612 11244 16640
rect 7616 16600 7622 16612
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11379 16612 11989 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 11977 16609 11989 16612
rect 12023 16609 12035 16643
rect 11977 16603 12035 16609
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 12877 16643 12935 16649
rect 12877 16640 12889 16643
rect 12400 16612 12889 16640
rect 12400 16600 12406 16612
rect 12877 16609 12889 16612
rect 12923 16609 12935 16643
rect 14274 16640 14280 16652
rect 14235 16612 14280 16640
rect 12877 16603 12935 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 6270 16572 6276 16584
rect 6231 16544 6276 16572
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 8665 16575 8723 16581
rect 8665 16541 8677 16575
rect 8711 16541 8723 16575
rect 8665 16535 8723 16541
rect 6288 16436 6316 16532
rect 7650 16504 7656 16516
rect 7563 16476 7656 16504
rect 7650 16464 7656 16476
rect 7708 16504 7714 16516
rect 8680 16504 8708 16535
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 10502 16572 10508 16584
rect 9272 16544 10364 16572
rect 10463 16544 10508 16572
rect 9272 16532 9278 16544
rect 7708 16476 8708 16504
rect 7708 16464 7714 16476
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10134 16504 10140 16516
rect 9640 16476 10140 16504
rect 9640 16464 9646 16476
rect 10134 16464 10140 16476
rect 10192 16464 10198 16516
rect 10336 16504 10364 16544
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11698 16572 11704 16584
rect 11655 16544 11704 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 12618 16572 12624 16584
rect 12579 16544 12624 16572
rect 12618 16532 12624 16544
rect 12676 16532 12682 16584
rect 11790 16504 11796 16516
rect 10336 16476 11796 16504
rect 11790 16464 11796 16476
rect 11848 16464 11854 16516
rect 13630 16464 13636 16516
rect 13688 16504 13694 16516
rect 14001 16507 14059 16513
rect 14001 16504 14013 16507
rect 13688 16476 14013 16504
rect 13688 16464 13694 16476
rect 14001 16473 14013 16476
rect 14047 16473 14059 16507
rect 14001 16467 14059 16473
rect 4632 16408 6316 16436
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 8113 16439 8171 16445
rect 8113 16436 8125 16439
rect 7800 16408 8125 16436
rect 7800 16396 7806 16408
rect 8113 16405 8125 16408
rect 8159 16405 8171 16439
rect 8113 16399 8171 16405
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 9122 16436 9128 16448
rect 8260 16408 9128 16436
rect 8260 16396 8266 16408
rect 9122 16396 9128 16408
rect 9180 16436 9186 16448
rect 12250 16436 12256 16448
rect 9180 16408 12256 16436
rect 9180 16396 9186 16408
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 6822 16232 6828 16244
rect 3007 16204 6828 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 8202 16232 8208 16244
rect 7248 16204 8208 16232
rect 7248 16192 7254 16204
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8352 16204 9045 16232
rect 8352 16192 8358 16204
rect 9033 16201 9045 16204
rect 9079 16201 9091 16235
rect 9033 16195 9091 16201
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 14274 16232 14280 16244
rect 10091 16204 14280 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 14274 16192 14280 16204
rect 14332 16192 14338 16244
rect 1026 16124 1032 16176
rect 1084 16164 1090 16176
rect 3418 16164 3424 16176
rect 1084 16136 3424 16164
rect 1084 16124 1090 16136
rect 3418 16124 3424 16136
rect 3476 16124 3482 16176
rect 3973 16167 4031 16173
rect 3973 16133 3985 16167
rect 4019 16164 4031 16167
rect 4246 16164 4252 16176
rect 4019 16136 4252 16164
rect 4019 16133 4031 16136
rect 3973 16127 4031 16133
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 6365 16167 6423 16173
rect 6365 16164 6377 16167
rect 4816 16136 6377 16164
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16096 2651 16099
rect 3605 16099 3663 16105
rect 3605 16096 3617 16099
rect 2639 16068 3617 16096
rect 2639 16065 2651 16068
rect 2593 16059 2651 16065
rect 3605 16065 3617 16068
rect 3651 16096 3663 16099
rect 3694 16096 3700 16108
rect 3651 16068 3700 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 3694 16056 3700 16068
rect 3752 16056 3758 16108
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16096 4675 16099
rect 4706 16096 4712 16108
rect 4663 16068 4712 16096
rect 4663 16065 4675 16068
rect 4617 16059 4675 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 16028 2375 16031
rect 2958 16028 2964 16040
rect 2363 16000 2964 16028
rect 2363 15997 2375 16000
rect 2317 15991 2375 15997
rect 2958 15988 2964 16000
rect 3016 15988 3022 16040
rect 3234 15988 3240 16040
rect 3292 16028 3298 16040
rect 4816 16028 4844 16136
rect 6365 16133 6377 16136
rect 6411 16133 6423 16167
rect 11057 16167 11115 16173
rect 11057 16164 11069 16167
rect 6365 16127 6423 16133
rect 8404 16136 11069 16164
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 5859 16068 7481 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 7469 16065 7481 16068
rect 7515 16096 7527 16099
rect 7558 16096 7564 16108
rect 7515 16068 7564 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8404 16105 8432 16136
rect 11057 16133 11069 16136
rect 11103 16133 11115 16167
rect 11057 16127 11115 16133
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 9306 16096 9312 16108
rect 8619 16068 9312 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 9582 16096 9588 16108
rect 9416 16068 9588 16096
rect 3292 16000 4844 16028
rect 5537 16031 5595 16037
rect 3292 15988 3298 16000
rect 5537 15997 5549 16031
rect 5583 15997 5595 16031
rect 6178 16028 6184 16040
rect 6139 16000 6184 16028
rect 5537 15991 5595 15997
rect 1762 15920 1768 15972
rect 1820 15960 1826 15972
rect 2409 15963 2467 15969
rect 1820 15932 2360 15960
rect 1820 15920 1826 15932
rect 1946 15892 1952 15904
rect 1907 15864 1952 15892
rect 1946 15852 1952 15864
rect 2004 15852 2010 15904
rect 2332 15892 2360 15932
rect 2409 15929 2421 15963
rect 2455 15960 2467 15963
rect 2866 15960 2872 15972
rect 2455 15932 2872 15960
rect 2455 15929 2467 15932
rect 2409 15923 2467 15929
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 3418 15960 3424 15972
rect 3379 15932 3424 15960
rect 3418 15920 3424 15932
rect 3476 15960 3482 15972
rect 3970 15960 3976 15972
rect 3476 15932 3976 15960
rect 3476 15920 3482 15932
rect 3970 15920 3976 15932
rect 4028 15920 4034 15972
rect 5552 15960 5580 15991
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 7190 16028 7196 16040
rect 7151 16000 7196 16028
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 9416 16028 9444 16068
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 10042 16096 10048 16108
rect 9723 16068 10048 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 10686 16096 10692 16108
rect 10647 16068 10692 16096
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 11609 16099 11667 16105
rect 11609 16096 11621 16099
rect 10796 16068 11621 16096
rect 7331 16000 9444 16028
rect 9493 16031 9551 16037
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 9493 15997 9505 16031
rect 9539 16028 9551 16031
rect 9950 16028 9956 16040
rect 9539 16000 9956 16028
rect 9539 15997 9551 16000
rect 9493 15991 9551 15997
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10796 16028 10824 16068
rect 11609 16065 11621 16068
rect 11655 16065 11667 16099
rect 11609 16059 11667 16065
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 11848 16068 13001 16096
rect 11848 16056 11854 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13814 16096 13820 16108
rect 13219 16068 13820 16096
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 11422 16028 11428 16040
rect 10284 16000 10824 16028
rect 11383 16000 11428 16028
rect 10284 15988 10290 16000
rect 11422 15988 11428 16000
rect 11480 15988 11486 16040
rect 11698 15988 11704 16040
rect 11756 16028 11762 16040
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 11756 16000 13553 16028
rect 11756 15988 11762 16000
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 13541 15991 13599 15997
rect 6270 15960 6276 15972
rect 5552 15932 6276 15960
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 9401 15963 9459 15969
rect 7944 15932 9260 15960
rect 3329 15895 3387 15901
rect 3329 15892 3341 15895
rect 2332 15864 3341 15892
rect 3329 15861 3341 15864
rect 3375 15892 3387 15895
rect 3602 15892 3608 15904
rect 3375 15864 3608 15892
rect 3375 15861 3387 15864
rect 3329 15855 3387 15861
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 4062 15852 4068 15904
rect 4120 15892 4126 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 4120 15864 4353 15892
rect 4120 15852 4126 15864
rect 4341 15861 4353 15864
rect 4387 15861 4399 15895
rect 4341 15855 4399 15861
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 4890 15892 4896 15904
rect 4479 15864 4896 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4890 15852 4896 15864
rect 4948 15852 4954 15904
rect 5169 15895 5227 15901
rect 5169 15861 5181 15895
rect 5215 15892 5227 15895
rect 5442 15892 5448 15904
rect 5215 15864 5448 15892
rect 5215 15861 5227 15864
rect 5169 15855 5227 15861
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 5902 15892 5908 15904
rect 5675 15864 5908 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 5902 15852 5908 15864
rect 5960 15852 5966 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7944 15901 7972 15932
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15861 7987 15895
rect 8294 15892 8300 15904
rect 8255 15864 8300 15892
rect 7929 15855 7987 15861
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 9232 15892 9260 15932
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 9674 15960 9680 15972
rect 9447 15932 9680 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 10505 15963 10563 15969
rect 10505 15960 10517 15963
rect 9784 15932 10517 15960
rect 9784 15892 9812 15932
rect 10505 15929 10517 15932
rect 10551 15929 10563 15963
rect 10505 15923 10563 15929
rect 13817 15963 13875 15969
rect 13817 15929 13829 15963
rect 13863 15960 13875 15963
rect 13906 15960 13912 15972
rect 13863 15932 13912 15960
rect 13863 15929 13875 15932
rect 13817 15923 13875 15929
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 9232 15864 9812 15892
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 9916 15864 10425 15892
rect 9916 15852 9922 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 10778 15852 10784 15904
rect 10836 15892 10842 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 10836 15864 11529 15892
rect 10836 15852 10842 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12032 15864 12541 15892
rect 12032 15852 12038 15864
rect 12529 15861 12541 15864
rect 12575 15861 12587 15895
rect 12894 15892 12900 15904
rect 12855 15864 12900 15892
rect 12529 15855 12587 15861
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2317 15691 2375 15697
rect 2317 15688 2329 15691
rect 2004 15660 2329 15688
rect 2004 15648 2010 15660
rect 2317 15657 2329 15660
rect 2363 15657 2375 15691
rect 3881 15691 3939 15697
rect 3881 15688 3893 15691
rect 2317 15651 2375 15657
rect 2608 15660 3893 15688
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1670 15552 1676 15564
rect 1443 15524 1676 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1670 15512 1676 15524
rect 1728 15512 1734 15564
rect 2406 15552 2412 15564
rect 2367 15524 2412 15552
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2608 15493 2636 15660
rect 3881 15657 3893 15660
rect 3927 15657 3939 15691
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 3881 15651 3939 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4522 15688 4528 15700
rect 4483 15660 4528 15688
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 5074 15688 5080 15700
rect 5035 15660 5080 15688
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5537 15691 5595 15697
rect 5537 15657 5549 15691
rect 5583 15688 5595 15691
rect 5905 15691 5963 15697
rect 5905 15688 5917 15691
rect 5583 15660 5917 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 5905 15657 5917 15660
rect 5951 15657 5963 15691
rect 5905 15651 5963 15657
rect 6089 15691 6147 15697
rect 6089 15657 6101 15691
rect 6135 15688 6147 15691
rect 6270 15688 6276 15700
rect 6135 15660 6276 15688
rect 6135 15657 6147 15660
rect 6089 15651 6147 15657
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 6730 15688 6736 15700
rect 6691 15660 6736 15688
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 7098 15688 7104 15700
rect 7059 15660 7104 15688
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 7193 15691 7251 15697
rect 7193 15657 7205 15691
rect 7239 15688 7251 15691
rect 7742 15688 7748 15700
rect 7239 15660 7748 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 9306 15688 9312 15700
rect 9267 15660 9312 15688
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 10686 15648 10692 15700
rect 10744 15688 10750 15700
rect 11057 15691 11115 15697
rect 11057 15688 11069 15691
rect 10744 15660 11069 15688
rect 10744 15648 10750 15660
rect 11057 15657 11069 15660
rect 11103 15657 11115 15691
rect 11057 15651 11115 15657
rect 11609 15691 11667 15697
rect 11609 15657 11621 15691
rect 11655 15688 11667 15691
rect 11698 15688 11704 15700
rect 11655 15660 11704 15688
rect 11655 15657 11667 15660
rect 11609 15651 11667 15657
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 11974 15688 11980 15700
rect 11935 15660 11980 15688
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 12952 15660 14289 15688
rect 12952 15648 12958 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 8294 15620 8300 15632
rect 2884 15592 8300 15620
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 1949 15351 2007 15357
rect 1949 15317 1961 15351
rect 1995 15348 2007 15351
rect 2884 15348 2912 15592
rect 8294 15580 8300 15592
rect 8352 15580 8358 15632
rect 9324 15620 9352 15648
rect 9922 15623 9980 15629
rect 9922 15620 9934 15623
rect 9324 15592 9934 15620
rect 9922 15589 9934 15592
rect 9968 15589 9980 15623
rect 9922 15583 9980 15589
rect 10410 15580 10416 15632
rect 10468 15620 10474 15632
rect 13262 15620 13268 15632
rect 10468 15592 13268 15620
rect 10468 15580 10474 15592
rect 13262 15580 13268 15592
rect 13320 15580 13326 15632
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 3375 15524 3801 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 4430 15552 4436 15564
rect 4391 15524 4436 15552
rect 3789 15515 3847 15521
rect 4430 15512 4436 15524
rect 4488 15512 4494 15564
rect 8202 15561 8208 15564
rect 8185 15555 8208 15561
rect 8185 15552 8197 15555
rect 4632 15524 8197 15552
rect 3142 15444 3148 15496
rect 3200 15484 3206 15496
rect 3421 15487 3479 15493
rect 3421 15484 3433 15487
rect 3200 15456 3433 15484
rect 3200 15444 3206 15456
rect 3421 15453 3433 15456
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 3694 15484 3700 15496
rect 3651 15456 3700 15484
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 3881 15487 3939 15493
rect 3881 15453 3893 15487
rect 3927 15484 3939 15487
rect 4632 15484 4660 15524
rect 8185 15521 8197 15524
rect 8260 15552 8266 15564
rect 9674 15552 9680 15564
rect 8260 15524 8333 15552
rect 9635 15524 9680 15552
rect 8185 15515 8208 15521
rect 8202 15512 8208 15515
rect 8260 15512 8266 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 12710 15552 12716 15564
rect 12115 15524 12716 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 12888 15555 12946 15561
rect 12888 15521 12900 15555
rect 12934 15552 12946 15555
rect 13814 15552 13820 15564
rect 12934 15524 13820 15552
rect 12934 15521 12946 15524
rect 12888 15515 12946 15521
rect 13814 15512 13820 15524
rect 13872 15552 13878 15564
rect 14550 15552 14556 15564
rect 13872 15524 14556 15552
rect 13872 15512 13878 15524
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 3927 15456 4660 15484
rect 4709 15487 4767 15493
rect 3927 15453 3939 15456
rect 3881 15447 3939 15453
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 4890 15484 4896 15496
rect 4755 15456 4896 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 5629 15487 5687 15493
rect 5629 15484 5641 15487
rect 5408 15456 5641 15484
rect 5408 15444 5414 15456
rect 5629 15453 5641 15456
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 5905 15487 5963 15493
rect 5905 15453 5917 15487
rect 5951 15484 5963 15487
rect 6822 15484 6828 15496
rect 5951 15456 6828 15484
rect 5951 15453 5963 15456
rect 5905 15447 5963 15453
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 7374 15484 7380 15496
rect 7335 15456 7380 15484
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15453 12311 15487
rect 12618 15484 12624 15496
rect 12579 15456 12624 15484
rect 12253 15447 12311 15453
rect 2961 15419 3019 15425
rect 2961 15385 2973 15419
rect 3007 15416 3019 15419
rect 3007 15388 7236 15416
rect 3007 15385 3019 15388
rect 2961 15379 3019 15385
rect 1995 15320 2912 15348
rect 3789 15351 3847 15357
rect 1995 15317 2007 15320
rect 1949 15311 2007 15317
rect 3789 15317 3801 15351
rect 3835 15348 3847 15351
rect 4154 15348 4160 15360
rect 3835 15320 4160 15348
rect 3835 15317 3847 15320
rect 3789 15311 3847 15317
rect 4154 15308 4160 15320
rect 4212 15348 4218 15360
rect 5442 15348 5448 15360
rect 4212 15320 5448 15348
rect 4212 15308 4218 15320
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 7208 15348 7236 15388
rect 7282 15376 7288 15428
rect 7340 15416 7346 15428
rect 7944 15416 7972 15447
rect 12268 15416 12296 15447
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 12342 15416 12348 15428
rect 7340 15388 7972 15416
rect 12255 15388 12348 15416
rect 7340 15376 7346 15388
rect 12342 15376 12348 15388
rect 12400 15416 12406 15428
rect 12400 15388 12664 15416
rect 12400 15376 12406 15388
rect 10778 15348 10784 15360
rect 7208 15320 10784 15348
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 12636 15348 12664 15388
rect 14001 15351 14059 15357
rect 14001 15348 14013 15351
rect 12636 15320 14013 15348
rect 14001 15317 14013 15320
rect 14047 15317 14059 15351
rect 14001 15311 14059 15317
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 3418 15144 3424 15156
rect 3379 15116 3424 15144
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 5074 15144 5080 15156
rect 3896 15116 5080 15144
rect 3896 15076 3924 15116
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 5718 15144 5724 15156
rect 5679 15116 5724 15144
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 6362 15104 6368 15156
rect 6420 15144 6426 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 6420 15116 8493 15144
rect 6420 15104 6426 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 8481 15107 8539 15113
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 9858 15144 9864 15156
rect 9171 15116 9864 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 14001 15147 14059 15153
rect 14001 15144 14013 15147
rect 12768 15116 14013 15144
rect 12768 15104 12774 15116
rect 14001 15113 14013 15116
rect 14047 15113 14059 15147
rect 15010 15144 15016 15156
rect 14971 15116 15016 15144
rect 14001 15107 14059 15113
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 1504 15048 3924 15076
rect 1504 14949 1532 15048
rect 5258 15036 5264 15088
rect 5316 15076 5322 15088
rect 5445 15079 5503 15085
rect 5445 15076 5457 15079
rect 5316 15048 5457 15076
rect 5316 15036 5322 15048
rect 5445 15045 5457 15048
rect 5491 15045 5503 15079
rect 8202 15076 8208 15088
rect 8163 15048 8208 15076
rect 5445 15039 5503 15045
rect 8202 15036 8208 15048
rect 8260 15076 8266 15088
rect 8260 15048 9260 15076
rect 8260 15036 8266 15048
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 1762 14968 1768 15020
rect 1820 15008 1826 15020
rect 2869 15011 2927 15017
rect 1820 14980 2636 15008
rect 1820 14968 1826 14980
rect 2608 14949 2636 14980
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3050 15008 3056 15020
rect 2915 14980 3056 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 3970 14968 3976 15020
rect 4028 15008 4034 15020
rect 6365 15011 6423 15017
rect 4028 14980 4200 15008
rect 4028 14968 4034 14980
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 3234 14940 3240 14952
rect 3195 14912 3240 14940
rect 2593 14903 2651 14909
rect 3234 14900 3240 14912
rect 3292 14900 3298 14952
rect 3694 14900 3700 14952
rect 3752 14940 3758 14952
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3752 14912 4077 14940
rect 3752 14900 3758 14912
rect 4065 14909 4077 14912
rect 4111 14909 4123 14943
rect 4172 14940 4200 14980
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 6411 14980 6960 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6089 14943 6147 14949
rect 6089 14940 6101 14943
rect 4172 14912 6101 14940
rect 4065 14903 4123 14909
rect 6089 14909 6101 14912
rect 6135 14940 6147 14943
rect 6270 14940 6276 14952
rect 6135 14912 6276 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6270 14900 6276 14912
rect 6328 14900 6334 14952
rect 4154 14872 4160 14884
rect 2240 14844 4160 14872
rect 2240 14813 2268 14844
rect 4154 14832 4160 14844
rect 4212 14832 4218 14884
rect 4332 14875 4390 14881
rect 4332 14841 4344 14875
rect 4378 14872 4390 14875
rect 4890 14872 4896 14884
rect 4378 14844 4896 14872
rect 4378 14841 4390 14844
rect 4332 14835 4390 14841
rect 4890 14832 4896 14844
rect 4948 14872 4954 14884
rect 6380 14872 6408 14971
rect 6730 14900 6736 14952
rect 6788 14940 6794 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6788 14912 6837 14940
rect 6788 14900 6794 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6932 14940 6960 14980
rect 8202 14940 8208 14952
rect 6932 14912 8208 14940
rect 6825 14903 6883 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8662 14940 8668 14952
rect 8623 14912 8668 14940
rect 8662 14900 8668 14912
rect 8720 14900 8726 14952
rect 9232 14940 9260 15048
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 9950 15076 9956 15088
rect 9640 15048 9956 15076
rect 9640 15036 9646 15048
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 11664 15048 15516 15076
rect 11664 15036 11670 15048
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9364 14980 9689 15008
rect 9364 14968 9370 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 10321 15011 10379 15017
rect 10321 15008 10333 15011
rect 9824 14980 10333 15008
rect 9824 14968 9830 14980
rect 10321 14977 10333 14980
rect 10367 14977 10379 15011
rect 13078 15008 13084 15020
rect 10321 14971 10379 14977
rect 11348 14980 13084 15008
rect 10226 14940 10232 14952
rect 9232 14912 10232 14940
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 11348 14940 11376 14980
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13262 15008 13268 15020
rect 13223 14980 13268 15008
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 13814 15008 13820 15020
rect 13495 14980 13820 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14550 15008 14556 15020
rect 14511 14980 14556 15008
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 15488 15017 15516 15048
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 15008 15715 15011
rect 15930 15008 15936 15020
rect 15703 14980 15936 15008
rect 15703 14977 15715 14980
rect 15657 14971 15715 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 12250 14940 12256 14952
rect 10336 14912 11376 14940
rect 11440 14912 12256 14940
rect 4948 14844 6408 14872
rect 7092 14875 7150 14881
rect 4948 14832 4954 14844
rect 7092 14841 7104 14875
rect 7138 14872 7150 14875
rect 7282 14872 7288 14884
rect 7138 14844 7288 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7282 14832 7288 14844
rect 7340 14832 7346 14884
rect 7374 14832 7380 14884
rect 7432 14872 7438 14884
rect 10336 14872 10364 14912
rect 7432 14844 10364 14872
rect 10588 14875 10646 14881
rect 7432 14832 7438 14844
rect 10588 14841 10600 14875
rect 10634 14872 10646 14875
rect 10686 14872 10692 14884
rect 10634 14844 10692 14872
rect 10634 14841 10646 14844
rect 10588 14835 10646 14841
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 2225 14807 2283 14813
rect 2225 14773 2237 14807
rect 2271 14773 2283 14807
rect 2682 14804 2688 14816
rect 2643 14776 2688 14804
rect 2225 14767 2283 14773
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 3200 14776 6193 14804
rect 3200 14764 3206 14776
rect 6181 14773 6193 14776
rect 6227 14804 6239 14807
rect 8478 14804 8484 14816
rect 6227 14776 8484 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9493 14807 9551 14813
rect 9493 14804 9505 14807
rect 9364 14776 9505 14804
rect 9364 14764 9370 14776
rect 9493 14773 9505 14776
rect 9539 14773 9551 14807
rect 9493 14767 9551 14773
rect 9585 14807 9643 14813
rect 9585 14773 9597 14807
rect 9631 14804 9643 14807
rect 9674 14804 9680 14816
rect 9631 14776 9680 14804
rect 9631 14773 9643 14776
rect 9585 14767 9643 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 11440 14804 11468 14912
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 13280 14940 13308 14968
rect 13630 14940 13636 14952
rect 13280 14912 13636 14940
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 14366 14940 14372 14952
rect 13955 14912 14372 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 14461 14875 14519 14881
rect 14461 14872 14473 14875
rect 12820 14844 14473 14872
rect 11698 14804 11704 14816
rect 9824 14776 11468 14804
rect 11659 14776 11704 14804
rect 9824 14764 9830 14776
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 12820 14813 12848 14844
rect 14461 14841 14473 14844
rect 14507 14841 14519 14875
rect 15378 14872 15384 14884
rect 15339 14844 15384 14872
rect 14461 14835 14519 14841
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 12805 14807 12863 14813
rect 12805 14773 12817 14807
rect 12851 14773 12863 14807
rect 12805 14767 12863 14773
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 13173 14807 13231 14813
rect 13173 14804 13185 14807
rect 12952 14776 13185 14804
rect 12952 14764 12958 14776
rect 13173 14773 13185 14776
rect 13219 14804 13231 14807
rect 18598 14804 18604 14816
rect 13219 14776 18604 14804
rect 13219 14773 13231 14776
rect 13173 14767 13231 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 4479 14572 5089 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 5077 14563 5135 14569
rect 5537 14603 5595 14609
rect 5537 14569 5549 14603
rect 5583 14600 5595 14603
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 5583 14572 8217 14600
rect 5583 14569 5595 14572
rect 5537 14563 5595 14569
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 8205 14563 8263 14569
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 9950 14560 9956 14612
rect 10008 14600 10014 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 10008 14572 10057 14600
rect 10008 14560 10014 14572
rect 10045 14569 10057 14572
rect 10091 14569 10103 14603
rect 10045 14563 10103 14569
rect 10137 14603 10195 14609
rect 10137 14569 10149 14603
rect 10183 14600 10195 14603
rect 15289 14603 15347 14609
rect 15289 14600 15301 14603
rect 10183 14572 15301 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 15289 14569 15301 14572
rect 15335 14569 15347 14603
rect 15289 14563 15347 14569
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 15657 14603 15715 14609
rect 15657 14600 15669 14603
rect 15528 14572 15669 14600
rect 15528 14560 15534 14572
rect 15657 14569 15669 14572
rect 15703 14569 15715 14603
rect 15657 14563 15715 14569
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 19426 14600 19432 14612
rect 15795 14572 19432 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 4246 14492 4252 14544
rect 4304 14532 4310 14544
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 4304 14504 4537 14532
rect 4304 14492 4310 14504
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 5445 14535 5503 14541
rect 5445 14501 5457 14535
rect 5491 14532 5503 14535
rect 5902 14532 5908 14544
rect 5491 14504 5908 14532
rect 5491 14501 5503 14504
rect 5445 14495 5503 14501
rect 5902 14492 5908 14504
rect 5960 14492 5966 14544
rect 5994 14492 6000 14544
rect 6052 14532 6058 14544
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 6052 14504 6469 14532
rect 6052 14492 6058 14504
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 6457 14495 6515 14501
rect 7374 14492 7380 14544
rect 7432 14492 7438 14544
rect 8665 14535 8723 14541
rect 8665 14501 8677 14535
rect 8711 14532 8723 14535
rect 10962 14532 10968 14544
rect 8711 14504 10968 14532
rect 8711 14501 8723 14504
rect 8665 14495 8723 14501
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 11416 14535 11474 14541
rect 11416 14501 11428 14535
rect 11462 14532 11474 14535
rect 11698 14532 11704 14544
rect 11462 14504 11704 14532
rect 11462 14501 11474 14504
rect 11416 14495 11474 14501
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 13596 14504 13952 14532
rect 13596 14492 13602 14504
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2130 14424 2136 14476
rect 2188 14464 2194 14476
rect 2297 14467 2355 14473
rect 2297 14464 2309 14467
rect 2188 14436 2309 14464
rect 2188 14424 2194 14436
rect 2297 14433 2309 14436
rect 2343 14464 2355 14467
rect 4706 14464 4712 14476
rect 2343 14436 4712 14464
rect 2343 14433 2355 14436
rect 2297 14427 2355 14433
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 6270 14424 6276 14476
rect 6328 14464 6334 14476
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 6328 14436 6561 14464
rect 6328 14424 6334 14436
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 2038 14396 2044 14408
rect 1999 14368 2044 14396
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 3436 14368 4629 14396
rect 3050 14288 3056 14340
rect 3108 14328 3114 14340
rect 3436 14337 3464 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4724 14396 4752 14424
rect 5350 14396 5356 14408
rect 4724 14368 5356 14396
rect 4617 14359 4675 14365
rect 5350 14356 5356 14368
rect 5408 14396 5414 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5408 14368 5641 14396
rect 5408 14356 5414 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 6638 14396 6644 14408
rect 6599 14368 6644 14396
rect 5629 14359 5687 14365
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 3108 14300 3433 14328
rect 3108 14288 3114 14300
rect 3421 14297 3433 14300
rect 3467 14297 3479 14331
rect 3421 14291 3479 14297
rect 7193 14331 7251 14337
rect 7193 14297 7205 14331
rect 7239 14328 7251 14331
rect 7392 14328 7420 14492
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 7834 14464 7840 14476
rect 7607 14436 7840 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8573 14467 8631 14473
rect 8573 14464 8585 14467
rect 8352 14436 8585 14464
rect 8352 14424 8358 14436
rect 8573 14433 8585 14436
rect 8619 14464 8631 14467
rect 9766 14464 9772 14476
rect 8619 14436 9772 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 9766 14424 9772 14436
rect 9824 14424 9830 14476
rect 10870 14464 10876 14476
rect 9876 14436 10364 14464
rect 10831 14436 10876 14464
rect 7650 14396 7656 14408
rect 7611 14368 7656 14396
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 7800 14368 7845 14396
rect 7800 14356 7806 14368
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 8849 14399 8907 14405
rect 8849 14396 8861 14399
rect 8260 14368 8861 14396
rect 8260 14356 8266 14368
rect 8849 14365 8861 14368
rect 8895 14396 8907 14399
rect 9398 14396 9404 14408
rect 8895 14368 9404 14396
rect 8895 14365 8907 14368
rect 8849 14359 8907 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 7239 14300 7420 14328
rect 7239 14297 7251 14300
rect 7193 14291 7251 14297
rect 7558 14288 7564 14340
rect 7616 14328 7622 14340
rect 9876 14328 9904 14436
rect 10226 14396 10232 14408
rect 10187 14368 10232 14396
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10336 14396 10364 14436
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11149 14467 11207 14473
rect 11149 14433 11161 14467
rect 11195 14464 11207 14467
rect 12434 14464 12440 14476
rect 11195 14436 12440 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 12434 14424 12440 14436
rect 12492 14464 12498 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12492 14436 12817 14464
rect 12492 14424 12498 14436
rect 12805 14433 12817 14436
rect 12851 14464 12863 14467
rect 12894 14464 12900 14476
rect 12851 14436 12900 14464
rect 12851 14433 12863 14436
rect 12805 14427 12863 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13072 14467 13130 14473
rect 13072 14433 13084 14467
rect 13118 14464 13130 14467
rect 13814 14464 13820 14476
rect 13118 14436 13820 14464
rect 13118 14433 13130 14436
rect 13072 14427 13130 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 13924 14464 13952 14504
rect 15856 14464 15884 14572
rect 19426 14560 19432 14572
rect 19484 14560 19490 14612
rect 13924 14436 15884 14464
rect 11054 14396 11060 14408
rect 10336 14368 11060 14396
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 7616 14300 9904 14328
rect 7616 14288 7622 14300
rect 12250 14288 12256 14340
rect 12308 14328 12314 14340
rect 14185 14331 14243 14337
rect 12308 14300 12848 14328
rect 12308 14288 12314 14300
rect 4062 14260 4068 14272
rect 4023 14232 4068 14260
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 4706 14220 4712 14272
rect 4764 14260 4770 14272
rect 5166 14260 5172 14272
rect 4764 14232 5172 14260
rect 4764 14220 4770 14232
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 6089 14263 6147 14269
rect 6089 14229 6101 14263
rect 6135 14260 6147 14263
rect 8386 14260 8392 14272
rect 6135 14232 8392 14260
rect 6135 14229 6147 14232
rect 6089 14223 6147 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 10410 14260 10416 14272
rect 8536 14232 10416 14260
rect 8536 14220 8542 14232
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 10689 14263 10747 14269
rect 10689 14229 10701 14263
rect 10735 14260 10747 14263
rect 11054 14260 11060 14272
rect 10735 14232 11060 14260
rect 10735 14229 10747 14232
rect 10689 14223 10747 14229
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 12820 14260 12848 14300
rect 14185 14297 14197 14331
rect 14231 14328 14243 14331
rect 14550 14328 14556 14340
rect 14231 14300 14556 14328
rect 14231 14297 14243 14300
rect 14185 14291 14243 14297
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 13998 14260 14004 14272
rect 12820 14232 14004 14260
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 1762 14056 1768 14068
rect 1535 14028 1768 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 2038 14016 2044 14068
rect 2096 14016 2102 14068
rect 3694 14056 3700 14068
rect 2516 14028 3700 14056
rect 2056 13988 2084 14016
rect 2516 13988 2544 14028
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 4157 14059 4215 14065
rect 4157 14025 4169 14059
rect 4203 14056 4215 14059
rect 4890 14056 4896 14068
rect 4203 14028 4896 14056
rect 4203 14025 4215 14028
rect 4157 14019 4215 14025
rect 4890 14016 4896 14028
rect 4948 14016 4954 14068
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7650 14056 7656 14068
rect 6871 14028 7656 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 7834 14056 7840 14068
rect 7795 14028 7840 14056
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 9306 14056 9312 14068
rect 9267 14028 9312 14056
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 13814 14056 13820 14068
rect 9456 14028 13676 14056
rect 13775 14028 13820 14056
rect 9456 14016 9462 14028
rect 2056 13960 2544 13988
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2516 13929 2544 13960
rect 3881 13991 3939 13997
rect 3881 13957 3893 13991
rect 3927 13988 3939 13991
rect 4338 13988 4344 14000
rect 3927 13960 4344 13988
rect 3927 13957 3939 13960
rect 3881 13951 3939 13957
rect 4338 13948 4344 13960
rect 4396 13988 4402 14000
rect 5169 13991 5227 13997
rect 4396 13960 4752 13988
rect 4396 13948 4402 13960
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 3602 13880 3608 13932
rect 3660 13920 3666 13932
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3660 13892 3985 13920
rect 3660 13880 3666 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4724 13929 4752 13960
rect 5169 13957 5181 13991
rect 5215 13988 5227 13991
rect 6270 13988 6276 14000
rect 5215 13960 6276 13988
rect 5215 13957 5227 13960
rect 5169 13951 5227 13957
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 8662 13948 8668 14000
rect 8720 13988 8726 14000
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8720 13960 8861 13988
rect 8720 13948 8726 13960
rect 8849 13957 8861 13960
rect 8895 13988 8907 13991
rect 10870 13988 10876 14000
rect 8895 13960 10876 13988
rect 8895 13957 8907 13960
rect 8849 13951 8907 13957
rect 10870 13948 10876 13960
rect 10928 13948 10934 14000
rect 10965 13991 11023 13997
rect 10965 13957 10977 13991
rect 11011 13988 11023 13991
rect 11790 13988 11796 14000
rect 11011 13960 11796 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 13648 13988 13676 14028
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 16025 14059 16083 14065
rect 16025 14056 16037 14059
rect 13924 14028 16037 14056
rect 13924 13988 13952 14028
rect 16025 14025 16037 14028
rect 16071 14025 16083 14059
rect 16025 14019 16083 14025
rect 13648 13960 13952 13988
rect 4617 13923 4675 13929
rect 4617 13920 4629 13923
rect 4120 13892 4629 13920
rect 4120 13880 4126 13892
rect 4617 13889 4629 13892
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13889 4767 13923
rect 5718 13920 5724 13932
rect 5679 13892 5724 13920
rect 4709 13883 4767 13889
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7650 13920 7656 13932
rect 7515 13892 7656 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7650 13880 7656 13892
rect 7708 13920 7714 13932
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 7708 13892 8401 13920
rect 7708 13880 7714 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8389 13883 8447 13889
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9858 13920 9864 13932
rect 8996 13892 9864 13920
rect 8996 13880 9002 13892
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10226 13920 10232 13932
rect 9999 13892 10232 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 10410 13880 10416 13932
rect 10468 13920 10474 13932
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 10468 13892 11437 13920
rect 10468 13880 10474 13892
rect 11425 13889 11437 13892
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 11609 13923 11667 13929
rect 11609 13889 11621 13923
rect 11655 13920 11667 13923
rect 11698 13920 11704 13932
rect 11655 13892 11704 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 12066 13880 12072 13932
rect 12124 13920 12130 13932
rect 12124 13892 12572 13920
rect 12124 13880 12130 13892
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 1949 13855 2007 13861
rect 1949 13852 1961 13855
rect 1452 13824 1961 13852
rect 1452 13812 1458 13824
rect 1949 13821 1961 13824
rect 1995 13821 2007 13855
rect 1949 13815 2007 13821
rect 2768 13855 2826 13861
rect 2768 13821 2780 13855
rect 2814 13852 2826 13855
rect 3050 13852 3056 13864
rect 2814 13824 3056 13852
rect 2814 13821 2826 13824
rect 2768 13815 2826 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4525 13855 4583 13861
rect 4525 13852 4537 13855
rect 4212 13824 4537 13852
rect 4212 13812 4218 13824
rect 4525 13821 4537 13824
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5500 13824 5641 13852
rect 5500 13812 5506 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 6362 13852 6368 13864
rect 6323 13824 6368 13852
rect 5629 13815 5687 13821
rect 6362 13812 6368 13824
rect 6420 13812 6426 13864
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 8297 13855 8355 13861
rect 8297 13852 8309 13855
rect 6972 13824 8309 13852
rect 6972 13812 6978 13824
rect 8297 13821 8309 13824
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9398 13852 9404 13864
rect 9079 13824 9404 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 10870 13852 10876 13864
rect 9508 13824 10876 13852
rect 1857 13787 1915 13793
rect 1857 13753 1869 13787
rect 1903 13784 1915 13787
rect 3418 13784 3424 13796
rect 1903 13756 3424 13784
rect 1903 13753 1915 13756
rect 1857 13747 1915 13753
rect 3418 13744 3424 13756
rect 3476 13744 3482 13796
rect 3786 13744 3792 13796
rect 3844 13784 3850 13796
rect 9508 13784 9536 13824
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 12158 13852 12164 13864
rect 11112 13824 12164 13852
rect 11112 13812 11118 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12544 13852 12572 13892
rect 12693 13855 12751 13861
rect 12693 13852 12705 13855
rect 12544 13824 12705 13852
rect 12693 13821 12705 13824
rect 12739 13821 12751 13855
rect 12693 13815 12751 13821
rect 12986 13812 12992 13864
rect 13044 13852 13050 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 13044 13824 14657 13852
rect 13044 13812 13050 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14912 13855 14970 13861
rect 14912 13821 14924 13855
rect 14958 13852 14970 13855
rect 18690 13852 18696 13864
rect 14958 13824 18696 13852
rect 14958 13821 14970 13824
rect 14912 13815 14970 13821
rect 18690 13812 18696 13824
rect 18748 13812 18754 13864
rect 3844 13756 9536 13784
rect 9677 13787 9735 13793
rect 3844 13744 3850 13756
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 10321 13787 10379 13793
rect 10321 13784 10333 13787
rect 9723 13756 10333 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 10321 13753 10333 13756
rect 10367 13753 10379 13787
rect 15930 13784 15936 13796
rect 10321 13747 10379 13753
rect 14936 13756 15936 13784
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 3878 13716 3884 13728
rect 3200 13688 3884 13716
rect 3200 13676 3206 13688
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 3973 13719 4031 13725
rect 3973 13685 3985 13719
rect 4019 13716 4031 13719
rect 5350 13716 5356 13728
rect 4019 13688 5356 13716
rect 4019 13685 4031 13688
rect 3973 13679 4031 13685
rect 5350 13676 5356 13688
rect 5408 13716 5414 13728
rect 5537 13719 5595 13725
rect 5537 13716 5549 13719
rect 5408 13688 5549 13716
rect 5408 13676 5414 13688
rect 5537 13685 5549 13688
rect 5583 13685 5595 13719
rect 5537 13679 5595 13685
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 6181 13719 6239 13725
rect 6181 13716 6193 13719
rect 5868 13688 6193 13716
rect 5868 13676 5874 13688
rect 6181 13685 6193 13688
rect 6227 13716 6239 13719
rect 6730 13716 6736 13728
rect 6227 13688 6736 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 7190 13716 7196 13728
rect 7151 13688 7196 13716
rect 7190 13676 7196 13688
rect 7248 13676 7254 13728
rect 7282 13676 7288 13728
rect 7340 13716 7346 13728
rect 7340 13688 7385 13716
rect 7340 13676 7346 13688
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7524 13688 8217 13716
rect 7524 13676 7530 13688
rect 8205 13685 8217 13688
rect 8251 13685 8263 13719
rect 9766 13716 9772 13728
rect 9727 13688 9772 13716
rect 8205 13679 8263 13685
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 11333 13719 11391 13725
rect 11333 13716 11345 13719
rect 9916 13688 11345 13716
rect 9916 13676 9922 13688
rect 11333 13685 11345 13688
rect 11379 13716 11391 13719
rect 11514 13716 11520 13728
rect 11379 13688 11520 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11977 13719 12035 13725
rect 11977 13685 11989 13719
rect 12023 13716 12035 13719
rect 12434 13716 12440 13728
rect 12023 13688 12440 13716
rect 12023 13685 12035 13688
rect 11977 13679 12035 13685
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 12802 13676 12808 13728
rect 12860 13716 12866 13728
rect 14936 13716 14964 13756
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 12860 13688 14964 13716
rect 12860 13676 12866 13688
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 16022 13716 16028 13728
rect 15068 13688 16028 13716
rect 15068 13676 15074 13688
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 2133 13515 2191 13521
rect 2133 13481 2145 13515
rect 2179 13512 2191 13515
rect 2682 13512 2688 13524
rect 2179 13484 2688 13512
rect 2179 13481 2191 13484
rect 2133 13475 2191 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 3326 13512 3332 13524
rect 3287 13484 3332 13512
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 5445 13515 5503 13521
rect 5445 13481 5457 13515
rect 5491 13512 5503 13515
rect 5718 13512 5724 13524
rect 5491 13484 5724 13512
rect 5491 13481 5503 13484
rect 5445 13475 5503 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 8757 13515 8815 13521
rect 8757 13512 8769 13515
rect 7800 13484 8769 13512
rect 7800 13472 7806 13484
rect 8757 13481 8769 13484
rect 8803 13481 8815 13515
rect 8757 13475 8815 13481
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 10502 13512 10508 13524
rect 8904 13484 10508 13512
rect 8904 13472 8910 13484
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 10594 13472 10600 13524
rect 10652 13512 10658 13524
rect 10870 13512 10876 13524
rect 10652 13484 10876 13512
rect 10652 13472 10658 13484
rect 10870 13472 10876 13484
rect 10928 13512 10934 13524
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 10928 13484 11069 13512
rect 10928 13472 10934 13484
rect 11057 13481 11069 13484
rect 11103 13481 11115 13515
rect 11057 13475 11115 13481
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 11848 13484 13369 13512
rect 11848 13472 11854 13484
rect 13357 13481 13369 13484
rect 13403 13481 13415 13515
rect 13357 13475 13415 13481
rect 14369 13515 14427 13521
rect 14369 13481 14381 13515
rect 14415 13512 14427 13515
rect 14550 13512 14556 13524
rect 14415 13484 14556 13512
rect 14415 13481 14427 13484
rect 14369 13475 14427 13481
rect 14550 13472 14556 13484
rect 14608 13512 14614 13524
rect 15010 13512 15016 13524
rect 14608 13484 15016 13512
rect 14608 13472 14614 13484
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 15160 13484 15301 13512
rect 15160 13472 15166 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 16301 13515 16359 13521
rect 16301 13481 16313 13515
rect 16347 13481 16359 13515
rect 16666 13512 16672 13524
rect 16627 13484 16672 13512
rect 16301 13475 16359 13481
rect 1486 13404 1492 13456
rect 1544 13444 1550 13456
rect 1673 13447 1731 13453
rect 1673 13444 1685 13447
rect 1544 13416 1685 13444
rect 1544 13404 1550 13416
rect 1673 13413 1685 13416
rect 1719 13413 1731 13447
rect 1673 13407 1731 13413
rect 2056 13416 3096 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2056 13376 2084 13416
rect 1443 13348 2084 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2314 13336 2320 13388
rect 2372 13376 2378 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2372 13348 2513 13376
rect 2372 13336 2378 13348
rect 2501 13345 2513 13348
rect 2547 13345 2559 13379
rect 2501 13339 2559 13345
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 2866 13376 2872 13388
rect 2639 13348 2872 13376
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2188 13280 2697 13308
rect 2188 13268 2194 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 3068 13308 3096 13416
rect 3418 13404 3424 13456
rect 3476 13444 3482 13456
rect 4062 13444 4068 13456
rect 3476 13416 4068 13444
rect 3476 13404 3482 13416
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 4338 13453 4344 13456
rect 4332 13444 4344 13453
rect 4299 13416 4344 13444
rect 4332 13407 4344 13416
rect 4338 13404 4344 13407
rect 4396 13404 4402 13456
rect 4540 13416 6215 13444
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3878 13376 3884 13388
rect 3191 13348 3884 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4540 13376 4568 13416
rect 3988 13348 4568 13376
rect 5721 13379 5779 13385
rect 3988 13308 4016 13348
rect 5721 13345 5733 13379
rect 5767 13376 5779 13379
rect 5810 13376 5816 13388
rect 5767 13348 5816 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 5994 13385 6000 13388
rect 5988 13339 6000 13385
rect 6052 13376 6058 13388
rect 6187 13376 6215 13416
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 16316 13444 16344 13475
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 9824 13416 16344 13444
rect 9824 13404 9830 13416
rect 7098 13376 7104 13388
rect 6052 13348 6088 13376
rect 6187 13348 7104 13376
rect 5994 13336 6000 13339
rect 6052 13336 6058 13348
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7650 13385 7656 13388
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 7644 13376 7656 13385
rect 7239 13348 7656 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 7644 13339 7656 13348
rect 7650 13336 7656 13339
rect 7708 13336 7714 13388
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 7984 13348 9628 13376
rect 7984 13336 7990 13348
rect 3068 13280 4016 13308
rect 4065 13311 4123 13317
rect 2685 13271 2743 13277
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 3694 13200 3700 13252
rect 3752 13240 3758 13252
rect 4080 13240 4108 13271
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 6788 13280 7389 13308
rect 6788 13268 6794 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 9600 13308 9628 13348
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9861 13379 9919 13385
rect 9861 13376 9873 13379
rect 9732 13348 9873 13376
rect 9732 13336 9738 13348
rect 9861 13345 9873 13348
rect 9907 13345 9919 13379
rect 10778 13376 10784 13388
rect 9861 13339 9919 13345
rect 9968 13348 10784 13376
rect 9968 13308 9996 13348
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11698 13376 11704 13388
rect 11011 13348 11704 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 11848 13348 11989 13376
rect 11848 13336 11854 13348
rect 11977 13345 11989 13348
rect 12023 13345 12035 13379
rect 12894 13376 12900 13388
rect 11977 13339 12035 13345
rect 12268 13348 12900 13376
rect 9600 13280 9996 13308
rect 7377 13271 7435 13277
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10100 13280 10145 13308
rect 10100 13268 10106 13280
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10284 13280 11192 13308
rect 10284 13268 10290 13280
rect 3752 13212 4108 13240
rect 7101 13243 7159 13249
rect 3752 13200 3758 13212
rect 7101 13209 7113 13243
rect 7147 13240 7159 13243
rect 7193 13243 7251 13249
rect 7193 13240 7205 13243
rect 7147 13212 7205 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 7193 13209 7205 13212
rect 7239 13209 7251 13243
rect 9950 13240 9956 13252
rect 7193 13203 7251 13209
rect 8312 13212 9956 13240
rect 3602 13132 3608 13184
rect 3660 13172 3666 13184
rect 8312 13172 8340 13212
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 11164 13240 11192 13280
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 12268 13317 12296 13348
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13265 13379 13323 13385
rect 13265 13345 13277 13379
rect 13311 13376 13323 13379
rect 13538 13376 13544 13388
rect 13311 13348 13544 13376
rect 13311 13345 13323 13348
rect 13265 13339 13323 13345
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 14182 13336 14188 13388
rect 14240 13376 14246 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 14240 13348 14289 13376
rect 14240 13336 14246 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 14277 13339 14335 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 11425 13311 11483 13317
rect 11296 13280 11341 13308
rect 11296 13268 11302 13280
rect 11425 13277 11437 13311
rect 11471 13308 11483 13311
rect 12069 13311 12127 13317
rect 12069 13308 12081 13311
rect 11471 13280 12081 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 12069 13277 12081 13280
rect 12115 13277 12127 13311
rect 12069 13271 12127 13277
rect 12253 13311 12311 13317
rect 12253 13277 12265 13311
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12584 13280 13461 13308
rect 12584 13268 12590 13280
rect 13449 13277 13461 13280
rect 13495 13308 13507 13311
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 13495 13280 14473 13308
rect 13495 13277 13507 13280
rect 13449 13271 13507 13277
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 14608 13280 15761 13308
rect 14608 13268 14614 13280
rect 15749 13277 15761 13280
rect 15795 13277 15807 13311
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15749 13271 15807 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16758 13308 16764 13320
rect 16719 13280 16764 13308
rect 16758 13268 16764 13280
rect 16816 13268 16822 13320
rect 16853 13311 16911 13317
rect 16853 13277 16865 13311
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 12802 13240 12808 13252
rect 11164 13212 12808 13240
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 12897 13243 12955 13249
rect 12897 13209 12909 13243
rect 12943 13240 12955 13243
rect 15010 13240 15016 13252
rect 12943 13212 15016 13240
rect 12943 13209 12955 13212
rect 12897 13203 12955 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 15948 13240 15976 13268
rect 16868 13240 16896 13271
rect 15948 13212 16896 13240
rect 3660 13144 8340 13172
rect 3660 13132 3666 13144
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10597 13175 10655 13181
rect 10597 13172 10609 13175
rect 10100 13144 10609 13172
rect 10100 13132 10106 13144
rect 10597 13141 10609 13144
rect 10643 13141 10655 13175
rect 10597 13135 10655 13141
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 10744 13144 11437 13172
rect 10744 13132 10750 13144
rect 11425 13141 11437 13144
rect 11471 13141 11483 13175
rect 11425 13135 11483 13141
rect 11609 13175 11667 13181
rect 11609 13141 11621 13175
rect 11655 13172 11667 13175
rect 13722 13172 13728 13184
rect 11655 13144 13728 13172
rect 11655 13141 11667 13144
rect 11609 13135 11667 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 13909 13175 13967 13181
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 14918 13172 14924 13184
rect 13955 13144 14924 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 3418 12928 3424 12980
rect 3476 12928 3482 12980
rect 3694 12928 3700 12980
rect 3752 12928 3758 12980
rect 3970 12968 3976 12980
rect 3931 12940 3976 12968
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 5810 12968 5816 12980
rect 4632 12940 5816 12968
rect 3142 12860 3148 12912
rect 3200 12900 3206 12912
rect 3436 12900 3464 12928
rect 3200 12872 3464 12900
rect 3712 12900 3740 12928
rect 4632 12900 4660 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 5994 12968 6000 12980
rect 5955 12940 6000 12968
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6825 12971 6883 12977
rect 6825 12937 6837 12971
rect 6871 12968 6883 12971
rect 7282 12968 7288 12980
rect 6871 12940 7288 12968
rect 6871 12937 6883 12940
rect 6825 12931 6883 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 9674 12968 9680 12980
rect 7432 12940 9260 12968
rect 9635 12940 9680 12968
rect 7432 12928 7438 12940
rect 3712 12872 4660 12900
rect 6012 12900 6040 12928
rect 6730 12900 6736 12912
rect 6012 12872 6736 12900
rect 3200 12860 3206 12872
rect 2406 12832 2412 12844
rect 2367 12804 2412 12832
rect 2406 12792 2412 12804
rect 2464 12792 2470 12844
rect 3252 12841 3280 12872
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12832 3479 12835
rect 3694 12832 3700 12844
rect 3467 12804 3700 12832
rect 3467 12801 3479 12804
rect 3421 12795 3479 12801
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4632 12841 4660 12872
rect 6730 12860 6736 12872
rect 6788 12900 6794 12912
rect 9232 12909 9260 12940
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 10226 12928 10232 12980
rect 10284 12928 10290 12980
rect 12066 12968 12072 12980
rect 10336 12940 12072 12968
rect 9217 12903 9275 12909
rect 6788 12872 7420 12900
rect 6788 12860 6794 12872
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 7392 12841 7420 12872
rect 9217 12869 9229 12903
rect 9263 12900 9275 12903
rect 10244 12900 10272 12928
rect 9263 12872 10272 12900
rect 9263 12869 9275 12872
rect 9217 12863 9275 12869
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 6328 12804 7297 12832
rect 6328 12792 6334 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 7650 12832 7656 12844
rect 7423 12804 7656 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 10336 12841 10364 12940
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12250 12928 12256 12980
rect 12308 12968 12314 12980
rect 12308 12940 12480 12968
rect 12308 12928 12314 12940
rect 12452 12900 12480 12940
rect 12618 12928 12624 12980
rect 12676 12968 12682 12980
rect 17126 12968 17132 12980
rect 12676 12940 17132 12968
rect 12676 12928 12682 12940
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 14274 12900 14280 12912
rect 12452 12872 12664 12900
rect 14187 12872 14280 12900
rect 10321 12835 10379 12841
rect 7800 12804 7972 12832
rect 7800 12792 7806 12804
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3191 12736 3617 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3786 12764 3792 12776
rect 3747 12736 3792 12764
rect 3605 12727 3663 12733
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 4884 12767 4942 12773
rect 4884 12733 4896 12767
rect 4930 12764 4942 12767
rect 5718 12764 5724 12776
rect 4930 12736 5724 12764
rect 4930 12733 4942 12736
rect 4884 12727 4942 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 6822 12724 6828 12776
rect 6880 12764 6886 12776
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 6880 12736 7849 12764
rect 6880 12724 6886 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7944 12764 7972 12804
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 12437 12835 12495 12841
rect 12437 12832 12449 12835
rect 11756 12804 12449 12832
rect 11756 12792 11762 12804
rect 12437 12801 12449 12804
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 8093 12767 8151 12773
rect 8093 12764 8105 12767
rect 7944 12736 8105 12764
rect 7837 12727 7895 12733
rect 8093 12733 8105 12736
rect 8139 12733 8151 12767
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 8093 12727 8151 12733
rect 10042 12724 10048 12736
rect 10100 12724 10106 12776
rect 10689 12767 10747 12773
rect 10689 12733 10701 12767
rect 10735 12764 10747 12767
rect 12636 12764 12664 12872
rect 14274 12860 14280 12872
rect 14332 12900 14338 12912
rect 14332 12872 16160 12900
rect 14332 12860 14338 12872
rect 12805 12835 12863 12841
rect 12805 12801 12817 12835
rect 12851 12832 12863 12835
rect 12897 12835 12955 12841
rect 12897 12832 12909 12835
rect 12851 12804 12909 12832
rect 12851 12801 12863 12804
rect 12805 12795 12863 12801
rect 12897 12801 12909 12804
rect 12943 12801 12955 12835
rect 14182 12832 14188 12844
rect 12897 12795 12955 12801
rect 13924 12804 14188 12832
rect 13924 12764 13952 12804
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 15102 12832 15108 12844
rect 15063 12804 15108 12832
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 16132 12841 16160 12872
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 14550 12764 14556 12776
rect 10735 12736 12480 12764
rect 12636 12736 13952 12764
rect 14108 12736 14556 12764
rect 10735 12733 10747 12736
rect 10689 12727 10747 12733
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12696 2283 12699
rect 4982 12696 4988 12708
rect 2271 12668 4988 12696
rect 2271 12665 2283 12668
rect 2225 12659 2283 12665
rect 4982 12656 4988 12668
rect 5040 12656 5046 12708
rect 7006 12656 7012 12708
rect 7064 12696 7070 12708
rect 7193 12699 7251 12705
rect 7193 12696 7205 12699
rect 7064 12668 7205 12696
rect 7064 12656 7070 12668
rect 7193 12665 7205 12668
rect 7239 12696 7251 12699
rect 8938 12696 8944 12708
rect 7239 12668 8944 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 10226 12656 10232 12708
rect 10284 12696 10290 12708
rect 10704 12696 10732 12727
rect 12452 12708 12480 12736
rect 10284 12668 10732 12696
rect 10956 12699 11014 12705
rect 10284 12656 10290 12668
rect 10956 12665 10968 12699
rect 11002 12696 11014 12699
rect 11238 12696 11244 12708
rect 11002 12668 11244 12696
rect 11002 12665 11014 12668
rect 10956 12659 11014 12665
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 12434 12656 12440 12708
rect 12492 12696 12498 12708
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12492 12668 12817 12696
rect 12492 12656 12498 12668
rect 12805 12665 12817 12668
rect 12851 12665 12863 12699
rect 12805 12659 12863 12665
rect 13164 12699 13222 12705
rect 13164 12665 13176 12699
rect 13210 12696 13222 12699
rect 13814 12696 13820 12708
rect 13210 12668 13820 12696
rect 13210 12665 13222 12668
rect 13164 12659 13222 12665
rect 13814 12656 13820 12668
rect 13872 12656 13878 12708
rect 1578 12588 1584 12640
rect 1636 12628 1642 12640
rect 1765 12631 1823 12637
rect 1765 12628 1777 12631
rect 1636 12600 1777 12628
rect 1636 12588 1642 12600
rect 1765 12597 1777 12600
rect 1811 12597 1823 12631
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 1765 12591 1823 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3605 12631 3663 12637
rect 2832 12600 2877 12628
rect 2832 12588 2838 12600
rect 3605 12597 3617 12631
rect 3651 12628 3663 12631
rect 5902 12628 5908 12640
rect 3651 12600 5908 12628
rect 3651 12597 3663 12600
rect 3605 12591 3663 12597
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 7374 12588 7380 12640
rect 7432 12628 7438 12640
rect 7742 12628 7748 12640
rect 7432 12600 7748 12628
rect 7432 12588 7438 12600
rect 7742 12588 7748 12600
rect 7800 12588 7806 12640
rect 10137 12631 10195 12637
rect 10137 12597 10149 12631
rect 10183 12628 10195 12631
rect 11422 12628 11428 12640
rect 10183 12600 11428 12628
rect 10183 12597 10195 12600
rect 10137 12591 10195 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 14108 12628 14136 12736
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 14918 12764 14924 12776
rect 14879 12736 14924 12764
rect 14918 12724 14924 12736
rect 14976 12724 14982 12776
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 15381 12767 15439 12773
rect 15068 12736 15113 12764
rect 15068 12724 15074 12736
rect 15381 12733 15393 12767
rect 15427 12764 15439 12767
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 15427 12736 15945 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15933 12733 15945 12736
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 16025 12699 16083 12705
rect 16025 12696 16037 12699
rect 14568 12668 16037 12696
rect 14568 12637 14596 12668
rect 16025 12665 16037 12668
rect 16071 12665 16083 12699
rect 16025 12659 16083 12665
rect 12032 12600 14136 12628
rect 14553 12631 14611 12637
rect 12032 12588 12038 12600
rect 14553 12597 14565 12631
rect 14599 12597 14611 12631
rect 14553 12591 14611 12597
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 15381 12631 15439 12637
rect 15381 12628 15393 12631
rect 15068 12600 15393 12628
rect 15068 12588 15074 12600
rect 15381 12597 15393 12600
rect 15427 12597 15439 12631
rect 15562 12628 15568 12640
rect 15523 12600 15568 12628
rect 15381 12591 15439 12597
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1765 12427 1823 12433
rect 1765 12393 1777 12427
rect 1811 12424 1823 12427
rect 2130 12424 2136 12436
rect 1811 12396 2136 12424
rect 1811 12393 1823 12396
rect 1765 12387 1823 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2271 12396 2789 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 3142 12424 3148 12436
rect 3055 12396 3148 12424
rect 2777 12387 2835 12393
rect 3142 12384 3148 12396
rect 3200 12424 3206 12436
rect 3326 12424 3332 12436
rect 3200 12396 3332 12424
rect 3200 12384 3206 12396
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 4246 12384 4252 12436
rect 4304 12424 4310 12436
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 4304 12396 4445 12424
rect 4304 12384 4310 12396
rect 4433 12393 4445 12396
rect 4479 12393 4491 12427
rect 4433 12387 4491 12393
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 4798 12424 4804 12436
rect 4571 12396 4804 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5261 12427 5319 12433
rect 5261 12393 5273 12427
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 5276 12356 5304 12387
rect 5718 12384 5724 12436
rect 5776 12424 5782 12436
rect 6546 12424 6552 12436
rect 5776 12396 6552 12424
rect 5776 12384 5782 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 6972 12396 7573 12424
rect 6972 12384 6978 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 8938 12424 8944 12436
rect 8899 12396 8944 12424
rect 7561 12387 7619 12393
rect 8938 12384 8944 12396
rect 8996 12424 9002 12436
rect 9582 12424 9588 12436
rect 8996 12396 9588 12424
rect 8996 12384 9002 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 10870 12424 10876 12436
rect 9732 12396 10876 12424
rect 9732 12384 9738 12396
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12342 12424 12348 12436
rect 12303 12396 12348 12424
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14550 12424 14556 12436
rect 14240 12396 14556 12424
rect 14240 12384 14246 12396
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 4212 12328 5304 12356
rect 8021 12359 8079 12365
rect 4212 12316 4218 12328
rect 8021 12325 8033 12359
rect 8067 12356 8079 12359
rect 9122 12356 9128 12368
rect 8067 12328 9128 12356
rect 8067 12325 8079 12328
rect 8021 12319 8079 12325
rect 9122 12316 9128 12328
rect 9180 12356 9186 12368
rect 10042 12356 10048 12368
rect 9180 12328 10048 12356
rect 9180 12316 9186 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10594 12356 10600 12368
rect 10152 12328 10600 12356
rect 2133 12291 2191 12297
rect 2133 12257 2145 12291
rect 2179 12288 2191 12291
rect 2774 12288 2780 12300
rect 2179 12260 2780 12288
rect 2179 12257 2191 12260
rect 2133 12251 2191 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 3237 12291 3295 12297
rect 3237 12257 3249 12291
rect 3283 12288 3295 12291
rect 3326 12288 3332 12300
rect 3283 12260 3332 12288
rect 3283 12257 3295 12260
rect 3237 12251 3295 12257
rect 3326 12248 3332 12260
rect 3384 12288 3390 12300
rect 3970 12288 3976 12300
rect 3384 12260 3976 12288
rect 3384 12248 3390 12260
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 5083 12291 5141 12297
rect 5083 12257 5095 12291
rect 5129 12257 5141 12291
rect 5083 12251 5141 12257
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2498 12220 2504 12232
rect 2455 12192 2504 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 3694 12220 3700 12232
rect 3467 12192 3700 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 3694 12180 3700 12192
rect 3752 12220 3758 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 3752 12192 4629 12220
rect 3752 12180 3758 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 5092 12152 5120 12251
rect 5810 12248 5816 12300
rect 5868 12288 5874 12300
rect 6178 12297 6184 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5868 12260 5917 12288
rect 5868 12248 5874 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 6172 12288 6184 12297
rect 6139 12260 6184 12288
rect 5905 12251 5963 12257
rect 6172 12251 6184 12260
rect 6178 12248 6184 12251
rect 6236 12248 6242 12300
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 7800 12260 7941 12288
rect 7800 12248 7806 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 10152 12288 10180 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 13808 12359 13866 12365
rect 10744 12328 11192 12356
rect 10744 12316 10750 12328
rect 8536 12260 10180 12288
rect 10496 12291 10554 12297
rect 8536 12248 8542 12260
rect 10496 12257 10508 12291
rect 10542 12288 10554 12291
rect 11054 12288 11060 12300
rect 10542 12260 11060 12288
rect 10542 12257 10554 12260
rect 10496 12251 10554 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11164 12288 11192 12328
rect 13808 12325 13820 12359
rect 13854 12356 13866 12359
rect 13906 12356 13912 12368
rect 13854 12328 13912 12356
rect 13854 12325 13866 12328
rect 13808 12319 13866 12325
rect 13906 12316 13912 12328
rect 13964 12316 13970 12368
rect 12253 12291 12311 12297
rect 12253 12288 12265 12291
rect 11164 12260 12265 12288
rect 12253 12257 12265 12260
rect 12299 12257 12311 12291
rect 12253 12251 12311 12257
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 12584 12260 13553 12288
rect 12584 12248 12590 12260
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 7708 12192 8125 12220
rect 7708 12180 7714 12192
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 9033 12223 9091 12229
rect 9033 12189 9045 12223
rect 9079 12189 9091 12223
rect 9033 12183 9091 12189
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9674 12220 9680 12232
rect 9635 12192 9680 12220
rect 9217 12183 9275 12189
rect 9048 12152 9076 12183
rect 1912 12124 5120 12152
rect 7208 12124 9076 12152
rect 9232 12152 9260 12183
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10226 12220 10232 12232
rect 9824 12192 10232 12220
rect 9824 12180 9830 12192
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 13078 12220 13084 12232
rect 13039 12192 13084 12220
rect 12437 12183 12495 12189
rect 10134 12152 10140 12164
rect 9232 12124 10140 12152
rect 1912 12112 1918 12124
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 4890 12084 4896 12096
rect 4111 12056 4896 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5442 12044 5448 12096
rect 5500 12084 5506 12096
rect 7208 12084 7236 12124
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 11238 12112 11244 12164
rect 11296 12112 11302 12164
rect 5500 12056 7236 12084
rect 7285 12087 7343 12093
rect 5500 12044 5506 12056
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 7374 12084 7380 12096
rect 7331 12056 7380 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 11146 12084 11152 12096
rect 8619 12056 11152 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11256 12084 11284 12112
rect 11609 12087 11667 12093
rect 11609 12084 11621 12087
rect 11256 12056 11621 12084
rect 11609 12053 11621 12056
rect 11655 12084 11667 12087
rect 12452 12084 12480 12183
rect 13078 12180 13084 12192
rect 13136 12180 13142 12232
rect 11655 12056 12480 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14458 12084 14464 12096
rect 13964 12056 14464 12084
rect 13964 12044 13970 12056
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14918 12084 14924 12096
rect 14879 12056 14924 12084
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 4982 11880 4988 11892
rect 2556 11852 3740 11880
rect 4943 11852 4988 11880
rect 2556 11840 2562 11852
rect 3712 11821 3740 11852
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 7377 11883 7435 11889
rect 7377 11880 7389 11883
rect 5132 11852 7389 11880
rect 5132 11840 5138 11852
rect 7377 11849 7389 11852
rect 7423 11849 7435 11883
rect 7377 11843 7435 11849
rect 10873 11883 10931 11889
rect 10873 11849 10885 11883
rect 10919 11880 10931 11883
rect 12342 11880 12348 11892
rect 10919 11852 12348 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 14918 11880 14924 11892
rect 13412 11852 14924 11880
rect 13412 11840 13418 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 3697 11815 3755 11821
rect 3697 11781 3709 11815
rect 3743 11812 3755 11815
rect 3743 11784 5580 11812
rect 3743 11781 3755 11784
rect 3697 11775 3755 11781
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 3712 11716 4537 11744
rect 3712 11688 3740 11716
rect 4525 11713 4537 11716
rect 4571 11713 4583 11747
rect 4525 11707 4583 11713
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5552 11753 5580 11784
rect 8662 11772 8668 11824
rect 8720 11812 8726 11824
rect 8720 11784 12388 11812
rect 8720 11772 8726 11784
rect 12360 11756 12388 11784
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 4948 11716 5457 11744
rect 4948 11704 4954 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5960 11716 6009 11744
rect 5960 11704 5966 11716
rect 5997 11713 6009 11716
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 9306 11744 9312 11756
rect 8067 11716 9312 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 9456 11716 10793 11744
rect 9456 11704 9462 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 1578 11676 1584 11688
rect 1539 11648 1584 11676
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 2096 11648 2329 11676
rect 2096 11636 2102 11648
rect 2317 11645 2329 11648
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2584 11679 2642 11685
rect 2584 11645 2596 11679
rect 2630 11676 2642 11679
rect 3694 11676 3700 11688
rect 2630 11648 3700 11676
rect 2630 11645 2642 11648
rect 2584 11639 2642 11645
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 8202 11676 8208 11688
rect 7576 11648 8208 11676
rect 5353 11611 5411 11617
rect 5353 11608 5365 11611
rect 3988 11580 5365 11608
rect 3988 11549 4016 11580
rect 5353 11577 5365 11580
rect 5399 11577 5411 11611
rect 5353 11571 5411 11577
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 7576 11608 7604 11648
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 10962 11676 10968 11688
rect 8435 11648 10968 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11532 11676 11560 11707
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 14642 11744 14648 11756
rect 12492 11716 12537 11744
rect 14603 11716 14648 11744
rect 12492 11704 12498 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11744 17003 11747
rect 17218 11744 17224 11756
rect 16991 11716 17224 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 11112 11648 11560 11676
rect 11112 11636 11118 11648
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 11940 11648 12931 11676
rect 11940 11636 11946 11648
rect 5500 11580 7604 11608
rect 7745 11611 7803 11617
rect 5500 11568 5506 11580
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 7791 11580 8432 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 3973 11543 4031 11549
rect 3973 11509 3985 11543
rect 4019 11509 4031 11543
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 3973 11503 4031 11509
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 4488 11512 4533 11540
rect 4488 11500 4494 11512
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7282 11540 7288 11552
rect 6972 11512 7288 11540
rect 6972 11500 6978 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 8202 11540 8208 11552
rect 7883 11512 8208 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8404 11540 8432 11580
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 10870 11608 10876 11620
rect 8536 11580 10876 11608
rect 8536 11568 8542 11580
rect 10870 11568 10876 11580
rect 10928 11568 10934 11620
rect 11238 11608 11244 11620
rect 11151 11580 11244 11608
rect 11238 11568 11244 11580
rect 11296 11608 11302 11620
rect 12704 11611 12762 11617
rect 11296 11580 12664 11608
rect 11296 11568 11302 11580
rect 12636 11552 12664 11580
rect 12704 11577 12716 11611
rect 12750 11608 12762 11611
rect 12802 11608 12808 11620
rect 12750 11580 12808 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 12903 11608 12931 11648
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 13136 11648 14473 11676
rect 13136 11636 13142 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 16666 11676 16672 11688
rect 16627 11648 16672 11676
rect 14461 11639 14519 11645
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 14553 11611 14611 11617
rect 14553 11608 14565 11611
rect 12903 11580 14565 11608
rect 14553 11577 14565 11580
rect 14599 11577 14611 11611
rect 14553 11571 14611 11577
rect 8846 11540 8852 11552
rect 8404 11512 8852 11540
rect 8846 11500 8852 11512
rect 8904 11500 8910 11552
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9548 11512 9689 11540
rect 9548 11500 9554 11512
rect 9677 11509 9689 11512
rect 9723 11509 9735 11543
rect 9677 11503 9735 11509
rect 10781 11543 10839 11549
rect 10781 11509 10793 11543
rect 10827 11540 10839 11543
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 10827 11512 11345 11540
rect 10827 11509 10839 11512
rect 10781 11503 10839 11509
rect 11333 11509 11345 11512
rect 11379 11509 11391 11543
rect 11333 11503 11391 11509
rect 12342 11500 12348 11552
rect 12400 11540 12406 11552
rect 12526 11540 12532 11552
rect 12400 11512 12532 11540
rect 12400 11500 12406 11512
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12618 11500 12624 11552
rect 12676 11500 12682 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 14274 11540 14280 11552
rect 14139 11512 14280 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2464 11308 2789 11336
rect 2464 11296 2470 11308
rect 2777 11305 2789 11308
rect 2823 11305 2835 11339
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 2777 11299 2835 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 5258 11336 5264 11348
rect 4488 11308 5264 11336
rect 4488 11296 4494 11308
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6178 11336 6184 11348
rect 6091 11308 6184 11336
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 7064 11308 7297 11336
rect 7064 11296 7070 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 10226 11336 10232 11348
rect 7285 11299 7343 11305
rect 7944 11308 10232 11336
rect 1664 11271 1722 11277
rect 1664 11237 1676 11271
rect 1710 11268 1722 11271
rect 2498 11268 2504 11280
rect 1710 11240 2504 11268
rect 1710 11237 1722 11240
rect 1664 11231 1722 11237
rect 2498 11228 2504 11240
rect 2556 11228 2562 11280
rect 3329 11271 3387 11277
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 3786 11268 3792 11280
rect 3375 11240 3792 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 3786 11228 3792 11240
rect 3844 11228 3850 11280
rect 6196 11268 6224 11296
rect 6196 11240 7880 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 2038 11200 2044 11212
rect 1443 11172 2044 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 2038 11160 2044 11172
rect 2096 11160 2102 11212
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 5068 11203 5126 11209
rect 5068 11169 5080 11203
rect 5114 11200 5126 11203
rect 5810 11200 5816 11212
rect 5114 11172 5816 11200
rect 5114 11169 5126 11172
rect 5068 11163 5126 11169
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6914 11200 6920 11212
rect 5920 11172 6920 11200
rect 4798 11132 4804 11144
rect 4759 11104 4804 11132
rect 4798 11092 4804 11104
rect 4856 11092 4862 11144
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 5920 11064 5948 11172
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 7064 11172 7205 11200
rect 7064 11160 7070 11172
rect 7193 11169 7205 11172
rect 7239 11200 7251 11203
rect 7650 11200 7656 11212
rect 7239 11172 7656 11200
rect 7239 11169 7251 11172
rect 7193 11163 7251 11169
rect 7650 11160 7656 11172
rect 7708 11160 7714 11212
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 7377 11135 7435 11141
rect 7377 11132 7389 11135
rect 6788 11104 7389 11132
rect 6788 11092 6794 11104
rect 7377 11101 7389 11104
rect 7423 11101 7435 11135
rect 7852 11132 7880 11240
rect 7944 11209 7972 11308
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 12434 11336 12440 11348
rect 11563 11308 12440 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 14093 11339 14151 11345
rect 14093 11305 14105 11339
rect 14139 11336 14151 11339
rect 16666 11336 16672 11348
rect 14139 11308 16672 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 8478 11268 8484 11280
rect 8128 11240 8484 11268
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11169 7987 11203
rect 8128 11200 8156 11240
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 8628 11240 9168 11268
rect 8628 11228 8634 11240
rect 9140 11212 9168 11240
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 9922 11271 9980 11277
rect 9922 11268 9934 11271
rect 9364 11240 9934 11268
rect 9364 11228 9370 11240
rect 9922 11237 9934 11240
rect 9968 11237 9980 11271
rect 9922 11231 9980 11237
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 11609 11271 11667 11277
rect 11609 11268 11621 11271
rect 11204 11240 11621 11268
rect 11204 11228 11210 11240
rect 11609 11237 11621 11240
rect 11655 11237 11667 11271
rect 11609 11231 11667 11237
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12526 11268 12532 11280
rect 12391 11240 12532 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12526 11228 12532 11240
rect 12584 11228 12590 11280
rect 7929 11163 7987 11169
rect 8036 11172 8156 11200
rect 8196 11203 8254 11209
rect 8036 11132 8064 11172
rect 8196 11169 8208 11203
rect 8242 11200 8254 11203
rect 8938 11200 8944 11212
rect 8242 11172 8944 11200
rect 8242 11169 8254 11172
rect 8196 11163 8254 11169
rect 8938 11160 8944 11172
rect 8996 11160 9002 11212
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9398 11200 9404 11212
rect 9180 11172 9404 11200
rect 9180 11160 9186 11172
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 13170 11200 13176 11212
rect 12360 11172 12572 11200
rect 13131 11172 13176 11200
rect 12360 11144 12388 11172
rect 7852 11104 8064 11132
rect 7377 11095 7435 11101
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11112 11104 11713 11132
rect 11112 11092 11118 11104
rect 11701 11101 11713 11104
rect 11747 11101 11759 11135
rect 11701 11095 11759 11101
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 12544 11141 12572 11172
rect 13170 11160 13176 11172
rect 13228 11160 13234 11212
rect 13265 11203 13323 11209
rect 13265 11169 13277 11203
rect 13311 11200 13323 11203
rect 14458 11200 14464 11212
rect 13311 11172 14228 11200
rect 14419 11172 14464 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11101 12495 11135
rect 12437 11095 12495 11101
rect 12529 11135 12587 11141
rect 12529 11101 12541 11135
rect 12575 11101 12587 11135
rect 12529 11095 12587 11101
rect 4396 11036 4844 11064
rect 4396 11024 4402 11036
rect 4816 10996 4844 11036
rect 5736 11036 5948 11064
rect 6825 11067 6883 11073
rect 5736 10996 5764 11036
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 7190 11064 7196 11076
rect 6871 11036 7196 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 9306 11064 9312 11076
rect 9267 11036 9312 11064
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 11149 11067 11207 11073
rect 11149 11033 11161 11067
rect 11195 11064 11207 11067
rect 12452 11064 12480 11095
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13280 11132 13308 11163
rect 12676 11104 13308 11132
rect 13357 11135 13415 11141
rect 12676 11092 12682 11104
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 12805 11067 12863 11073
rect 12805 11064 12817 11067
rect 11195 11036 12480 11064
rect 12544 11036 12817 11064
rect 11195 11033 11207 11036
rect 11149 11027 11207 11033
rect 4816 10968 5764 10996
rect 6270 10956 6276 11008
rect 6328 10996 6334 11008
rect 9674 10996 9680 11008
rect 6328 10968 9680 10996
rect 6328 10956 6334 10968
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 11974 10996 11980 11008
rect 11935 10968 11980 10996
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12158 10956 12164 11008
rect 12216 10996 12222 11008
rect 12544 10996 12572 11036
rect 12805 11033 12817 11036
rect 12851 11033 12863 11067
rect 12805 11027 12863 11033
rect 12894 11024 12900 11076
rect 12952 11064 12958 11076
rect 13372 11064 13400 11095
rect 12952 11036 13400 11064
rect 14200 11064 14228 11172
rect 14458 11160 14464 11172
rect 14516 11160 14522 11212
rect 14550 11132 14556 11144
rect 14511 11104 14556 11132
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 14700 11104 14745 11132
rect 14700 11092 14706 11104
rect 16850 11064 16856 11076
rect 14200 11036 16856 11064
rect 12952 11024 12958 11036
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 12216 10968 12572 10996
rect 12216 10956 12222 10968
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 16574 10996 16580 11008
rect 13136 10968 16580 10996
rect 13136 10956 13142 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 3421 10795 3479 10801
rect 3421 10761 3433 10795
rect 3467 10792 3479 10795
rect 4706 10792 4712 10804
rect 3467 10764 4712 10792
rect 3467 10761 3479 10764
rect 3421 10755 3479 10761
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 7466 10792 7472 10804
rect 5951 10764 7472 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7576 10764 8524 10792
rect 5810 10724 5816 10736
rect 5723 10696 5816 10724
rect 5810 10684 5816 10696
rect 5868 10724 5874 10736
rect 7576 10724 7604 10764
rect 5868 10696 7604 10724
rect 8496 10724 8524 10764
rect 8846 10752 8852 10804
rect 8904 10792 8910 10804
rect 9217 10795 9275 10801
rect 9217 10792 9229 10795
rect 8904 10764 9229 10792
rect 8904 10752 8910 10764
rect 9217 10761 9229 10764
rect 9263 10761 9275 10795
rect 9217 10755 9275 10761
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10134 10792 10140 10804
rect 10008 10764 10140 10792
rect 10008 10752 10014 10764
rect 10134 10752 10140 10764
rect 10192 10792 10198 10804
rect 11977 10795 12035 10801
rect 10192 10764 11560 10792
rect 10192 10752 10198 10764
rect 8938 10724 8944 10736
rect 8496 10696 8800 10724
rect 8899 10696 8944 10724
rect 5868 10684 5874 10696
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6730 10656 6736 10668
rect 6595 10628 6736 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 2038 10588 2044 10600
rect 1999 10560 2044 10588
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 6270 10588 6276 10600
rect 4479 10560 4936 10588
rect 6231 10560 6276 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 2308 10523 2366 10529
rect 2308 10489 2320 10523
rect 2354 10520 2366 10523
rect 2406 10520 2412 10532
rect 2354 10492 2412 10520
rect 2354 10489 2366 10492
rect 2308 10483 2366 10489
rect 2406 10480 2412 10492
rect 2464 10480 2470 10532
rect 4614 10480 4620 10532
rect 4672 10529 4678 10532
rect 4672 10523 4736 10529
rect 4672 10489 4690 10523
rect 4724 10489 4736 10523
rect 4672 10483 4736 10489
rect 4672 10480 4678 10483
rect 4798 10480 4804 10532
rect 4856 10520 4862 10532
rect 4908 10520 4936 10560
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 6420 10560 7573 10588
rect 6420 10548 6426 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7828 10591 7886 10597
rect 7828 10557 7840 10591
rect 7874 10588 7886 10591
rect 8662 10588 8668 10600
rect 7874 10560 8668 10588
rect 7874 10557 7886 10560
rect 7828 10551 7886 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8772 10588 8800 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 9306 10684 9312 10736
rect 9364 10724 9370 10736
rect 10226 10724 10232 10736
rect 9364 10696 10088 10724
rect 10187 10696 10232 10724
rect 9364 10684 9370 10696
rect 8956 10656 8984 10684
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 8956 10628 9781 10656
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 10060 10656 10088 10696
rect 10226 10684 10232 10696
rect 10284 10724 10290 10736
rect 11532 10724 11560 10764
rect 11977 10761 11989 10795
rect 12023 10792 12035 10795
rect 12342 10792 12348 10804
rect 12023 10764 12348 10792
rect 12023 10761 12035 10764
rect 11977 10755 12035 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 13449 10795 13507 10801
rect 12492 10764 12537 10792
rect 12492 10752 12498 10764
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 14458 10792 14464 10804
rect 13495 10764 14464 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 10284 10696 10640 10724
rect 11532 10696 13124 10724
rect 10284 10684 10290 10696
rect 10612 10665 10640 10696
rect 13096 10665 13124 10696
rect 13814 10684 13820 10736
rect 13872 10724 13878 10736
rect 14277 10727 14335 10733
rect 13872 10696 14136 10724
rect 13872 10684 13878 10696
rect 10597 10659 10655 10665
rect 10060 10628 10539 10656
rect 9769 10619 9827 10625
rect 9306 10588 9312 10600
rect 8772 10560 9312 10588
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9456 10560 9689 10588
rect 9456 10548 9462 10560
rect 9677 10557 9689 10560
rect 9723 10557 9735 10591
rect 9677 10551 9735 10557
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 9916 10560 10425 10588
rect 9916 10548 9922 10560
rect 10413 10557 10425 10560
rect 10459 10557 10471 10591
rect 10511 10588 10539 10628
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13354 10656 13360 10668
rect 13127 10628 13360 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13354 10616 13360 10628
rect 13412 10616 13418 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13556 10628 14013 10656
rect 13556 10588 13584 10628
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 14108 10656 14136 10696
rect 14277 10693 14289 10727
rect 14323 10724 14335 10727
rect 15010 10724 15016 10736
rect 14323 10696 15016 10724
rect 14323 10693 14335 10696
rect 14277 10687 14335 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 14108 10628 14841 10656
rect 14001 10619 14059 10625
rect 14829 10625 14841 10628
rect 14875 10656 14887 10659
rect 15102 10656 15108 10668
rect 14875 10628 15108 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 10511 10560 13584 10588
rect 13817 10591 13875 10597
rect 10413 10551 10471 10557
rect 13817 10557 13829 10591
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 5074 10520 5080 10532
rect 4856 10492 5080 10520
rect 4856 10480 4862 10492
rect 5074 10480 5080 10492
rect 5132 10520 5138 10532
rect 6380 10520 6408 10548
rect 9585 10523 9643 10529
rect 9585 10520 9597 10523
rect 5132 10492 6408 10520
rect 8200 10492 9597 10520
rect 5132 10480 5138 10492
rect 3973 10455 4031 10461
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 5626 10452 5632 10464
rect 4019 10424 5632 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6328 10424 6377 10452
rect 6328 10412 6334 10424
rect 6365 10421 6377 10424
rect 6411 10452 6423 10455
rect 6914 10452 6920 10464
rect 6411 10424 6920 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 7101 10455 7159 10461
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 8200 10452 8228 10492
rect 9585 10489 9597 10492
rect 9631 10489 9643 10523
rect 10134 10520 10140 10532
rect 9585 10483 9643 10489
rect 9692 10492 10140 10520
rect 7147 10424 8228 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9692 10452 9720 10492
rect 10134 10480 10140 10492
rect 10192 10480 10198 10532
rect 10864 10523 10922 10529
rect 10864 10489 10876 10523
rect 10910 10520 10922 10523
rect 11054 10520 11060 10532
rect 10910 10492 11060 10520
rect 10910 10489 10922 10492
rect 10864 10483 10922 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 13832 10520 13860 10551
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 14645 10591 14703 10597
rect 14645 10588 14657 10591
rect 14332 10560 14657 10588
rect 14332 10548 14338 10560
rect 14645 10557 14657 10560
rect 14691 10557 14703 10591
rect 14645 10551 14703 10557
rect 12636 10492 13860 10520
rect 8352 10424 9720 10452
rect 8352 10412 8358 10424
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 12636 10452 12664 10492
rect 10376 10424 12664 10452
rect 10376 10412 10382 10424
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12768 10424 12817 10452
rect 12768 10412 12774 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13078 10452 13084 10464
rect 12943 10424 13084 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 13909 10455 13967 10461
rect 13909 10452 13921 10455
rect 13872 10424 13921 10452
rect 13872 10412 13878 10424
rect 13909 10421 13921 10424
rect 13955 10421 13967 10455
rect 13909 10415 13967 10421
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 14424 10424 14749 10452
rect 14424 10412 14430 10424
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14737 10415 14795 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 3234 10248 3240 10260
rect 2179 10220 3240 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 3694 10248 3700 10260
rect 3655 10220 3700 10248
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4433 10251 4491 10257
rect 4433 10217 4445 10251
rect 4479 10248 4491 10251
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4479 10220 4905 10248
rect 4479 10217 4491 10220
rect 4433 10211 4491 10217
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 4893 10211 4951 10217
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10217 5135 10251
rect 8202 10248 8208 10260
rect 8163 10220 8208 10248
rect 5077 10211 5135 10217
rect 4985 10183 5043 10189
rect 4985 10180 4997 10183
rect 1596 10152 4997 10180
rect 1596 10121 1624 10152
rect 4985 10149 4997 10152
rect 5031 10149 5043 10183
rect 5092 10180 5120 10211
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 10318 10248 10324 10260
rect 8312 10220 10324 10248
rect 8312 10180 8340 10220
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 12894 10248 12900 10260
rect 12851 10220 12900 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 14366 10248 14372 10260
rect 13127 10220 14372 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 5092 10152 8340 10180
rect 8573 10183 8631 10189
rect 4985 10143 5043 10149
rect 8573 10149 8585 10183
rect 8619 10180 8631 10183
rect 8846 10180 8852 10192
rect 8619 10152 8852 10180
rect 8619 10149 8631 10152
rect 8573 10143 8631 10149
rect 8846 10140 8852 10152
rect 8904 10140 8910 10192
rect 9766 10180 9772 10192
rect 9508 10152 9772 10180
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 2133 10115 2191 10121
rect 2133 10112 2145 10115
rect 1903 10084 2145 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 2133 10081 2145 10084
rect 2179 10081 2191 10115
rect 2133 10075 2191 10081
rect 2584 10115 2642 10121
rect 2584 10081 2596 10115
rect 2630 10112 2642 10115
rect 2866 10112 2872 10124
rect 2630 10084 2872 10112
rect 2630 10081 2642 10084
rect 2584 10075 2642 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5445 10115 5503 10121
rect 5445 10081 5457 10115
rect 5491 10112 5503 10115
rect 5626 10112 5632 10124
rect 5491 10084 5632 10112
rect 5491 10081 5503 10084
rect 5445 10075 5503 10081
rect 5626 10072 5632 10084
rect 5684 10072 5690 10124
rect 6362 10112 6368 10124
rect 6323 10084 6368 10112
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 6454 10072 6460 10124
rect 6512 10072 6518 10124
rect 6638 10121 6644 10124
rect 6632 10112 6644 10121
rect 6599 10084 6644 10112
rect 6632 10075 6644 10084
rect 6638 10072 6644 10075
rect 6696 10072 6702 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 9398 10112 9404 10124
rect 6972 10084 9404 10112
rect 6972 10072 6978 10084
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 2038 10004 2044 10056
rect 2096 10044 2102 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 2096 10016 2329 10044
rect 2096 10004 2102 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 2317 10007 2375 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5224 10016 5549 10044
rect 5224 10004 5230 10016
rect 5537 10013 5549 10016
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5810 10044 5816 10056
rect 5767 10016 5816 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5810 10004 5816 10016
rect 5868 10044 5874 10056
rect 6472 10044 6500 10072
rect 5868 10016 6500 10044
rect 5868 10004 5874 10016
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8352 10016 8677 10044
rect 8352 10004 8358 10016
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 8849 10047 8907 10053
rect 8849 10013 8861 10047
rect 8895 10044 8907 10047
rect 8938 10044 8944 10056
rect 8895 10016 8944 10044
rect 8895 10013 8907 10016
rect 8849 10007 8907 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 4893 9979 4951 9985
rect 4893 9945 4905 9979
rect 4939 9976 4951 9979
rect 5626 9976 5632 9988
rect 4939 9948 5632 9976
rect 4939 9945 4951 9948
rect 4893 9939 4951 9945
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 7466 9936 7472 9988
rect 7524 9976 7530 9988
rect 9508 9976 9536 10152
rect 9766 10140 9772 10152
rect 9824 10140 9830 10192
rect 9950 10189 9956 10192
rect 9944 10180 9956 10189
rect 9911 10152 9956 10180
rect 9944 10143 9956 10152
rect 9950 10140 9956 10143
rect 10008 10140 10014 10192
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 11692 10183 11750 10189
rect 10192 10152 11560 10180
rect 10192 10140 10198 10152
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10226 10112 10232 10124
rect 9723 10084 10232 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10226 10072 10232 10084
rect 10284 10112 10290 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 10284 10084 11437 10112
rect 10284 10072 10290 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11532 10112 11560 10152
rect 11692 10149 11704 10183
rect 11738 10180 11750 10183
rect 12342 10180 12348 10192
rect 11738 10152 12348 10180
rect 11738 10149 11750 10152
rect 11692 10143 11750 10149
rect 12342 10140 12348 10152
rect 12400 10140 12406 10192
rect 12894 10112 12900 10124
rect 11532 10084 12900 10112
rect 11425 10075 11483 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 13446 10112 13452 10124
rect 13407 10084 13452 10112
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12710 10044 12716 10056
rect 12492 10016 12716 10044
rect 12492 10004 12498 10016
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13228 10016 13553 10044
rect 13228 10004 13234 10016
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 14090 10044 14096 10056
rect 13771 10016 14096 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 7524 9948 9536 9976
rect 7524 9936 7530 9948
rect 4062 9908 4068 9920
rect 4023 9880 4068 9908
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9908 5043 9911
rect 7650 9908 7656 9920
rect 5031 9880 7656 9908
rect 5031 9877 5043 9880
rect 4985 9871 5043 9877
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8662 9908 8668 9920
rect 7791 9880 8668 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 10318 9908 10324 9920
rect 9456 9880 10324 9908
rect 9456 9868 9462 9880
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 11054 9908 11060 9920
rect 10967 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9908 11118 9920
rect 12710 9908 12716 9920
rect 11112 9880 12716 9908
rect 11112 9868 11118 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 10410 9704 10416 9716
rect 4028 9676 10416 9704
rect 4028 9664 4034 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 10520 9676 10824 9704
rect 1949 9639 2007 9645
rect 1949 9605 1961 9639
rect 1995 9636 2007 9639
rect 3050 9636 3056 9648
rect 1995 9608 3056 9636
rect 1995 9605 2007 9608
rect 1949 9599 2007 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 4985 9639 5043 9645
rect 4448 9608 4752 9636
rect 2590 9568 2596 9580
rect 2551 9540 2596 9568
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 3510 9568 3516 9580
rect 3471 9540 3516 9568
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 4448 9577 4476 9608
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4614 9568 4620 9580
rect 4575 9540 4620 9568
rect 4433 9531 4491 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 4724 9568 4752 9608
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 8113 9639 8171 9645
rect 5031 9608 7972 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5629 9571 5687 9577
rect 4724 9540 5580 9568
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3418 9500 3424 9512
rect 2740 9472 3424 9500
rect 2740 9460 2746 9472
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5316 9472 5457 9500
rect 5316 9460 5322 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5552 9500 5580 9540
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5810 9568 5816 9580
rect 5675 9540 5816 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 7006 9568 7012 9580
rect 6564 9540 7012 9568
rect 6564 9500 6592 9540
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 7374 9568 7380 9580
rect 7335 9540 7380 9568
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 5552 9472 6592 9500
rect 6641 9503 6699 9509
rect 5445 9463 5503 9469
rect 5644 9444 5672 9472
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 6687 9472 7880 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 3329 9435 3387 9441
rect 3329 9401 3341 9435
rect 3375 9432 3387 9435
rect 3375 9404 4016 9432
rect 3375 9401 3387 9404
rect 3329 9395 3387 9401
rect 2314 9364 2320 9376
rect 2275 9336 2320 9364
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9364 2467 9367
rect 2961 9367 3019 9373
rect 2961 9364 2973 9367
rect 2455 9336 2973 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 2961 9333 2973 9336
rect 3007 9333 3019 9367
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 2961 9327 3019 9333
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3988 9373 4016 9404
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 5166 9432 5172 9444
rect 4212 9404 5172 9432
rect 4212 9392 4218 9404
rect 5166 9392 5172 9404
rect 5224 9432 5230 9444
rect 5224 9404 5479 9432
rect 5224 9392 5230 9404
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9333 4031 9367
rect 3973 9327 4031 9333
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4706 9364 4712 9376
rect 4387 9336 4712 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 5350 9364 5356 9376
rect 5311 9336 5356 9364
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5451 9364 5479 9404
rect 5626 9392 5632 9444
rect 5684 9392 5690 9444
rect 5997 9435 6055 9441
rect 5997 9401 6009 9435
rect 6043 9432 6055 9435
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6043 9404 7205 9432
rect 6043 9401 6055 9404
rect 5997 9395 6055 9401
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7340 9404 7385 9432
rect 7340 9392 7346 9404
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 5451 9336 6469 9364
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 7098 9364 7104 9376
rect 6871 9336 7104 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7852 9373 7880 9472
rect 7944 9432 7972 9608
rect 8113 9605 8125 9639
rect 8159 9636 8171 9639
rect 8294 9636 8300 9648
rect 8159 9608 8300 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 9585 9639 9643 9645
rect 9585 9605 9597 9639
rect 9631 9636 9643 9639
rect 10520 9636 10548 9676
rect 9631 9608 10548 9636
rect 9631 9605 9643 9608
rect 9585 9599 9643 9605
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 10796 9636 10824 9676
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 16758 9704 16764 9716
rect 11112 9676 16764 9704
rect 11112 9664 11118 9676
rect 16758 9664 16764 9676
rect 16816 9664 16822 9716
rect 10652 9608 10697 9636
rect 10796 9608 11284 9636
rect 10652 9596 10658 9608
rect 8662 9568 8668 9580
rect 8623 9540 8668 9568
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10008 9540 10149 9568
rect 10008 9528 10014 9540
rect 10137 9537 10149 9540
rect 10183 9568 10195 9571
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10183 9540 11161 9568
rect 10183 9537 10195 9540
rect 10137 9531 10195 9537
rect 11149 9537 11161 9540
rect 11195 9537 11207 9571
rect 11256 9568 11284 9608
rect 11698 9596 11704 9648
rect 11756 9636 11762 9648
rect 11882 9636 11888 9648
rect 11756 9608 11888 9636
rect 11756 9596 11762 9608
rect 11882 9596 11888 9608
rect 11940 9596 11946 9648
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 12526 9636 12532 9648
rect 12483 9608 12532 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 14277 9639 14335 9645
rect 14277 9636 14289 9639
rect 12768 9608 13032 9636
rect 12768 9596 12774 9608
rect 13004 9577 13032 9608
rect 13648 9608 14289 9636
rect 13648 9580 13676 9608
rect 14277 9605 14289 9608
rect 14323 9605 14335 9639
rect 14277 9599 14335 9605
rect 14461 9639 14519 9645
rect 14461 9605 14473 9639
rect 14507 9636 14519 9639
rect 17954 9636 17960 9648
rect 14507 9608 17960 9636
rect 14507 9605 14519 9608
rect 14461 9599 14519 9605
rect 17954 9596 17960 9608
rect 18012 9596 18018 9648
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 11256 9540 12909 9568
rect 11149 9531 11207 9537
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13630 9528 13636 9580
rect 13688 9528 13694 9580
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 9490 9500 9496 9512
rect 8067 9472 9496 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10505 9503 10563 9509
rect 10505 9500 10517 9503
rect 9732 9472 10517 9500
rect 9732 9460 9738 9472
rect 10505 9469 10517 9472
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 10652 9472 12817 9500
rect 10652 9460 10658 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 12805 9463 12863 9469
rect 12912 9472 13829 9500
rect 10870 9432 10876 9444
rect 7944 9404 10876 9432
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 10965 9435 11023 9441
rect 10965 9401 10977 9435
rect 11011 9432 11023 9435
rect 11609 9435 11667 9441
rect 11609 9432 11621 9435
rect 11011 9404 11621 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 11609 9401 11621 9404
rect 11655 9401 11667 9435
rect 11609 9395 11667 9401
rect 7837 9367 7895 9373
rect 7837 9333 7849 9367
rect 7883 9364 7895 9367
rect 8294 9364 8300 9376
rect 7883 9336 8300 9364
rect 7883 9333 7895 9336
rect 7837 9327 7895 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 8573 9367 8631 9373
rect 8573 9333 8585 9367
rect 8619 9364 8631 9367
rect 8754 9364 8760 9376
rect 8619 9336 8760 9364
rect 8619 9333 8631 9336
rect 8573 9327 8631 9333
rect 8754 9324 8760 9336
rect 8812 9324 8818 9376
rect 9950 9364 9956 9376
rect 9911 9336 9956 9364
rect 9950 9324 9956 9336
rect 10008 9324 10014 9376
rect 10045 9367 10103 9373
rect 10045 9333 10057 9367
rect 10091 9364 10103 9367
rect 10134 9364 10140 9376
rect 10091 9336 10140 9364
rect 10091 9333 10103 9336
rect 10045 9327 10103 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10505 9367 10563 9373
rect 10505 9333 10517 9367
rect 10551 9364 10563 9367
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 10551 9336 11069 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11057 9327 11115 9333
rect 11514 9324 11520 9376
rect 11572 9364 11578 9376
rect 12912 9364 12940 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 14016 9500 14044 9531
rect 14090 9528 14096 9580
rect 14148 9568 14154 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14148 9540 15025 9568
rect 14148 9528 14154 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15013 9531 15071 9537
rect 14182 9500 14188 9512
rect 14016 9472 14188 9500
rect 13817 9463 13875 9469
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 15102 9500 15108 9512
rect 14323 9472 15108 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 15102 9460 15108 9472
rect 15160 9460 15166 9512
rect 14829 9435 14887 9441
rect 14829 9432 14841 9435
rect 13464 9404 14841 9432
rect 13464 9373 13492 9404
rect 14829 9401 14841 9404
rect 14875 9401 14887 9435
rect 14829 9395 14887 9401
rect 11572 9336 12940 9364
rect 13449 9367 13507 9373
rect 11572 9324 11578 9336
rect 13449 9333 13461 9367
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 13964 9336 14009 9364
rect 13964 9324 13970 9336
rect 14550 9324 14556 9376
rect 14608 9364 14614 9376
rect 14921 9367 14979 9373
rect 14921 9364 14933 9367
rect 14608 9336 14933 9364
rect 14608 9324 14614 9336
rect 14921 9333 14933 9336
rect 14967 9333 14979 9367
rect 14921 9327 14979 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3476 9132 4077 9160
rect 3476 9120 3482 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 5534 9160 5540 9172
rect 4571 9132 5540 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 5534 9120 5540 9132
rect 5592 9160 5598 9172
rect 6730 9160 6736 9172
rect 5592 9132 6736 9160
rect 5592 9120 5598 9132
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 8297 9163 8355 9169
rect 8297 9160 8309 9163
rect 6871 9132 8309 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 8297 9129 8309 9132
rect 8343 9129 8355 9163
rect 8297 9123 8355 9129
rect 9217 9163 9275 9169
rect 9217 9129 9229 9163
rect 9263 9160 9275 9163
rect 9950 9160 9956 9172
rect 9263 9132 9956 9160
rect 9263 9129 9275 9132
rect 9217 9123 9275 9129
rect 9950 9120 9956 9132
rect 10008 9160 10014 9172
rect 10137 9163 10195 9169
rect 10137 9160 10149 9163
rect 10008 9132 10149 9160
rect 10008 9120 10014 9132
rect 10137 9129 10149 9132
rect 10183 9129 10195 9163
rect 10137 9123 10195 9129
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 11054 9160 11060 9172
rect 10468 9132 11060 9160
rect 10468 9120 10474 9132
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 11664 9132 12020 9160
rect 11664 9120 11670 9132
rect 2308 9095 2366 9101
rect 2308 9061 2320 9095
rect 2354 9092 2366 9095
rect 2498 9092 2504 9104
rect 2354 9064 2504 9092
rect 2354 9061 2366 9064
rect 2308 9055 2366 9061
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 7098 9052 7104 9104
rect 7156 9092 7162 9104
rect 8205 9095 8263 9101
rect 8205 9092 8217 9095
rect 7156 9064 8217 9092
rect 7156 9052 7162 9064
rect 8205 9061 8217 9064
rect 8251 9061 8263 9095
rect 8205 9055 8263 9061
rect 8849 9095 8907 9101
rect 8849 9061 8861 9095
rect 8895 9092 8907 9095
rect 11514 9092 11520 9104
rect 8895 9064 11520 9092
rect 8895 9061 8907 9064
rect 8849 9055 8907 9061
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 11992 9092 12020 9132
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 13173 9163 13231 9169
rect 13173 9160 13185 9163
rect 12400 9132 13185 9160
rect 12400 9120 12406 9132
rect 13173 9129 13185 9132
rect 13219 9129 13231 9163
rect 13173 9123 13231 9129
rect 13725 9163 13783 9169
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 13906 9160 13912 9172
rect 13771 9132 13912 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14366 9160 14372 9172
rect 14139 9132 14372 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 12069 9095 12127 9101
rect 12069 9092 12081 9095
rect 11992 9064 12081 9092
rect 12069 9061 12081 9064
rect 12115 9061 12127 9095
rect 13081 9095 13139 9101
rect 13081 9092 13093 9095
rect 12069 9055 12127 9061
rect 12176 9064 13093 9092
rect 2516 9024 2544 9052
rect 3881 9027 3939 9033
rect 2516 8996 3832 9024
rect 1578 8956 1584 8968
rect 1539 8928 1584 8956
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 2038 8956 2044 8968
rect 1951 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2056 8820 2084 8916
rect 3804 8888 3832 8996
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4154 9024 4160 9036
rect 3927 8996 4160 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4430 9024 4436 9036
rect 4391 8996 4436 9024
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 5074 8984 5080 9036
rect 5132 9024 5138 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 5132 8996 5181 9024
rect 5132 8984 5138 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 5258 8984 5264 9036
rect 5316 8984 5322 9036
rect 5436 9027 5494 9033
rect 5436 8993 5448 9027
rect 5482 9024 5494 9027
rect 5482 8996 6684 9024
rect 5482 8993 5494 8996
rect 5436 8987 5494 8993
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 4672 8928 4765 8956
rect 4672 8916 4678 8928
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 5276 8956 5304 8984
rect 4856 8928 5304 8956
rect 4856 8916 4862 8928
rect 4632 8888 4660 8916
rect 3252 8860 3740 8888
rect 3804 8860 4660 8888
rect 6656 8888 6684 8996
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 7064 8996 7205 9024
rect 7064 8984 7070 8996
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8352 8996 9505 9024
rect 8352 8984 8358 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9732 8996 10057 9024
rect 9732 8984 9738 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 12176 9024 12204 9064
rect 13081 9061 13093 9064
rect 13127 9061 13139 9095
rect 13081 9055 13139 9061
rect 10045 8987 10103 8993
rect 12084 8996 12204 9024
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 8389 8959 8447 8965
rect 7432 8928 7477 8956
rect 7432 8916 7438 8928
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 7392 8888 7420 8916
rect 8404 8888 8432 8919
rect 8662 8916 8668 8968
rect 8720 8956 8726 8968
rect 10229 8959 10287 8965
rect 8720 8928 9996 8956
rect 8720 8916 8726 8928
rect 6656 8860 7420 8888
rect 7484 8860 8432 8888
rect 9309 8891 9367 8897
rect 3252 8820 3280 8860
rect 3418 8820 3424 8832
rect 2056 8792 3280 8820
rect 3379 8792 3424 8820
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 3712 8829 3740 8860
rect 3697 8823 3755 8829
rect 3697 8789 3709 8823
rect 3743 8820 3755 8823
rect 5074 8820 5080 8832
rect 3743 8792 5080 8820
rect 3743 8789 3755 8792
rect 3697 8783 3755 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 6549 8823 6607 8829
rect 6549 8789 6561 8823
rect 6595 8820 6607 8823
rect 6638 8820 6644 8832
rect 6595 8792 6644 8820
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 6638 8780 6644 8792
rect 6696 8820 6702 8832
rect 7484 8820 7512 8860
rect 9309 8857 9321 8891
rect 9355 8888 9367 8891
rect 9858 8888 9864 8900
rect 9355 8860 9864 8888
rect 9355 8857 9367 8860
rect 9309 8851 9367 8857
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 6696 8792 7512 8820
rect 6696 8780 6702 8792
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7708 8792 7849 8820
rect 7708 8780 7714 8792
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 7926 8780 7932 8832
rect 7984 8820 7990 8832
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 7984 8792 9229 8820
rect 7984 8780 7990 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 9766 8820 9772 8832
rect 9723 8792 9772 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 9968 8820 9996 8928
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 10042 8848 10048 8900
rect 10100 8888 10106 8900
rect 10244 8888 10272 8919
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 10560 8928 11161 8956
rect 10560 8916 10566 8928
rect 11149 8925 11161 8928
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12084 8956 12112 8996
rect 11296 8928 11341 8956
rect 11716 8928 12112 8956
rect 12161 8959 12219 8965
rect 11296 8916 11302 8928
rect 10100 8860 10272 8888
rect 10689 8891 10747 8897
rect 10100 8848 10106 8860
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 11422 8888 11428 8900
rect 10735 8860 11428 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 11422 8848 11428 8860
rect 11480 8848 11486 8900
rect 11716 8897 11744 8928
rect 12161 8925 12173 8959
rect 12207 8925 12219 8959
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 12161 8919 12219 8925
rect 11701 8891 11759 8897
rect 11701 8857 11713 8891
rect 11747 8857 11759 8891
rect 12176 8888 12204 8919
rect 12342 8916 12348 8928
rect 12400 8956 12406 8968
rect 13078 8956 13084 8968
rect 12400 8928 13084 8956
rect 12400 8916 12406 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13814 8916 13820 8968
rect 13872 8956 13878 8968
rect 14185 8959 14243 8965
rect 14185 8956 14197 8959
rect 13872 8928 14197 8956
rect 13872 8916 13878 8928
rect 14185 8925 14197 8928
rect 14231 8925 14243 8959
rect 14185 8919 14243 8925
rect 14274 8916 14280 8968
rect 14332 8956 14338 8968
rect 14332 8928 14377 8956
rect 14332 8916 14338 8928
rect 12434 8888 12440 8900
rect 12176 8860 12440 8888
rect 11701 8851 11759 8857
rect 12434 8848 12440 8860
rect 12492 8848 12498 8900
rect 12618 8888 12624 8900
rect 12531 8860 12624 8888
rect 12544 8820 12572 8860
rect 12618 8848 12624 8860
rect 12676 8888 12682 8900
rect 13446 8888 13452 8900
rect 12676 8860 13452 8888
rect 12676 8848 12682 8860
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 12710 8820 12716 8832
rect 9968 8792 12572 8820
rect 12671 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2038 8616 2044 8628
rect 1412 8588 2044 8616
rect 1412 8489 1440 8588
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 3053 8619 3111 8625
rect 3053 8616 3065 8619
rect 2372 8588 3065 8616
rect 2372 8576 2378 8588
rect 3053 8585 3065 8588
rect 3099 8585 3111 8619
rect 3053 8579 3111 8585
rect 3970 8576 3976 8628
rect 4028 8616 4034 8628
rect 6457 8619 6515 8625
rect 4028 8588 6408 8616
rect 4028 8576 4034 8588
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 2777 8551 2835 8557
rect 2777 8548 2789 8551
rect 2648 8520 2789 8548
rect 2648 8508 2654 8520
rect 2777 8517 2789 8520
rect 2823 8517 2835 8551
rect 2777 8511 2835 8517
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8449 1455 8483
rect 3418 8480 3424 8492
rect 1397 8443 1455 8449
rect 3068 8452 3424 8480
rect 1664 8415 1722 8421
rect 1664 8381 1676 8415
rect 1710 8412 1722 8415
rect 3068 8412 3096 8452
rect 3418 8440 3424 8452
rect 3476 8480 3482 8492
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 3476 8452 3617 8480
rect 3476 8440 3482 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4525 8483 4583 8489
rect 4525 8480 4537 8483
rect 4212 8452 4537 8480
rect 4212 8440 4218 8452
rect 4525 8449 4537 8452
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 4890 8480 4896 8492
rect 4755 8452 4896 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 5074 8480 5080 8492
rect 5035 8452 5080 8480
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 6380 8480 6408 8588
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 7374 8616 7380 8628
rect 6503 8588 7380 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 10134 8616 10140 8628
rect 10047 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8616 10198 8628
rect 14090 8616 14096 8628
rect 10192 8588 14096 8616
rect 10192 8576 10198 8588
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14550 8616 14556 8628
rect 14507 8588 14556 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 12066 8548 12072 8560
rect 12027 8520 12072 8548
rect 12066 8508 12072 8520
rect 12124 8508 12130 8560
rect 12253 8551 12311 8557
rect 12253 8517 12265 8551
rect 12299 8548 12311 8551
rect 12342 8548 12348 8560
rect 12299 8520 12348 8548
rect 12299 8517 12311 8520
rect 12253 8511 12311 8517
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 13449 8551 13507 8557
rect 13004 8520 13400 8548
rect 6380 8452 7236 8480
rect 1710 8384 3096 8412
rect 3513 8415 3571 8421
rect 1710 8381 1722 8384
rect 1664 8375 1722 8381
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 4062 8412 4068 8424
rect 3559 8384 4068 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7208 8412 7236 8452
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 13004 8480 13032 8520
rect 11940 8452 13032 8480
rect 13081 8483 13139 8489
rect 11940 8440 11946 8452
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13262 8480 13268 8492
rect 13127 8452 13268 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 13372 8480 13400 8520
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 13495 8520 14872 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13372 8452 13921 8480
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8480 14151 8483
rect 14274 8480 14280 8492
rect 14139 8452 14280 8480
rect 14139 8449 14151 8452
rect 14093 8443 14151 8449
rect 14274 8440 14280 8452
rect 14332 8440 14338 8492
rect 7926 8412 7932 8424
rect 7208 8384 7932 8412
rect 7101 8375 7159 8381
rect 5344 8347 5402 8353
rect 5344 8313 5356 8347
rect 5390 8344 5402 8347
rect 5534 8344 5540 8356
rect 5390 8316 5540 8344
rect 5390 8313 5402 8316
rect 5344 8307 5402 8313
rect 5534 8304 5540 8316
rect 5592 8304 5598 8356
rect 7116 8344 7144 8375
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8036 8384 8769 8412
rect 7374 8353 7380 8356
rect 7368 8344 7380 8353
rect 7116 8316 7236 8344
rect 7335 8316 7380 8344
rect 3418 8276 3424 8288
rect 3379 8248 3424 8276
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 4062 8276 4068 8288
rect 4023 8248 4068 8276
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4433 8279 4491 8285
rect 4433 8276 4445 8279
rect 4212 8248 4445 8276
rect 4212 8236 4218 8248
rect 4433 8245 4445 8248
rect 4479 8245 4491 8279
rect 4433 8239 4491 8245
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5166 8276 5172 8288
rect 4764 8248 5172 8276
rect 4764 8236 4770 8248
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 7208 8276 7236 8316
rect 7368 8307 7380 8316
rect 7374 8304 7380 8307
rect 7432 8304 7438 8356
rect 8036 8344 8064 8384
rect 8757 8381 8769 8384
rect 8803 8412 8815 8415
rect 10226 8412 10232 8424
rect 8803 8384 10232 8412
rect 8803 8381 8815 8384
rect 8757 8375 8815 8381
rect 10226 8372 10232 8384
rect 10284 8412 10290 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10284 8384 10701 8412
rect 10284 8372 10290 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 14182 8412 14188 8424
rect 10689 8375 10747 8381
rect 10796 8384 14188 8412
rect 9024 8347 9082 8353
rect 9024 8344 9036 8347
rect 7484 8316 8064 8344
rect 8496 8316 9036 8344
rect 7484 8276 7512 8316
rect 8496 8285 8524 8316
rect 9024 8313 9036 8316
rect 9070 8344 9082 8347
rect 10796 8344 10824 8384
rect 14182 8372 14188 8384
rect 14240 8412 14246 8424
rect 14844 8421 14872 8520
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14936 8452 15025 8480
rect 14829 8415 14887 8421
rect 14240 8384 14780 8412
rect 14240 8372 14246 8384
rect 9070 8316 10824 8344
rect 9070 8313 9082 8316
rect 9024 8307 9082 8313
rect 10870 8304 10876 8356
rect 10928 8353 10934 8356
rect 10928 8347 10992 8353
rect 10928 8313 10946 8347
rect 10980 8344 10992 8347
rect 11146 8344 11152 8356
rect 10980 8316 11152 8344
rect 10980 8313 10992 8316
rect 10928 8307 10992 8313
rect 10928 8304 10934 8307
rect 11146 8304 11152 8316
rect 11204 8344 11210 8356
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 11204 8316 12265 8344
rect 11204 8304 11210 8316
rect 12253 8313 12265 8316
rect 12299 8313 12311 8347
rect 12802 8344 12808 8356
rect 12763 8316 12808 8344
rect 12253 8307 12311 8313
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 14752 8344 14780 8384
rect 14829 8381 14841 8415
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 14936 8344 14964 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 13780 8316 14412 8344
rect 14752 8316 14964 8344
rect 13780 8304 13786 8316
rect 7208 8248 7512 8276
rect 8481 8279 8539 8285
rect 8481 8245 8493 8279
rect 8527 8245 8539 8279
rect 8481 8239 8539 8245
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 12158 8276 12164 8288
rect 9180 8248 12164 8276
rect 9180 8236 9186 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 12492 8248 12537 8276
rect 12492 8236 12498 8248
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13817 8279 13875 8285
rect 12952 8248 12997 8276
rect 12952 8236 12958 8248
rect 13817 8245 13829 8279
rect 13863 8276 13875 8279
rect 13906 8276 13912 8288
rect 13863 8248 13912 8276
rect 13863 8245 13875 8248
rect 13817 8239 13875 8245
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 14384 8276 14412 8316
rect 14921 8279 14979 8285
rect 14921 8276 14933 8279
rect 14384 8248 14933 8276
rect 14921 8245 14933 8248
rect 14967 8245 14979 8279
rect 14921 8239 14979 8245
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 1636 8044 2329 8072
rect 1636 8032 1642 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 3467 8044 4261 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 4982 8072 4988 8084
rect 4396 8044 4988 8072
rect 4396 8032 4402 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 7193 8075 7251 8081
rect 7193 8072 7205 8075
rect 5592 8044 7205 8072
rect 5592 8032 5598 8044
rect 7193 8041 7205 8044
rect 7239 8041 7251 8075
rect 7193 8035 7251 8041
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7340 8044 7481 8072
rect 7340 8032 7346 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7708 8044 7849 8072
rect 7708 8032 7714 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 8527 8044 10456 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 3329 8007 3387 8013
rect 3329 7973 3341 8007
rect 3375 8004 3387 8007
rect 4062 8004 4068 8016
rect 3375 7976 4068 8004
rect 3375 7973 3387 7976
rect 3329 7967 3387 7973
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 4709 8007 4767 8013
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 4798 8004 4804 8016
rect 4755 7976 4804 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 6733 8007 6791 8013
rect 6733 7973 6745 8007
rect 6779 8004 6791 8007
rect 8294 8004 8300 8016
rect 6779 7976 8300 8004
rect 6779 7973 6791 7976
rect 6733 7967 6791 7973
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 8444 7976 8953 8004
rect 8444 7964 8450 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 9122 8004 9128 8016
rect 8941 7967 8999 7973
rect 9048 7976 9128 8004
rect 2409 7939 2467 7945
rect 2409 7905 2421 7939
rect 2455 7936 2467 7939
rect 2455 7908 3924 7936
rect 2455 7905 2467 7908
rect 2409 7899 2467 7905
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 3605 7871 3663 7877
rect 2556 7840 2601 7868
rect 2556 7828 2562 7840
rect 3605 7837 3617 7871
rect 3651 7837 3663 7871
rect 3896 7868 3924 7908
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 4617 7939 4675 7945
rect 4617 7936 4629 7939
rect 4028 7908 4629 7936
rect 4028 7896 4034 7908
rect 4617 7905 4629 7908
rect 4663 7936 4675 7939
rect 5350 7936 5356 7948
rect 4663 7908 5356 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7936 5963 7939
rect 6362 7936 6368 7948
rect 5951 7908 6368 7936
rect 5951 7905 5963 7908
rect 5905 7899 5963 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 6638 7936 6644 7948
rect 6599 7908 6644 7936
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7650 7936 7656 7948
rect 7156 7908 7656 7936
rect 7156 7896 7162 7908
rect 7650 7896 7656 7908
rect 7708 7896 7714 7948
rect 8849 7939 8907 7945
rect 7760 7908 8064 7936
rect 4338 7868 4344 7880
rect 3896 7840 4344 7868
rect 3605 7831 3663 7837
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7800 2007 7803
rect 3418 7800 3424 7812
rect 1995 7772 3424 7800
rect 1995 7769 2007 7772
rect 1949 7763 2007 7769
rect 3418 7760 3424 7772
rect 3476 7760 3482 7812
rect 2958 7732 2964 7744
rect 2919 7704 2964 7732
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3620 7732 3648 7831
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4890 7868 4896 7880
rect 4803 7840 4896 7868
rect 4890 7828 4896 7840
rect 4948 7868 4954 7880
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 4948 7840 6101 7868
rect 4948 7828 4954 7840
rect 6089 7837 6101 7840
rect 6135 7868 6147 7871
rect 6178 7868 6184 7880
rect 6135 7840 6184 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6788 7840 6837 7868
rect 6788 7828 6794 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 7760 7868 7788 7908
rect 7926 7868 7932 7880
rect 7239 7840 7788 7868
rect 7887 7840 7932 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8036 7877 8064 7908
rect 8849 7905 8861 7939
rect 8895 7936 8907 7939
rect 9048 7936 9076 7976
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 9944 8007 10002 8013
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 10134 8004 10140 8016
rect 9990 7976 10140 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10428 8004 10456 8044
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10870 8072 10876 8084
rect 10652 8044 10876 8072
rect 10652 8032 10658 8044
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 11333 8075 11391 8081
rect 11333 8041 11345 8075
rect 11379 8072 11391 8075
rect 11606 8072 11612 8084
rect 11379 8044 11612 8072
rect 11379 8041 11391 8044
rect 11333 8035 11391 8041
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 14458 8072 14464 8084
rect 11716 8044 14464 8072
rect 11716 8004 11744 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 13814 8004 13820 8016
rect 10428 7976 11744 8004
rect 11900 7976 13820 8004
rect 9674 7936 9680 7948
rect 8895 7908 9076 7936
rect 9587 7908 9680 7936
rect 8895 7905 8907 7908
rect 8849 7899 8907 7905
rect 9674 7896 9680 7908
rect 9732 7936 9738 7948
rect 10226 7936 10232 7948
rect 9732 7908 10232 7936
rect 9732 7896 9738 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11606 7896 11612 7948
rect 11664 7936 11670 7948
rect 11793 7939 11851 7945
rect 11793 7936 11805 7939
rect 11664 7908 11805 7936
rect 11664 7896 11670 7908
rect 11793 7905 11805 7908
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7868 9183 7871
rect 9306 7868 9312 7880
rect 9171 7840 9312 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 11900 7868 11928 7976
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 12066 7945 12072 7948
rect 12060 7899 12072 7945
rect 12124 7936 12130 7948
rect 13722 7945 13728 7948
rect 13716 7936 13728 7945
rect 12124 7908 12160 7936
rect 13683 7908 13728 7936
rect 12066 7896 12072 7899
rect 12124 7896 12130 7908
rect 13716 7899 13728 7908
rect 13722 7896 13728 7899
rect 13780 7896 13786 7948
rect 13446 7868 13452 7880
rect 10888 7840 11928 7868
rect 13407 7840 13452 7868
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 4120 7772 8064 7800
rect 4120 7760 4126 7772
rect 4706 7732 4712 7744
rect 3620 7704 4712 7732
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 5442 7732 5448 7744
rect 5403 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 6270 7732 6276 7744
rect 6231 7704 6276 7732
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7377 7735 7435 7741
rect 7377 7701 7389 7735
rect 7423 7732 7435 7735
rect 7558 7732 7564 7744
rect 7423 7704 7564 7732
rect 7423 7701 7435 7704
rect 7377 7695 7435 7701
rect 7558 7692 7564 7704
rect 7616 7732 7622 7744
rect 7926 7732 7932 7744
rect 7616 7704 7932 7732
rect 7616 7692 7622 7704
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8036 7732 8064 7772
rect 10888 7732 10916 7840
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 11054 7732 11060 7744
rect 8036 7704 10916 7732
rect 11015 7704 11060 7732
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 12032 7704 13185 7732
rect 12032 7692 12038 7704
rect 13173 7701 13185 7704
rect 13219 7732 13231 7735
rect 13722 7732 13728 7744
rect 13219 7704 13728 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14240 7704 14841 7732
rect 14240 7692 14246 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 14829 7695 14887 7701
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 5810 7528 5816 7540
rect 3292 7500 5816 7528
rect 3292 7488 3298 7500
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7248 7500 7849 7528
rect 7248 7488 7254 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 12437 7531 12495 7537
rect 7837 7491 7895 7497
rect 8864 7500 12388 7528
rect 6270 7420 6276 7472
rect 6328 7460 6334 7472
rect 6328 7432 7512 7460
rect 6328 7420 6334 7432
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3513 7395 3571 7401
rect 3513 7392 3525 7395
rect 2924 7364 3525 7392
rect 2924 7352 2930 7364
rect 3513 7361 3525 7364
rect 3559 7361 3571 7395
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 3513 7355 3571 7361
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 1394 7284 1400 7336
rect 1452 7324 1458 7336
rect 2317 7327 2375 7333
rect 2317 7324 2329 7327
rect 1452 7296 2329 7324
rect 1452 7284 1458 7296
rect 2317 7293 2329 7296
rect 2363 7293 2375 7327
rect 2317 7287 2375 7293
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 4617 7327 4675 7333
rect 2464 7296 2509 7324
rect 2464 7284 2470 7296
rect 4617 7293 4629 7327
rect 4663 7293 4675 7327
rect 4617 7287 4675 7293
rect 4632 7256 4660 7287
rect 4706 7284 4712 7336
rect 4764 7324 4770 7336
rect 4873 7327 4931 7333
rect 4873 7324 4885 7327
rect 4764 7296 4885 7324
rect 4764 7284 4770 7296
rect 4873 7293 4885 7296
rect 4919 7324 4931 7327
rect 4919 7296 5396 7324
rect 4919 7293 4931 7296
rect 4873 7287 4931 7293
rect 5074 7256 5080 7268
rect 4632 7228 5080 7256
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 5368 7256 5396 7296
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 5500 7296 7205 7324
rect 5500 7284 5506 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 7392 7256 7420 7355
rect 7484 7324 7512 7432
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 8864 7401 8892 7500
rect 10597 7463 10655 7469
rect 10597 7429 10609 7463
rect 10643 7460 10655 7463
rect 11606 7460 11612 7472
rect 10643 7432 11612 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 12360 7460 12388 7500
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 12894 7528 12900 7540
rect 12483 7500 12900 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13449 7463 13507 7469
rect 11808 7432 12296 7460
rect 12360 7432 13308 7460
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 7708 7364 8401 7392
rect 7708 7352 7714 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7361 8907 7395
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 8849 7355 8907 7361
rect 8956 7364 10057 7392
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 7484 7296 8217 7324
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8956 7324 8984 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10226 7392 10232 7404
rect 10187 7364 10232 7392
rect 10045 7355 10103 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 11808 7401 11836 7432
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11974 7392 11980 7404
rect 11935 7364 11980 7392
rect 11793 7355 11851 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 8205 7287 8263 7293
rect 8312 7296 8984 7324
rect 5368 7228 7420 7256
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 8312 7256 8340 7296
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 9916 7296 10793 7324
rect 9916 7284 9922 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 12268 7324 12296 7432
rect 13078 7392 13084 7404
rect 13039 7364 13084 7392
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 12434 7324 12440 7336
rect 11747 7296 12112 7324
rect 12268 7296 12440 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 7800 7228 8340 7256
rect 9953 7259 10011 7265
rect 7800 7216 7806 7228
rect 9953 7225 9965 7259
rect 9999 7256 10011 7259
rect 10318 7256 10324 7268
rect 9999 7228 10324 7256
rect 9999 7225 10011 7228
rect 9953 7219 10011 7225
rect 10318 7216 10324 7228
rect 10376 7216 10382 7268
rect 12084 7256 12112 7296
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 13280 7324 13308 7432
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 15746 7460 15752 7472
rect 13495 7432 15752 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 13722 7392 13728 7404
rect 13596 7364 13728 7392
rect 13596 7352 13602 7364
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 14090 7392 14096 7404
rect 14003 7364 14096 7392
rect 14090 7352 14096 7364
rect 14148 7392 14154 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 14148 7364 15117 7392
rect 14148 7352 14154 7364
rect 15105 7361 15117 7364
rect 15151 7392 15163 7395
rect 16942 7392 16948 7404
rect 15151 7364 16948 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 13280 7296 14841 7324
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 12710 7256 12716 7268
rect 11348 7228 11928 7256
rect 12084 7228 12716 7256
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 2961 7191 3019 7197
rect 2961 7157 2973 7191
rect 3007 7188 3019 7191
rect 3142 7188 3148 7200
rect 3007 7160 3148 7188
rect 3007 7157 3019 7160
rect 2961 7151 3019 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3326 7188 3332 7200
rect 3287 7160 3332 7188
rect 3326 7148 3332 7160
rect 3384 7148 3390 7200
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 5994 7188 6000 7200
rect 3476 7160 3521 7188
rect 5955 7160 6000 7188
rect 3476 7148 3482 7160
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6825 7191 6883 7197
rect 6825 7157 6837 7191
rect 6871 7188 6883 7191
rect 7190 7188 7196 7200
rect 6871 7160 7196 7188
rect 6871 7157 6883 7160
rect 6825 7151 6883 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7282 7148 7288 7200
rect 7340 7188 7346 7200
rect 8294 7188 8300 7200
rect 7340 7160 7385 7188
rect 8255 7160 8300 7188
rect 7340 7148 7346 7160
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7188 9643 7191
rect 10134 7188 10140 7200
rect 9631 7160 10140 7188
rect 9631 7157 9643 7160
rect 9585 7151 9643 7157
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 11348 7197 11376 7228
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7157 11391 7191
rect 11900 7188 11928 7228
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 12805 7259 12863 7265
rect 12805 7225 12817 7259
rect 12851 7256 12863 7259
rect 12986 7256 12992 7268
rect 12851 7228 12992 7256
rect 12851 7225 12863 7228
rect 12805 7219 12863 7225
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 13814 7256 13820 7268
rect 13775 7228 13820 7256
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14366 7216 14372 7268
rect 14424 7256 14430 7268
rect 14921 7259 14979 7265
rect 14921 7256 14933 7259
rect 14424 7228 14933 7256
rect 14424 7216 14430 7228
rect 14921 7225 14933 7228
rect 14967 7225 14979 7259
rect 14921 7219 14979 7225
rect 12526 7188 12532 7200
rect 11900 7160 12532 7188
rect 11333 7151 11391 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12894 7188 12900 7200
rect 12807 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7188 12958 7200
rect 13354 7188 13360 7200
rect 12952 7160 13360 7188
rect 12952 7148 12958 7160
rect 13354 7148 13360 7160
rect 13412 7148 13418 7200
rect 13906 7188 13912 7200
rect 13867 7160 13912 7188
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14458 7188 14464 7200
rect 14419 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 3016 6956 7941 6984
rect 3016 6944 3022 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 9033 6987 9091 6993
rect 9033 6953 9045 6987
rect 9079 6984 9091 6987
rect 9582 6984 9588 6996
rect 9079 6956 9588 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 13078 6984 13084 6996
rect 13039 6956 13084 6984
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 14274 6984 14280 6996
rect 13771 6956 14280 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 14516 6956 15669 6984
rect 14516 6944 14522 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 1940 6919 1998 6925
rect 1940 6885 1952 6919
rect 1986 6916 1998 6919
rect 2130 6916 2136 6928
rect 1986 6888 2136 6916
rect 1986 6885 1998 6888
rect 1940 6879 1998 6885
rect 2130 6876 2136 6888
rect 2188 6876 2194 6928
rect 2682 6876 2688 6928
rect 2740 6876 2746 6928
rect 4332 6919 4390 6925
rect 4332 6885 4344 6919
rect 4378 6916 4390 6919
rect 4890 6916 4896 6928
rect 4378 6888 4896 6916
rect 4378 6885 4390 6888
rect 4332 6879 4390 6885
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 6362 6916 6368 6928
rect 5960 6888 6368 6916
rect 5960 6876 5966 6888
rect 6362 6876 6368 6888
rect 6420 6916 6426 6928
rect 8941 6919 8999 6925
rect 8941 6916 8953 6919
rect 6420 6888 8953 6916
rect 6420 6876 6426 6888
rect 8941 6885 8953 6888
rect 8987 6885 8999 6919
rect 10042 6916 10048 6928
rect 8941 6879 8999 6885
rect 9039 6888 10048 6916
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 1762 6848 1768 6860
rect 1719 6820 1768 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2700 6848 2728 6876
rect 2958 6848 2964 6860
rect 2700 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6808 3022 6860
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 4111 6820 5396 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 5368 6792 5396 6820
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6172 6851 6230 6857
rect 6172 6848 6184 6851
rect 6052 6820 6184 6848
rect 6052 6808 6058 6820
rect 6172 6817 6184 6820
rect 6218 6848 6230 6851
rect 7377 6851 7435 6857
rect 6218 6820 6960 6848
rect 6218 6817 6230 6820
rect 6172 6811 6230 6817
rect 2682 6740 2688 6792
rect 2740 6780 2746 6792
rect 3329 6783 3387 6789
rect 3329 6780 3341 6783
rect 2740 6752 3341 6780
rect 2740 6740 2746 6752
rect 3329 6749 3341 6752
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5408 6752 5917 6780
rect 5408 6740 5414 6752
rect 5905 6749 5917 6752
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 2866 6672 2872 6724
rect 2924 6712 2930 6724
rect 3053 6715 3111 6721
rect 3053 6712 3065 6715
rect 2924 6684 3065 6712
rect 2924 6672 2930 6684
rect 3053 6681 3065 6684
rect 3099 6681 3111 6715
rect 6932 6712 6960 6820
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 9039 6848 9067 6888
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 10962 6916 10968 6928
rect 10744 6888 10968 6916
rect 10744 6876 10750 6888
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11054 6876 11060 6928
rect 11112 6916 11118 6928
rect 12342 6916 12348 6928
rect 11112 6888 12348 6916
rect 11112 6876 11118 6888
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 13354 6876 13360 6928
rect 13412 6916 13418 6928
rect 16574 6916 16580 6928
rect 13412 6888 16580 6916
rect 13412 6876 13418 6888
rect 16574 6876 16580 6888
rect 16632 6876 16638 6928
rect 9674 6848 9680 6860
rect 7423 6820 9067 6848
rect 9635 6820 9680 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 9674 6808 9680 6820
rect 9732 6808 9738 6860
rect 9944 6851 10002 6857
rect 9944 6817 9956 6851
rect 9990 6848 10002 6851
rect 11072 6848 11100 6876
rect 9990 6820 11100 6848
rect 9990 6817 10002 6820
rect 9944 6811 10002 6817
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 11968 6851 12026 6857
rect 11968 6848 11980 6851
rect 11204 6820 11980 6848
rect 11204 6808 11210 6820
rect 11968 6817 11980 6820
rect 12014 6848 12026 6851
rect 12894 6848 12900 6860
rect 12014 6820 12900 6848
rect 12014 6817 12026 6820
rect 11968 6811 12026 6817
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13780 6820 13829 6848
rect 13780 6808 13786 6820
rect 13817 6817 13829 6820
rect 13863 6848 13875 6851
rect 15010 6848 15016 6860
rect 13863 6820 15016 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15746 6848 15752 6860
rect 15707 6820 15752 6848
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7248 6752 8033 6780
rect 7248 6740 7254 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 8128 6712 8156 6743
rect 6932 6684 8156 6712
rect 3053 6675 3111 6681
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 4764 6616 5457 6644
rect 4764 6604 4770 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7374 6644 7380 6656
rect 7331 6616 7380 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7558 6644 7564 6656
rect 7519 6616 7564 6644
rect 7558 6604 7564 6616
rect 7616 6604 7622 6656
rect 8570 6644 8576 6656
rect 8531 6616 8576 6644
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 9232 6644 9260 6743
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11664 6752 11713 6780
rect 11664 6740 11670 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13262 6780 13268 6792
rect 13044 6752 13268 6780
rect 13044 6740 13050 6752
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 10686 6672 10692 6724
rect 10744 6712 10750 6724
rect 11054 6712 11060 6724
rect 10744 6684 11060 6712
rect 10744 6672 10750 6684
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 13357 6715 13415 6721
rect 13357 6681 13369 6715
rect 13403 6712 13415 6715
rect 13814 6712 13820 6724
rect 13403 6684 13820 6712
rect 13403 6681 13415 6684
rect 13357 6675 13415 6681
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 10594 6644 10600 6656
rect 9232 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 13262 6644 13268 6656
rect 12400 6616 13268 6644
rect 12400 6604 12406 6616
rect 13262 6604 13268 6616
rect 13320 6644 13326 6656
rect 13924 6644 13952 6743
rect 14550 6740 14556 6792
rect 14608 6780 14614 6792
rect 14737 6783 14795 6789
rect 14737 6780 14749 6783
rect 14608 6752 14749 6780
rect 14608 6740 14614 6752
rect 14737 6749 14749 6752
rect 14783 6749 14795 6783
rect 15838 6780 15844 6792
rect 15799 6752 15844 6780
rect 14737 6743 14795 6749
rect 15838 6740 15844 6752
rect 15896 6740 15902 6792
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 15102 6712 15108 6724
rect 14332 6684 15108 6712
rect 14332 6672 14338 6684
rect 15102 6672 15108 6684
rect 15160 6712 15166 6724
rect 17126 6712 17132 6724
rect 15160 6684 17132 6712
rect 15160 6672 15166 6684
rect 17126 6672 17132 6684
rect 17184 6672 17190 6724
rect 13320 6616 13952 6644
rect 15289 6647 15347 6653
rect 13320 6604 13326 6616
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 17310 6644 17316 6656
rect 15335 6616 17316 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2280 6412 2973 6440
rect 2280 6400 2286 6412
rect 2961 6409 2973 6412
rect 3007 6409 3019 6443
rect 2961 6403 3019 6409
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 3418 6440 3424 6452
rect 3283 6412 3424 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 2976 6372 3004 6403
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 7282 6440 7288 6452
rect 5767 6412 7288 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 12802 6440 12808 6452
rect 8628 6412 12808 6440
rect 8628 6400 8634 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 15746 6440 15752 6452
rect 13872 6412 15752 6440
rect 13872 6400 13878 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 2976 6344 3832 6372
rect 3804 6313 3832 6344
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 7742 6372 7748 6384
rect 4120 6344 7748 6372
rect 4120 6332 4126 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 9306 6372 9312 6384
rect 9219 6344 9312 6372
rect 9306 6332 9312 6344
rect 9364 6372 9370 6384
rect 9364 6344 10916 6372
rect 9364 6332 9370 6344
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4028 6276 4905 6304
rect 4028 6264 4034 6276
rect 4893 6273 4905 6276
rect 4939 6304 4951 6307
rect 6270 6304 6276 6316
rect 4939 6276 5580 6304
rect 6231 6276 6276 6304
rect 4939 6273 4951 6276
rect 4893 6267 4951 6273
rect 1581 6239 1639 6245
rect 1581 6205 1593 6239
rect 1627 6205 1639 6239
rect 1581 6199 1639 6205
rect 1848 6239 1906 6245
rect 1848 6205 1860 6239
rect 1894 6236 1906 6239
rect 3988 6236 4016 6264
rect 1894 6208 4016 6236
rect 4617 6239 4675 6245
rect 1894 6205 1906 6208
rect 1848 6199 1906 6205
rect 1596 6100 1624 6199
rect 2516 6180 2544 6208
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 4982 6236 4988 6248
rect 4663 6208 4988 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5445 6239 5503 6245
rect 5445 6236 5457 6239
rect 5316 6208 5457 6236
rect 5316 6196 5322 6208
rect 5445 6205 5457 6208
rect 5491 6205 5503 6239
rect 5552 6236 5580 6276
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 6972 6276 7297 6304
rect 6972 6264 6978 6276
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7285 6267 7343 6273
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7374 6236 7380 6248
rect 5552 6208 7380 6236
rect 5445 6199 5503 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8018 6236 8024 6248
rect 7975 6208 8024 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8196 6239 8254 6245
rect 8196 6205 8208 6239
rect 8242 6236 8254 6239
rect 10502 6236 10508 6248
rect 8242 6208 10508 6236
rect 8242 6205 8254 6208
rect 8196 6199 8254 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 10888 6236 10916 6344
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6304 11023 6307
rect 11146 6304 11152 6316
rect 11011 6276 11152 6304
rect 11011 6273 11023 6276
rect 10965 6267 11023 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12066 6304 12072 6316
rect 12023 6276 12072 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12066 6264 12072 6276
rect 12124 6304 12130 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12124 6276 13001 6304
rect 12124 6264 12130 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 16393 6307 16451 6313
rect 12989 6267 13047 6273
rect 13556 6276 14320 6304
rect 13556 6236 13584 6276
rect 10888 6208 13584 6236
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14185 6239 14243 6245
rect 14185 6236 14197 6239
rect 13688 6208 14197 6236
rect 13688 6196 13694 6208
rect 14185 6205 14197 6208
rect 14231 6205 14243 6239
rect 14292 6236 14320 6276
rect 16393 6273 16405 6307
rect 16439 6273 16451 6307
rect 16393 6267 16451 6273
rect 15838 6236 15844 6248
rect 14292 6208 15844 6236
rect 14185 6199 14243 6205
rect 2498 6128 2504 6180
rect 2556 6128 2562 6180
rect 4522 6128 4528 6180
rect 4580 6168 4586 6180
rect 10594 6168 10600 6180
rect 4580 6140 10600 6168
rect 4580 6128 4586 6140
rect 10594 6128 10600 6140
rect 10652 6128 10658 6180
rect 10781 6171 10839 6177
rect 10781 6137 10793 6171
rect 10827 6168 10839 6171
rect 11054 6168 11060 6180
rect 10827 6140 11060 6168
rect 10827 6137 10839 6140
rect 10781 6131 10839 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 11701 6171 11759 6177
rect 11701 6137 11713 6171
rect 11747 6168 11759 6171
rect 13449 6171 13507 6177
rect 13449 6168 13461 6171
rect 11747 6140 13461 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 13449 6137 13461 6140
rect 13495 6137 13507 6171
rect 14200 6168 14228 6199
rect 15838 6196 15844 6208
rect 15896 6236 15902 6248
rect 16408 6236 16436 6267
rect 15896 6208 16436 6236
rect 15896 6196 15902 6208
rect 14458 6177 14464 6180
rect 14452 6168 14464 6177
rect 14200 6140 14320 6168
rect 14419 6140 14464 6168
rect 13449 6131 13507 6137
rect 1762 6100 1768 6112
rect 1596 6072 1768 6100
rect 1762 6060 1768 6072
rect 1820 6060 1826 6112
rect 3602 6100 3608 6112
rect 3563 6072 3608 6100
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3697 6103 3755 6109
rect 3697 6069 3709 6103
rect 3743 6100 3755 6103
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 3743 6072 4261 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 4249 6063 4307 6069
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 5074 6100 5080 6112
rect 4755 6072 5080 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6100 5319 6103
rect 5350 6100 5356 6112
rect 5307 6072 5356 6100
rect 5307 6069 5319 6072
rect 5261 6063 5319 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6181 6103 6239 6109
rect 6181 6069 6193 6103
rect 6227 6100 6239 6103
rect 6825 6103 6883 6109
rect 6825 6100 6837 6103
rect 6227 6072 6837 6100
rect 6227 6069 6239 6072
rect 6181 6063 6239 6069
rect 6825 6069 6837 6072
rect 6871 6069 6883 6103
rect 6825 6063 6883 6069
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 6972 6072 7205 6100
rect 6972 6060 6978 6072
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 7193 6063 7251 6069
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 10042 6100 10048 6112
rect 7432 6072 10048 6100
rect 7432 6060 7438 6072
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10318 6100 10324 6112
rect 10279 6072 10324 6100
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 10560 6072 10701 6100
rect 10560 6060 10566 6072
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 10928 6072 11345 6100
rect 10928 6060 10934 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11793 6103 11851 6109
rect 11793 6100 11805 6103
rect 11572 6072 11805 6100
rect 11572 6060 11578 6072
rect 11793 6069 11805 6072
rect 11839 6069 11851 6103
rect 11793 6063 11851 6069
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 11940 6072 12449 6100
rect 11940 6060 11946 6072
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12676 6072 12817 6100
rect 12676 6060 12682 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 12897 6103 12955 6109
rect 12897 6069 12909 6103
rect 12943 6100 12955 6103
rect 13170 6100 13176 6112
rect 12943 6072 13176 6100
rect 12943 6069 12955 6072
rect 12897 6063 12955 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14182 6100 14188 6112
rect 13872 6072 14188 6100
rect 13872 6060 13878 6072
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14292 6100 14320 6140
rect 14452 6131 14464 6140
rect 14458 6128 14464 6131
rect 14516 6128 14522 6180
rect 15286 6100 15292 6112
rect 14292 6072 15292 6100
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 15838 6100 15844 6112
rect 15799 6072 15844 6100
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 16206 6100 16212 6112
rect 16167 6072 16212 6100
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16298 6060 16304 6112
rect 16356 6100 16362 6112
rect 16356 6072 16401 6100
rect 16356 6060 16362 6072
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2041 5899 2099 5905
rect 2041 5896 2053 5899
rect 2004 5868 2053 5896
rect 2004 5856 2010 5868
rect 2041 5865 2053 5868
rect 2087 5865 2099 5899
rect 2041 5859 2099 5865
rect 2593 5899 2651 5905
rect 2593 5865 2605 5899
rect 2639 5896 2651 5899
rect 3602 5896 3608 5908
rect 2639 5868 3608 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 6181 5899 6239 5905
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 6270 5896 6276 5908
rect 6227 5868 6276 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 9858 5896 9864 5908
rect 6880 5868 9864 5896
rect 6880 5856 6886 5868
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10502 5896 10508 5908
rect 10463 5868 10508 5896
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 10870 5896 10876 5908
rect 10831 5868 10876 5896
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 10965 5899 11023 5905
rect 10965 5865 10977 5899
rect 11011 5896 11023 5899
rect 11882 5896 11888 5908
rect 11011 5868 11888 5896
rect 11011 5865 11023 5868
rect 10965 5859 11023 5865
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12032 5868 15700 5896
rect 12032 5856 12038 5868
rect 5068 5831 5126 5837
rect 5068 5797 5080 5831
rect 5114 5828 5126 5831
rect 7466 5828 7472 5840
rect 5114 5800 7472 5828
rect 5114 5797 5126 5800
rect 5068 5791 5126 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 7644 5831 7702 5837
rect 7644 5797 7656 5831
rect 7690 5828 7702 5831
rect 9306 5828 9312 5840
rect 7690 5800 9312 5828
rect 7690 5797 7702 5800
rect 7644 5791 7702 5797
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 10318 5788 10324 5840
rect 10376 5828 10382 5840
rect 10376 5800 11928 5828
rect 10376 5788 10382 5800
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2682 5760 2688 5772
rect 1995 5732 2688 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 2961 5763 3019 5769
rect 2961 5760 2973 5763
rect 2832 5732 2973 5760
rect 2832 5720 2838 5732
rect 2961 5729 2973 5732
rect 3007 5729 3019 5763
rect 2961 5723 3019 5729
rect 4706 5720 4712 5772
rect 4764 5760 4770 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4764 5732 4813 5760
rect 4764 5720 4770 5732
rect 4801 5729 4813 5732
rect 4847 5760 4859 5763
rect 5350 5760 5356 5772
rect 4847 5732 5356 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 5350 5720 5356 5732
rect 5408 5760 5414 5772
rect 6822 5760 6828 5772
rect 5408 5732 6828 5760
rect 5408 5720 5414 5732
rect 6822 5720 6828 5732
rect 6880 5760 6886 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 6880 5732 7389 5760
rect 6880 5720 6886 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 9214 5760 9220 5772
rect 7377 5723 7435 5729
rect 7484 5732 9220 5760
rect 2130 5692 2136 5704
rect 2091 5664 2136 5692
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3142 5692 3148 5704
rect 3099 5664 3148 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3142 5652 3148 5664
rect 3200 5652 3206 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3970 5692 3976 5704
rect 3283 5664 3976 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 7484 5692 7512 5732
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 11790 5769 11796 5772
rect 11784 5760 11796 5769
rect 11164 5732 11796 5760
rect 11164 5701 11192 5732
rect 11784 5723 11796 5732
rect 11790 5720 11796 5723
rect 11848 5720 11854 5772
rect 11900 5760 11928 5800
rect 13262 5788 13268 5840
rect 13320 5828 13326 5840
rect 15562 5837 15568 5840
rect 15556 5828 15568 5837
rect 13320 5800 13952 5828
rect 15523 5800 15568 5828
rect 13320 5788 13326 5800
rect 13538 5760 13544 5772
rect 11900 5732 12664 5760
rect 13499 5732 13544 5760
rect 6472 5664 7512 5692
rect 11149 5695 11207 5701
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 3326 5624 3332 5636
rect 1627 5596 3332 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 5074 5516 5080 5568
rect 5132 5556 5138 5568
rect 6472 5556 6500 5664
rect 11149 5661 11161 5695
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5661 11575 5695
rect 12636 5692 12664 5732
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 13814 5769 13820 5772
rect 13808 5760 13820 5769
rect 13775 5732 13820 5760
rect 13808 5723 13820 5732
rect 13814 5720 13820 5723
rect 13872 5720 13878 5772
rect 13924 5760 13952 5800
rect 15556 5791 15568 5800
rect 15562 5788 15568 5791
rect 15620 5788 15626 5840
rect 15672 5828 15700 5868
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 17405 5899 17463 5905
rect 17405 5896 17417 5899
rect 15896 5868 17417 5896
rect 15896 5856 15902 5868
rect 17405 5865 17417 5868
rect 17451 5865 17463 5899
rect 17405 5859 17463 5865
rect 16761 5831 16819 5837
rect 16761 5828 16773 5831
rect 15672 5800 16773 5828
rect 16761 5797 16773 5800
rect 16807 5797 16819 5831
rect 17310 5828 17316 5840
rect 17271 5800 17316 5828
rect 16761 5791 16819 5797
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 13924 5732 17540 5760
rect 13446 5692 13452 5704
rect 12636 5664 13452 5692
rect 11517 5655 11575 5661
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 11422 5624 11428 5636
rect 10928 5596 11428 5624
rect 10928 5584 10934 5596
rect 11422 5584 11428 5596
rect 11480 5624 11486 5636
rect 11532 5624 11560 5655
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 17512 5701 17540 5732
rect 17954 5720 17960 5772
rect 18012 5760 18018 5772
rect 18877 5763 18935 5769
rect 18877 5760 18889 5763
rect 18012 5732 18889 5760
rect 18012 5720 18018 5732
rect 18877 5729 18889 5732
rect 18923 5729 18935 5763
rect 18877 5723 18935 5729
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 19153 5695 19211 5701
rect 19153 5661 19165 5695
rect 19199 5692 19211 5695
rect 19794 5692 19800 5704
rect 19199 5664 19800 5692
rect 19199 5661 19211 5664
rect 19153 5655 19211 5661
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 12894 5624 12900 5636
rect 11480 5596 11560 5624
rect 12855 5596 12900 5624
rect 11480 5584 11486 5596
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 16669 5627 16727 5633
rect 16669 5593 16681 5627
rect 16715 5624 16727 5627
rect 16761 5627 16819 5633
rect 16761 5624 16773 5627
rect 16715 5596 16773 5624
rect 16715 5593 16727 5596
rect 16669 5587 16727 5593
rect 16761 5593 16773 5596
rect 16807 5593 16819 5627
rect 16761 5587 16819 5593
rect 5132 5528 6500 5556
rect 5132 5516 5138 5528
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6730 5556 6736 5568
rect 6604 5528 6736 5556
rect 6604 5516 6610 5528
rect 6730 5516 6736 5528
rect 6788 5556 6794 5568
rect 8018 5556 8024 5568
rect 6788 5528 8024 5556
rect 6788 5516 6794 5528
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8754 5556 8760 5568
rect 8667 5528 8760 5556
rect 8754 5516 8760 5528
rect 8812 5556 8818 5568
rect 13262 5556 13268 5568
rect 8812 5528 13268 5556
rect 8812 5516 8818 5528
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 14918 5556 14924 5568
rect 14879 5528 14924 5556
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 16945 5559 17003 5565
rect 16945 5556 16957 5559
rect 15344 5528 16957 5556
rect 15344 5516 15350 5528
rect 16945 5525 16957 5528
rect 16991 5525 17003 5559
rect 16945 5519 17003 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4798 5352 4804 5364
rect 4120 5324 4804 5352
rect 4120 5312 4126 5324
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5592 5324 6009 5352
rect 5592 5312 5598 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 5997 5315 6055 5321
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 7524 5324 7788 5352
rect 7524 5312 7530 5324
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 6178 5284 6184 5296
rect 5776 5256 6184 5284
rect 5776 5244 5782 5256
rect 6178 5244 6184 5256
rect 6236 5244 6242 5296
rect 7760 5284 7788 5324
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8481 5355 8539 5361
rect 8481 5352 8493 5355
rect 8352 5324 8493 5352
rect 8352 5312 8358 5324
rect 8481 5321 8493 5324
rect 8527 5321 8539 5355
rect 8481 5315 8539 5321
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 11112 5324 11345 5352
rect 11112 5312 11118 5324
rect 11333 5321 11345 5324
rect 11379 5321 11391 5355
rect 14182 5352 14188 5364
rect 11333 5315 11391 5321
rect 11808 5324 14188 5352
rect 7760 5256 8984 5284
rect 3878 5216 3884 5228
rect 3839 5188 3884 5216
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8956 5225 8984 5256
rect 8941 5219 8999 5225
rect 8076 5188 8892 5216
rect 8076 5176 8082 5188
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 2041 5151 2099 5157
rect 2041 5148 2053 5151
rect 1820 5120 2053 5148
rect 1820 5108 1826 5120
rect 2041 5117 2053 5120
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 2308 5151 2366 5157
rect 2308 5117 2320 5151
rect 2354 5148 2366 5151
rect 2590 5148 2596 5160
rect 2354 5120 2596 5148
rect 2354 5117 2366 5120
rect 2308 5111 2366 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 4154 5148 4160 5160
rect 3743 5120 4160 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4706 5148 4712 5160
rect 4663 5120 4712 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 6454 5148 6460 5160
rect 4816 5120 6460 5148
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 4816 5080 4844 5120
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6822 5148 6828 5160
rect 6783 5120 6828 5148
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7092 5151 7150 5157
rect 7092 5117 7104 5151
rect 7138 5148 7150 5151
rect 8754 5148 8760 5160
rect 7138 5120 8760 5148
rect 7138 5117 7150 5120
rect 7092 5111 7150 5117
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8864 5148 8892 5188
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 9048 5148 9076 5179
rect 10226 5176 10232 5228
rect 10284 5216 10290 5228
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10284 5188 10517 5216
rect 10284 5176 10290 5188
rect 10505 5185 10517 5188
rect 10551 5216 10563 5219
rect 11808 5216 11836 5324
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14277 5355 14335 5361
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 14323 5324 14381 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 14369 5321 14381 5324
rect 14415 5321 14427 5355
rect 14369 5315 14427 5321
rect 16206 5312 16212 5364
rect 16264 5352 16270 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 16264 5324 16405 5352
rect 16264 5312 16270 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 13357 5287 13415 5293
rect 13357 5253 13369 5287
rect 13403 5284 13415 5287
rect 13403 5256 15056 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 11974 5216 11980 5228
rect 10551 5188 11836 5216
rect 11935 5188 11980 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 14001 5219 14059 5225
rect 14001 5185 14013 5219
rect 14047 5216 14059 5219
rect 14458 5216 14464 5228
rect 14047 5188 14464 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14458 5176 14464 5188
rect 14516 5216 14522 5228
rect 14918 5216 14924 5228
rect 14516 5188 14924 5216
rect 14516 5176 14522 5188
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 8864 5120 9076 5148
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 12805 5151 12863 5157
rect 12805 5148 12817 5151
rect 9732 5120 12817 5148
rect 9732 5108 9738 5120
rect 12805 5117 12817 5120
rect 12851 5117 12863 5151
rect 12805 5111 12863 5117
rect 14277 5151 14335 5157
rect 14277 5117 14289 5151
rect 14323 5148 14335 5151
rect 14323 5120 14504 5148
rect 14323 5117 14335 5120
rect 14277 5111 14335 5117
rect 4028 5052 4844 5080
rect 4884 5083 4942 5089
rect 4028 5040 4034 5052
rect 4884 5049 4896 5083
rect 4930 5080 4942 5083
rect 5534 5080 5540 5092
rect 4930 5052 5540 5080
rect 4930 5049 4942 5052
rect 4884 5043 4942 5049
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 6362 5040 6368 5092
rect 6420 5080 6426 5092
rect 8849 5083 8907 5089
rect 8849 5080 8861 5083
rect 6420 5052 8861 5080
rect 6420 5040 6426 5052
rect 8849 5049 8861 5052
rect 8895 5049 8907 5083
rect 13725 5083 13783 5089
rect 13725 5080 13737 5083
rect 8849 5043 8907 5049
rect 9876 5052 13737 5080
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 3292 4984 3433 5012
rect 3292 4972 3298 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3421 4975 3479 4981
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 9876 5021 9904 5052
rect 13725 5049 13737 5052
rect 13771 5049 13783 5083
rect 14476 5080 14504 5120
rect 14550 5108 14556 5160
rect 14608 5148 14614 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 14608 5120 14749 5148
rect 14608 5108 14614 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15028 5148 15056 5256
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15620 5188 15945 5216
rect 15620 5176 15626 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 16942 5216 16948 5228
rect 16903 5188 16948 5216
rect 15933 5179 15991 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 15841 5151 15899 5157
rect 15841 5148 15853 5151
rect 14884 5120 14929 5148
rect 15028 5120 15853 5148
rect 14884 5108 14890 5120
rect 15841 5117 15853 5120
rect 15887 5117 15899 5151
rect 19794 5148 19800 5160
rect 19755 5120 19800 5148
rect 15841 5111 15899 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 14476 5052 15761 5080
rect 13725 5043 13783 5049
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 15749 5043 15807 5049
rect 15930 5040 15936 5092
rect 15988 5080 15994 5092
rect 16853 5083 16911 5089
rect 16853 5080 16865 5083
rect 15988 5052 16865 5080
rect 15988 5040 15994 5052
rect 16853 5049 16865 5052
rect 16899 5049 16911 5083
rect 16853 5043 16911 5049
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 7432 4984 8217 5012
rect 7432 4972 7438 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 4981 9919 5015
rect 9861 4975 9919 4981
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10229 5015 10287 5021
rect 10229 5012 10241 5015
rect 10192 4984 10241 5012
rect 10192 4972 10198 4984
rect 10229 4981 10241 4984
rect 10275 4981 10287 5015
rect 10229 4975 10287 4981
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10410 5012 10416 5024
rect 10367 4984 10416 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 11054 4972 11060 5024
rect 11112 5012 11118 5024
rect 11701 5015 11759 5021
rect 11701 5012 11713 5015
rect 11112 4984 11713 5012
rect 11112 4972 11118 4984
rect 11701 4981 11713 4984
rect 11747 4981 11759 5015
rect 11701 4975 11759 4981
rect 11793 5015 11851 5021
rect 11793 4981 11805 5015
rect 11839 5012 11851 5015
rect 12894 5012 12900 5024
rect 11839 4984 12900 5012
rect 11839 4981 11851 4984
rect 11793 4975 11851 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13630 5012 13636 5024
rect 13035 4984 13636 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 14182 5012 14188 5024
rect 13863 4984 14188 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16758 5012 16764 5024
rect 16719 4984 16764 5012
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 19981 5015 20039 5021
rect 19981 4981 19993 5015
rect 20027 5012 20039 5015
rect 20622 5012 20628 5024
rect 20027 4984 20628 5012
rect 20027 4981 20039 4984
rect 19981 4975 20039 4981
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 4706 4808 4712 4820
rect 1903 4780 4712 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5626 4808 5632 4820
rect 5000 4780 5632 4808
rect 4424 4743 4482 4749
rect 4424 4709 4436 4743
rect 4470 4740 4482 4743
rect 5000 4740 5028 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 6144 4780 6285 4808
rect 6144 4768 6150 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 6273 4771 6331 4777
rect 7377 4811 7435 4817
rect 7377 4777 7389 4811
rect 7423 4808 7435 4811
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 7423 4780 10149 4808
rect 7423 4777 7435 4780
rect 7377 4771 7435 4777
rect 10137 4777 10149 4780
rect 10183 4777 10195 4811
rect 10137 4771 10195 4777
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 11698 4808 11704 4820
rect 10744 4780 11704 4808
rect 10744 4768 10750 4780
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 12032 4780 12633 4808
rect 12032 4768 12038 4780
rect 12621 4777 12633 4780
rect 12667 4777 12679 4811
rect 12894 4808 12900 4820
rect 12855 4780 12900 4808
rect 12621 4771 12679 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 14182 4808 14188 4820
rect 14143 4780 14188 4808
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15289 4811 15347 4817
rect 15289 4777 15301 4811
rect 15335 4808 15347 4811
rect 16298 4808 16304 4820
rect 15335 4780 16304 4808
rect 15335 4777 15347 4780
rect 15289 4771 15347 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 7742 4740 7748 4752
rect 4470 4712 5028 4740
rect 7703 4712 7748 4740
rect 4470 4709 4482 4712
rect 4424 4703 4482 4709
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 7926 4700 7932 4752
rect 7984 4740 7990 4752
rect 13906 4740 13912 4752
rect 7984 4712 13912 4740
rect 7984 4700 7990 4712
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 13998 4700 14004 4752
rect 14056 4740 14062 4752
rect 14553 4743 14611 4749
rect 14553 4740 14565 4743
rect 14056 4712 14565 4740
rect 14056 4700 14062 4712
rect 14553 4709 14565 4712
rect 14599 4740 14611 4743
rect 15102 4740 15108 4752
rect 14599 4712 15108 4740
rect 14599 4709 14611 4712
rect 14553 4703 14611 4709
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 15378 4700 15384 4752
rect 15436 4740 15442 4752
rect 15436 4712 17080 4740
rect 15436 4700 15442 4712
rect 2222 4672 2228 4684
rect 2183 4644 2228 4672
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 3237 4675 3295 4681
rect 2372 4644 2417 4672
rect 2372 4632 2378 4644
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 4062 4672 4068 4684
rect 3283 4644 4068 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 4798 4672 4804 4684
rect 4203 4644 4804 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4982 4632 4988 4684
rect 5040 4672 5046 4684
rect 6270 4672 6276 4684
rect 5040 4644 6276 4672
rect 5040 4632 5046 4644
rect 6270 4632 6276 4644
rect 6328 4672 6334 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6328 4644 6653 4672
rect 6328 4632 6334 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 7374 4672 7380 4684
rect 6641 4635 6699 4641
rect 6932 4644 7380 4672
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3326 4604 3332 4616
rect 3287 4576 3332 4604
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 3421 4607 3479 4613
rect 3421 4573 3433 4607
rect 3467 4573 3479 4607
rect 3421 4567 3479 4573
rect 2424 4536 2452 4564
rect 3436 4536 3464 4567
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 6932 4613 6960 4644
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4641 8815 4675
rect 8757 4635 8815 4641
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 5500 4576 6745 4604
rect 5500 4564 5506 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7156 4576 7849 4604
rect 7156 4564 7162 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8202 4604 8208 4616
rect 8067 4576 8208 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8772 4604 8800 4635
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 8904 4644 8949 4672
rect 8904 4632 8910 4644
rect 9306 4632 9312 4684
rect 9364 4672 9370 4684
rect 10045 4675 10103 4681
rect 10045 4672 10057 4675
rect 9364 4644 10057 4672
rect 9364 4632 9370 4644
rect 10045 4641 10057 4644
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 11508 4675 11566 4681
rect 11508 4641 11520 4675
rect 11554 4672 11566 4675
rect 11790 4672 11796 4684
rect 11554 4644 11796 4672
rect 11554 4641 11566 4644
rect 11508 4635 11566 4641
rect 11790 4632 11796 4644
rect 11848 4672 11854 4684
rect 12066 4672 12072 4684
rect 11848 4644 12072 4672
rect 11848 4632 11854 4644
rect 12066 4632 12072 4644
rect 12124 4672 12130 4684
rect 13262 4672 13268 4684
rect 12124 4644 12296 4672
rect 13223 4644 13268 4672
rect 12124 4632 12130 4644
rect 8312 4576 8800 4604
rect 8941 4607 8999 4613
rect 5534 4536 5540 4548
rect 2424 4508 3464 4536
rect 5447 4508 5540 4536
rect 5534 4496 5540 4508
rect 5592 4536 5598 4548
rect 7650 4536 7656 4548
rect 5592 4508 7656 4536
rect 5592 4496 5598 4508
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7926 4496 7932 4548
rect 7984 4536 7990 4548
rect 8312 4536 8340 4576
rect 8941 4573 8953 4607
rect 8987 4573 8999 4607
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 8941 4567 8999 4573
rect 7984 4508 8340 4536
rect 7984 4496 7990 4508
rect 8386 4496 8392 4548
rect 8444 4536 8450 4548
rect 8444 4508 8489 4536
rect 8444 4496 8450 4508
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 5074 4468 5080 4480
rect 2915 4440 5080 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 6178 4428 6184 4480
rect 6236 4468 6242 4480
rect 8956 4468 8984 4567
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10689 4607 10747 4613
rect 10689 4604 10701 4607
rect 10376 4576 10701 4604
rect 10376 4564 10382 4576
rect 10689 4573 10701 4576
rect 10735 4573 10747 4607
rect 10689 4567 10747 4573
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 10928 4576 11253 4604
rect 10928 4564 10934 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11241 4567 11299 4573
rect 6236 4440 8984 4468
rect 9677 4471 9735 4477
rect 6236 4428 6242 4440
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 11146 4468 11152 4480
rect 9723 4440 11152 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 12268 4468 12296 4644
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 13823 4644 14657 4672
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 13823 4536 13851 4644
rect 14645 4641 14657 4644
rect 14691 4672 14703 4675
rect 14691 4644 15148 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 14737 4607 14795 4613
rect 14737 4604 14749 4607
rect 14332 4576 14749 4604
rect 14332 4564 14338 4576
rect 14737 4573 14749 4576
rect 14783 4573 14795 4607
rect 14737 4567 14795 4573
rect 12492 4508 13851 4536
rect 15120 4536 15148 4644
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15252 4644 15669 4672
rect 15252 4632 15258 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 15746 4632 15752 4684
rect 15804 4672 15810 4684
rect 17052 4681 17080 4712
rect 17037 4675 17095 4681
rect 15804 4644 15849 4672
rect 15804 4632 15810 4644
rect 17037 4641 17049 4675
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 17313 4675 17371 4681
rect 17313 4641 17325 4675
rect 17359 4672 17371 4675
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17359 4644 17877 4672
rect 17359 4641 17371 4644
rect 17313 4635 17371 4641
rect 17865 4641 17877 4644
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 15933 4607 15991 4613
rect 15933 4573 15945 4607
rect 15979 4604 15991 4607
rect 16942 4604 16948 4616
rect 15979 4576 16948 4604
rect 15979 4573 15991 4576
rect 15933 4567 15991 4573
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17034 4536 17040 4548
rect 15120 4508 17040 4536
rect 12492 4496 12498 4508
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 13538 4468 13544 4480
rect 12268 4440 13544 4468
rect 13538 4428 13544 4440
rect 13596 4428 13602 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 18782 4468 18788 4480
rect 18095 4440 18788 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 2406 4224 2412 4276
rect 2464 4264 2470 4276
rect 3145 4267 3203 4273
rect 3145 4264 3157 4267
rect 2464 4236 3157 4264
rect 2464 4224 2470 4236
rect 3145 4233 3157 4236
rect 3191 4233 3203 4267
rect 3145 4227 3203 4233
rect 5629 4267 5687 4273
rect 5629 4233 5641 4267
rect 5675 4264 5687 4267
rect 6362 4264 6368 4276
rect 5675 4236 6368 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7098 4264 7104 4276
rect 7059 4236 7104 4264
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 8113 4267 8171 4273
rect 8113 4264 8125 4267
rect 7800 4236 8125 4264
rect 7800 4224 7806 4236
rect 8113 4233 8125 4236
rect 8159 4233 8171 4267
rect 9306 4264 9312 4276
rect 9267 4236 9312 4264
rect 8113 4227 8171 4233
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 11440 4236 11928 4264
rect 4801 4199 4859 4205
rect 4801 4165 4813 4199
rect 4847 4165 4859 4199
rect 4801 4159 4859 4165
rect 4816 4128 4844 4159
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 10597 4199 10655 4205
rect 6512 4168 8800 4196
rect 6512 4156 6518 4168
rect 6178 4128 6184 4140
rect 4816 4100 6184 4128
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7340 4100 7665 4128
rect 7340 4088 7346 4100
rect 7653 4097 7665 4100
rect 7699 4128 7711 4131
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 7699 4100 8677 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 1762 4060 1768 4072
rect 1675 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4060 1826 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 1820 4032 3433 4060
rect 1820 4020 1826 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 4798 4060 4804 4072
rect 3467 4032 4804 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6730 4060 6736 4072
rect 6135 4032 6736 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 6730 4020 6736 4032
rect 6788 4020 6794 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8772 4060 8800 4168
rect 10597 4165 10609 4199
rect 10643 4196 10655 4199
rect 10781 4199 10839 4205
rect 10781 4196 10793 4199
rect 10643 4168 10793 4196
rect 10643 4165 10655 4168
rect 10597 4159 10655 4165
rect 10781 4165 10793 4168
rect 10827 4165 10839 4199
rect 10781 4159 10839 4165
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 11054 4196 11060 4208
rect 11011 4168 11060 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 9766 4128 9772 4140
rect 9727 4100 9772 4128
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4128 10011 4131
rect 10502 4128 10508 4140
rect 9999 4100 10508 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11440 4137 11468 4236
rect 11790 4196 11796 4208
rect 11532 4168 11796 4196
rect 11532 4137 11560 4168
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 11425 4131 11483 4137
rect 11425 4128 11437 4131
rect 11296 4100 11437 4128
rect 11296 4088 11302 4100
rect 11425 4097 11437 4100
rect 11471 4097 11483 4131
rect 11425 4091 11483 4097
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4097 11575 4131
rect 11900 4128 11928 4236
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13817 4267 13875 4273
rect 13817 4264 13829 4267
rect 13596 4236 13829 4264
rect 13596 4224 13602 4236
rect 13817 4233 13829 4236
rect 13863 4233 13875 4267
rect 13817 4227 13875 4233
rect 14016 4236 14596 4264
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 14016 4196 14044 4236
rect 13504 4168 14044 4196
rect 14093 4199 14151 4205
rect 13504 4156 13510 4168
rect 14093 4165 14105 4199
rect 14139 4165 14151 4199
rect 14568 4196 14596 4236
rect 14568 4168 14688 4196
rect 14093 4159 14151 4165
rect 14108 4128 14136 4159
rect 14660 4137 14688 4168
rect 14645 4131 14703 4137
rect 11900 4100 12572 4128
rect 14108 4100 14596 4128
rect 11517 4091 11575 4097
rect 9490 4060 9496 4072
rect 8527 4032 9496 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4060 9735 4063
rect 10318 4060 10324 4072
rect 9723 4032 10324 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 10318 4020 10324 4032
rect 10376 4020 10382 4072
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4060 10471 4063
rect 11698 4060 11704 4072
rect 10459 4032 11704 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12124 4032 12449 4060
rect 12124 4020 12130 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12544 4060 12572 4100
rect 14458 4060 14464 4072
rect 12544 4032 12940 4060
rect 14419 4032 14464 4060
rect 12437 4023 12495 4029
rect 2032 3995 2090 4001
rect 2032 3961 2044 3995
rect 2078 3992 2090 3995
rect 3234 3992 3240 4004
rect 2078 3964 3240 3992
rect 2078 3961 2090 3964
rect 2032 3955 2090 3961
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 3688 3995 3746 4001
rect 3688 3961 3700 3995
rect 3734 3992 3746 3995
rect 3734 3964 3832 3992
rect 3734 3961 3746 3964
rect 3688 3955 3746 3961
rect 3804 3924 3832 3964
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 4246 3992 4252 4004
rect 3936 3964 4252 3992
rect 3936 3952 3942 3964
rect 4246 3952 4252 3964
rect 4304 3952 4310 4004
rect 10134 3992 10140 4004
rect 7760 3964 10140 3992
rect 7760 3936 7788 3964
rect 10134 3952 10140 3964
rect 10192 3992 10198 4004
rect 10594 3992 10600 4004
rect 10192 3964 10600 3992
rect 10192 3952 10198 3964
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10781 3995 10839 4001
rect 10781 3961 10793 3995
rect 10827 3992 10839 3995
rect 12704 3995 12762 4001
rect 10827 3964 12664 3992
rect 10827 3961 10839 3964
rect 10781 3955 10839 3961
rect 3970 3924 3976 3936
rect 3804 3896 3976 3924
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 5166 3924 5172 3936
rect 5127 3896 5172 3924
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5534 3924 5540 3936
rect 5316 3896 5540 3924
rect 5316 3884 5322 3896
rect 5534 3884 5540 3896
rect 5592 3924 5598 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5592 3896 6009 3924
rect 5592 3884 5598 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7469 3927 7527 3933
rect 7469 3924 7481 3927
rect 7156 3896 7481 3924
rect 7156 3884 7162 3896
rect 7469 3893 7481 3896
rect 7515 3893 7527 3927
rect 7469 3887 7527 3893
rect 7561 3927 7619 3933
rect 7561 3893 7573 3927
rect 7607 3924 7619 3927
rect 7742 3924 7748 3936
rect 7607 3896 7748 3924
rect 7607 3893 7619 3896
rect 7561 3887 7619 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8570 3924 8576 3936
rect 8531 3896 8576 3924
rect 8570 3884 8576 3896
rect 8628 3924 8634 3936
rect 11330 3924 11336 3936
rect 8628 3896 11336 3924
rect 8628 3884 8634 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 11790 3924 11796 3936
rect 11664 3896 11796 3924
rect 11664 3884 11670 3896
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12636 3924 12664 3964
rect 12704 3961 12716 3995
rect 12750 3992 12762 3995
rect 12802 3992 12808 4004
rect 12750 3964 12808 3992
rect 12750 3961 12762 3964
rect 12704 3955 12762 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 12912 3992 12940 4032
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 14568 4060 14596 4100
rect 14645 4097 14657 4131
rect 14691 4097 14703 4131
rect 15930 4128 15936 4140
rect 14645 4091 14703 4097
rect 15028 4100 15936 4128
rect 15028 4060 15056 4100
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 14568 4032 15056 4060
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 14553 3995 14611 4001
rect 14553 3992 14565 3995
rect 12912 3964 14565 3992
rect 14553 3961 14565 3964
rect 14599 3961 14611 3995
rect 14553 3955 14611 3961
rect 14642 3952 14648 4004
rect 14700 3952 14706 4004
rect 15010 3952 15016 4004
rect 15068 3992 15074 4004
rect 15120 3992 15148 4023
rect 15068 3964 15148 3992
rect 15068 3952 15074 3964
rect 13170 3924 13176 3936
rect 12636 3896 13176 3924
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 14660 3924 14688 3952
rect 15289 3927 15347 3933
rect 15289 3924 15301 3927
rect 14660 3896 15301 3924
rect 15289 3893 15301 3896
rect 15335 3893 15347 3927
rect 15289 3887 15347 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 3568 3692 5120 3720
rect 3568 3680 3574 3692
rect 2032 3655 2090 3661
rect 2032 3621 2044 3655
rect 2078 3652 2090 3655
rect 2406 3652 2412 3664
rect 2078 3624 2412 3652
rect 2078 3621 2090 3624
rect 2032 3615 2090 3621
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 4798 3652 4804 3664
rect 4172 3624 4804 3652
rect 4172 3593 4200 3624
rect 4798 3612 4804 3624
rect 4856 3612 4862 3664
rect 5092 3652 5120 3692
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5224 3692 6193 3720
rect 5224 3680 5230 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 10410 3720 10416 3732
rect 7156 3692 10416 3720
rect 7156 3680 7162 3692
rect 10410 3680 10416 3692
rect 10468 3720 10474 3732
rect 11054 3720 11060 3732
rect 10468 3692 11060 3720
rect 10468 3680 10474 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 13081 3723 13139 3729
rect 13081 3689 13093 3723
rect 13127 3720 13139 3723
rect 13354 3720 13360 3732
rect 13127 3692 13360 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 8570 3652 8576 3664
rect 5092 3624 8576 3652
rect 8570 3612 8576 3624
rect 8628 3612 8634 3664
rect 8941 3655 8999 3661
rect 8941 3621 8953 3655
rect 8987 3652 8999 3655
rect 9674 3652 9680 3664
rect 8987 3624 9680 3652
rect 8987 3621 8999 3624
rect 8941 3615 8999 3621
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 10036 3655 10094 3661
rect 10036 3621 10048 3655
rect 10082 3652 10094 3655
rect 10226 3652 10232 3664
rect 10082 3624 10232 3652
rect 10082 3621 10094 3624
rect 10036 3615 10094 3621
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 11164 3652 11192 3683
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 16758 3720 16764 3732
rect 13740 3692 16764 3720
rect 11606 3652 11612 3664
rect 11164 3624 11612 3652
rect 11606 3612 11612 3624
rect 11664 3661 11670 3664
rect 11664 3655 11728 3661
rect 11664 3621 11682 3655
rect 11716 3621 11728 3655
rect 11664 3615 11728 3621
rect 11664 3612 11670 3615
rect 11790 3612 11796 3664
rect 11848 3652 11854 3664
rect 13740 3652 13768 3692
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 11848 3624 13768 3652
rect 11848 3612 11854 3624
rect 13814 3612 13820 3664
rect 13872 3652 13878 3664
rect 13872 3624 14136 3652
rect 13872 3612 13878 3624
rect 4157 3587 4215 3593
rect 4157 3553 4169 3587
rect 4203 3553 4215 3587
rect 4157 3547 4215 3553
rect 4424 3587 4482 3593
rect 4424 3553 4436 3587
rect 4470 3584 4482 3587
rect 4470 3556 6408 3584
rect 4470 3553 4482 3556
rect 4424 3547 4482 3553
rect 6380 3528 6408 3556
rect 6822 3544 6828 3596
rect 6880 3584 6886 3596
rect 7282 3593 7288 3596
rect 7009 3587 7067 3593
rect 7009 3584 7021 3587
rect 6880 3556 7021 3584
rect 6880 3544 6886 3556
rect 7009 3553 7021 3556
rect 7055 3553 7067 3587
rect 7276 3584 7288 3593
rect 7243 3556 7288 3584
rect 7009 3547 7067 3553
rect 7276 3547 7288 3556
rect 7282 3544 7288 3547
rect 7340 3544 7346 3596
rect 7558 3544 7564 3596
rect 7616 3584 7622 3596
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 7616 3556 8677 3584
rect 7616 3544 7622 3556
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 11238 3584 11244 3596
rect 8665 3547 8723 3553
rect 9692 3556 11244 3584
rect 1762 3516 1768 3528
rect 1723 3488 1768 3516
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 3418 3516 3424 3528
rect 3379 3488 3424 3516
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 5224 3488 6285 3516
rect 5224 3476 5230 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6362 3476 6368 3528
rect 6420 3516 6426 3528
rect 6420 3488 6465 3516
rect 6420 3476 6426 3488
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9692 3516 9720 3556
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 12066 3584 12072 3596
rect 11440 3556 12072 3584
rect 11440 3528 11468 3556
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12250 3544 12256 3596
rect 12308 3584 12314 3596
rect 12308 3556 12480 3584
rect 12308 3544 12314 3556
rect 8996 3488 9720 3516
rect 8996 3476 9002 3488
rect 9766 3476 9772 3528
rect 9824 3516 9830 3528
rect 11422 3516 11428 3528
rect 9824 3488 9917 3516
rect 11383 3488 11428 3516
rect 9824 3476 9830 3488
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 12452 3516 12480 3556
rect 12526 3544 12532 3596
rect 12584 3584 12590 3596
rect 13449 3587 13507 3593
rect 13449 3584 13461 3587
rect 12584 3556 13461 3584
rect 12584 3544 12590 3556
rect 13449 3553 13461 3556
rect 13495 3584 13507 3587
rect 13906 3584 13912 3596
rect 13495 3556 13912 3584
rect 13495 3553 13507 3556
rect 13449 3547 13507 3553
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 14108 3593 14136 3624
rect 14093 3587 14151 3593
rect 14093 3553 14105 3587
rect 14139 3553 14151 3587
rect 14093 3547 14151 3553
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 12894 3516 12900 3528
rect 12452 3488 12900 3516
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 6638 3448 6644 3460
rect 5859 3420 6644 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 9784 3448 9812 3476
rect 12802 3448 12808 3460
rect 8260 3420 9812 3448
rect 12715 3420 12808 3448
rect 8260 3408 8266 3420
rect 12802 3408 12808 3420
rect 12860 3448 12866 3460
rect 13648 3448 13676 3479
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14056 3488 14289 3516
rect 14056 3476 14062 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 15304 3448 15332 3547
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15436 3556 16037 3584
rect 15436 3544 15442 3556
rect 16025 3553 16037 3556
rect 16071 3553 16083 3587
rect 16025 3547 16083 3553
rect 15565 3519 15623 3525
rect 15565 3485 15577 3519
rect 15611 3516 15623 3519
rect 16114 3516 16120 3528
rect 15611 3488 16120 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 12860 3420 13676 3448
rect 13740 3420 15332 3448
rect 12860 3408 12866 3420
rect 3145 3383 3203 3389
rect 3145 3349 3157 3383
rect 3191 3380 3203 3383
rect 3970 3380 3976 3392
rect 3191 3352 3976 3380
rect 3191 3349 3203 3352
rect 3145 3343 3203 3349
rect 3970 3340 3976 3352
rect 4028 3380 4034 3392
rect 5258 3380 5264 3392
rect 4028 3352 5264 3380
rect 4028 3340 4034 3352
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5537 3383 5595 3389
rect 5537 3349 5549 3383
rect 5583 3380 5595 3383
rect 5626 3380 5632 3392
rect 5583 3352 5632 3380
rect 5583 3349 5595 3352
rect 5537 3343 5595 3349
rect 5626 3340 5632 3352
rect 5684 3380 5690 3392
rect 6546 3380 6552 3392
rect 5684 3352 6552 3380
rect 5684 3340 5690 3352
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 8294 3340 8300 3392
rect 8352 3380 8358 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 8352 3352 8401 3380
rect 8352 3340 8358 3352
rect 8389 3349 8401 3352
rect 8435 3380 8447 3383
rect 10502 3380 10508 3392
rect 8435 3352 10508 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 11790 3340 11796 3392
rect 11848 3380 11854 3392
rect 12526 3380 12532 3392
rect 11848 3352 12532 3380
rect 11848 3340 11854 3352
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 13740 3380 13768 3420
rect 12676 3352 13768 3380
rect 12676 3340 12682 3352
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 16209 3383 16267 3389
rect 16209 3380 16221 3383
rect 14148 3352 16221 3380
rect 14148 3340 14154 3352
rect 16209 3349 16221 3352
rect 16255 3349 16267 3383
rect 16209 3343 16267 3349
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3384 3148 3709 3176
rect 3384 3136 3390 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 4212 3148 4721 3176
rect 4212 3136 4218 3148
rect 4709 3145 4721 3148
rect 4755 3145 4767 3179
rect 4709 3139 4767 3145
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5350 3176 5356 3188
rect 4856 3148 5356 3176
rect 4856 3136 4862 3148
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 8386 3176 8392 3188
rect 5767 3148 8392 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 9364 3148 9597 3176
rect 9364 3136 9370 3148
rect 9585 3145 9597 3148
rect 9631 3176 9643 3179
rect 10226 3176 10232 3188
rect 9631 3148 10232 3176
rect 9631 3145 9643 3148
rect 9585 3139 9643 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 13357 3179 13415 3185
rect 13357 3176 13369 3179
rect 12483 3148 13369 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 13357 3145 13369 3148
rect 13403 3145 13415 3179
rect 13357 3139 13415 3145
rect 14369 3179 14427 3185
rect 14369 3145 14381 3179
rect 14415 3176 14427 3179
rect 21082 3176 21088 3188
rect 14415 3148 21088 3176
rect 14415 3145 14427 3148
rect 14369 3139 14427 3145
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 7282 3068 7288 3120
rect 7340 3108 7346 3120
rect 7340 3080 7604 3108
rect 7340 3068 7346 3080
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 2961 3043 3019 3049
rect 2961 3040 2973 3043
rect 2924 3012 2973 3040
rect 2924 3000 2930 3012
rect 2961 3009 2973 3012
rect 3007 3040 3019 3043
rect 3234 3040 3240 3052
rect 3007 3012 3240 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3234 3000 3240 3012
rect 3292 3040 3298 3052
rect 3970 3040 3976 3052
rect 3292 3012 3976 3040
rect 3292 3000 3298 3012
rect 3970 3000 3976 3012
rect 4028 3040 4034 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4028 3012 4261 3040
rect 4028 3000 4034 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 5258 3040 5264 3052
rect 5219 3012 5264 3040
rect 4249 3003 4307 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 3050 2972 3056 2984
rect 2731 2944 3056 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 5166 2972 5172 2984
rect 5127 2944 5172 2972
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6380 2972 6408 3003
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7576 3049 7604 3080
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 11112 3080 11551 3108
rect 11112 3068 11118 3080
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7156 3012 7481 3040
rect 7156 3000 7162 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 9214 3000 9220 3052
rect 9272 3040 9278 3052
rect 9858 3040 9864 3052
rect 9272 3012 9864 3040
rect 9272 3000 9278 3012
rect 9858 3000 9864 3012
rect 9916 3040 9922 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 9916 3012 10425 3040
rect 9916 3000 9922 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 11425 3043 11483 3049
rect 11425 3040 11437 3043
rect 10560 3012 11437 3040
rect 10560 3000 10566 3012
rect 11425 3009 11437 3012
rect 11471 3009 11483 3043
rect 11523 3040 11551 3080
rect 12710 3068 12716 3120
rect 12768 3108 12774 3120
rect 14274 3108 14280 3120
rect 12768 3080 14280 3108
rect 12768 3068 12774 3080
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 14921 3111 14979 3117
rect 14921 3077 14933 3111
rect 14967 3108 14979 3111
rect 16022 3108 16028 3120
rect 14967 3080 16028 3108
rect 14967 3077 14979 3080
rect 14921 3071 14979 3077
rect 16022 3068 16028 3080
rect 16080 3068 16086 3120
rect 18509 3111 18567 3117
rect 18509 3077 18521 3111
rect 18555 3108 18567 3111
rect 19242 3108 19248 3120
rect 18555 3080 19248 3108
rect 18555 3077 18567 3080
rect 18509 3071 18567 3077
rect 19242 3068 19248 3080
rect 19300 3068 19306 3120
rect 13081 3043 13139 3049
rect 11523 3012 12848 3040
rect 11425 3003 11483 3009
rect 8202 2972 8208 2984
rect 6380 2944 8064 2972
rect 8163 2944 8208 2972
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 4246 2904 4252 2916
rect 4111 2876 4252 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 4706 2864 4712 2916
rect 4764 2904 4770 2916
rect 5077 2907 5135 2913
rect 5077 2904 5089 2907
rect 4764 2876 5089 2904
rect 4764 2864 4770 2876
rect 5077 2873 5089 2876
rect 5123 2873 5135 2907
rect 5810 2904 5816 2916
rect 5077 2867 5135 2873
rect 5368 2876 5816 2904
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3602 2836 3608 2848
rect 2832 2808 3608 2836
rect 2832 2796 2838 2808
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 5368 2836 5396 2876
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 6089 2907 6147 2913
rect 6089 2873 6101 2907
rect 6135 2904 6147 2907
rect 7558 2904 7564 2916
rect 6135 2876 7564 2904
rect 6135 2873 6147 2876
rect 6089 2867 6147 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8036 2904 8064 2944
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 10778 2972 10784 2984
rect 10275 2944 10784 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 10778 2932 10784 2944
rect 10836 2932 10842 2984
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 12820 2981 12848 3012
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13354 3040 13360 3052
rect 13127 3012 13360 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 15378 3040 15384 3052
rect 13771 3012 15384 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 22462 3040 22468 3052
rect 15488 3012 22468 3040
rect 12805 2975 12863 2981
rect 11112 2944 11468 2972
rect 11112 2932 11118 2944
rect 8294 2904 8300 2916
rect 8036 2876 8300 2904
rect 8294 2864 8300 2876
rect 8352 2904 8358 2916
rect 8450 2907 8508 2913
rect 8450 2904 8462 2907
rect 8352 2876 8462 2904
rect 8352 2864 8358 2876
rect 8450 2873 8462 2876
rect 8496 2873 8508 2907
rect 11333 2907 11391 2913
rect 11333 2904 11345 2907
rect 8450 2867 8508 2873
rect 9876 2876 11345 2904
rect 4203 2808 5396 2836
rect 6181 2839 6239 2845
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 7009 2839 7067 2845
rect 7009 2836 7021 2839
rect 6227 2808 7021 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 7009 2805 7021 2808
rect 7055 2805 7067 2839
rect 7009 2799 7067 2805
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 7377 2839 7435 2845
rect 7377 2836 7389 2839
rect 7340 2808 7389 2836
rect 7340 2796 7346 2808
rect 7377 2805 7389 2808
rect 7423 2805 7435 2839
rect 7377 2799 7435 2805
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 8754 2836 8760 2848
rect 8260 2808 8760 2836
rect 8260 2796 8266 2808
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 9876 2845 9904 2876
rect 11333 2873 11345 2876
rect 11379 2873 11391 2907
rect 11440 2904 11468 2944
rect 12805 2941 12817 2975
rect 12851 2941 12863 2975
rect 13449 2975 13507 2981
rect 13449 2972 13461 2975
rect 12805 2935 12863 2941
rect 12912 2944 13461 2972
rect 12912 2904 12940 2944
rect 13449 2941 13461 2944
rect 13495 2941 13507 2975
rect 13449 2935 13507 2941
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13964 2944 14197 2972
rect 13964 2932 13970 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 14185 2935 14243 2941
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 15102 2932 15108 2984
rect 15160 2972 15166 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 15160 2944 15301 2972
rect 15160 2932 15166 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15488 2972 15516 3012
rect 22462 3000 22468 3012
rect 22520 3000 22526 3052
rect 16114 2972 16120 2984
rect 15289 2935 15347 2941
rect 15396 2944 15516 2972
rect 16075 2944 16120 2972
rect 11440 2876 12940 2904
rect 13357 2907 13415 2913
rect 11333 2867 11391 2873
rect 13357 2873 13369 2907
rect 13403 2904 13415 2907
rect 15194 2904 15200 2916
rect 13403 2876 15200 2904
rect 13403 2873 13415 2876
rect 13357 2867 13415 2873
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2805 9919 2839
rect 10318 2836 10324 2848
rect 10279 2808 10324 2836
rect 9861 2799 9919 2805
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 10410 2796 10416 2848
rect 10468 2836 10474 2848
rect 10873 2839 10931 2845
rect 10873 2836 10885 2839
rect 10468 2808 10885 2836
rect 10468 2796 10474 2808
rect 10873 2805 10885 2808
rect 10919 2805 10931 2839
rect 11238 2836 11244 2848
rect 11199 2808 11244 2836
rect 10873 2799 10931 2805
rect 11238 2796 11244 2808
rect 11296 2796 11302 2848
rect 12894 2836 12900 2848
rect 12807 2808 12900 2836
rect 12894 2796 12900 2808
rect 12952 2836 12958 2848
rect 13262 2836 13268 2848
rect 12952 2808 13268 2836
rect 12952 2796 12958 2808
rect 13262 2796 13268 2808
rect 13320 2836 13326 2848
rect 15396 2836 15424 2944
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 17034 2972 17040 2984
rect 16995 2944 17040 2972
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17126 2932 17132 2984
rect 17184 2972 17190 2984
rect 18325 2975 18383 2981
rect 18325 2972 18337 2975
rect 17184 2944 18337 2972
rect 17184 2932 17190 2944
rect 18325 2941 18337 2944
rect 18371 2941 18383 2975
rect 18874 2972 18880 2984
rect 18835 2944 18880 2972
rect 18325 2935 18383 2941
rect 18874 2932 18880 2944
rect 18932 2932 18938 2984
rect 22002 2904 22008 2916
rect 15488 2876 22008 2904
rect 15488 2845 15516 2876
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 13320 2808 15424 2836
rect 15473 2839 15531 2845
rect 13320 2796 13326 2808
rect 15473 2805 15485 2839
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 16942 2836 16948 2848
rect 16347 2808 16948 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2836 17279 2839
rect 17862 2836 17868 2848
rect 17267 2808 17868 2836
rect 17267 2805 17279 2808
rect 17221 2799 17279 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 19061 2839 19119 2845
rect 19061 2805 19073 2839
rect 19107 2836 19119 2839
rect 19702 2836 19708 2848
rect 19107 2808 19708 2836
rect 19107 2805 19119 2808
rect 19061 2799 19119 2805
rect 19702 2796 19708 2808
rect 19760 2796 19766 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 21542 2836 21548 2848
rect 19852 2808 21548 2836
rect 19852 2796 19858 2808
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 2222 2632 2228 2644
rect 2183 2604 2228 2632
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2593 2635 2651 2641
rect 2593 2601 2605 2635
rect 2639 2632 2651 2635
rect 3418 2632 3424 2644
rect 2639 2604 3424 2632
rect 2639 2601 2651 2604
rect 2593 2595 2651 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 4062 2632 4068 2644
rect 4023 2604 4068 2632
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2632 5411 2635
rect 7374 2632 7380 2644
rect 5399 2604 7380 2632
rect 5399 2601 5411 2604
rect 5353 2595 5411 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 7558 2632 7564 2644
rect 7519 2604 7564 2632
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 9033 2635 9091 2641
rect 9033 2632 9045 2635
rect 8444 2604 9045 2632
rect 8444 2592 8450 2604
rect 9033 2601 9045 2604
rect 9079 2601 9091 2635
rect 9033 2595 9091 2601
rect 9125 2635 9183 2641
rect 9125 2601 9137 2635
rect 9171 2632 9183 2635
rect 10410 2632 10416 2644
rect 9171 2604 10416 2632
rect 9171 2601 9183 2604
rect 9125 2595 9183 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11977 2635 12035 2641
rect 11977 2601 11989 2635
rect 12023 2601 12035 2635
rect 11977 2595 12035 2601
rect 13541 2635 13599 2641
rect 13541 2601 13553 2635
rect 13587 2632 13599 2635
rect 19794 2632 19800 2644
rect 13587 2604 19800 2632
rect 13587 2601 13599 2604
rect 13541 2595 13599 2601
rect 2685 2567 2743 2573
rect 2685 2533 2697 2567
rect 2731 2564 2743 2567
rect 2958 2564 2964 2576
rect 2731 2536 2964 2564
rect 2731 2533 2743 2536
rect 2685 2527 2743 2533
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 3970 2524 3976 2576
rect 4028 2564 4034 2576
rect 5994 2564 6000 2576
rect 4028 2536 4660 2564
rect 4028 2524 4034 2536
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 4154 2496 4160 2508
rect 3844 2468 4160 2496
rect 3844 2456 3850 2468
rect 4154 2456 4160 2468
rect 4212 2496 4218 2508
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 4212 2468 4445 2496
rect 4212 2456 4218 2468
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 2866 2428 2872 2440
rect 2827 2400 2872 2428
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 4632 2437 4660 2536
rect 5828 2536 6000 2564
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 5721 2499 5779 2505
rect 5721 2496 5733 2499
rect 5316 2468 5733 2496
rect 5316 2456 5322 2468
rect 5721 2465 5733 2468
rect 5767 2465 5779 2499
rect 5721 2459 5779 2465
rect 5828 2440 5856 2536
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 8110 2524 8116 2576
rect 8168 2564 8174 2576
rect 9582 2564 9588 2576
rect 8168 2536 9588 2564
rect 8168 2524 8174 2536
rect 9582 2524 9588 2536
rect 9640 2564 9646 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9640 2536 10149 2564
rect 9640 2524 9646 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 10778 2524 10784 2576
rect 10836 2564 10842 2576
rect 11992 2564 12020 2595
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 20162 2564 20168 2576
rect 10836 2536 11836 2564
rect 11992 2536 20168 2564
rect 10836 2524 10842 2536
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 11808 2505 11836 2536
rect 20162 2524 20168 2536
rect 20220 2524 20226 2576
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 5960 2468 7941 2496
rect 5960 2456 5966 2468
rect 7929 2465 7941 2468
rect 7975 2465 7987 2499
rect 10229 2499 10287 2505
rect 7929 2459 7987 2465
rect 8220 2468 9720 2496
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 4617 2391 4675 2397
rect 4540 2360 4568 2391
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6362 2428 6368 2440
rect 6043 2400 6368 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7558 2428 7564 2440
rect 7064 2400 7564 2428
rect 7064 2388 7070 2400
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 8018 2428 8024 2440
rect 7979 2400 8024 2428
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8220 2437 8248 2468
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8938 2428 8944 2440
rect 8205 2391 8263 2397
rect 8588 2400 8944 2428
rect 6178 2360 6184 2372
rect 4540 2332 6184 2360
rect 6178 2320 6184 2332
rect 6236 2320 6242 2372
rect 8036 2360 8064 2388
rect 8588 2360 8616 2400
rect 8938 2388 8944 2400
rect 8996 2388 9002 2440
rect 9306 2428 9312 2440
rect 9267 2400 9312 2428
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9692 2428 9720 2468
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 11793 2499 11851 2505
rect 10275 2468 11376 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 9858 2428 9864 2440
rect 9692 2400 9864 2428
rect 9858 2388 9864 2400
rect 9916 2428 9922 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9916 2400 10333 2428
rect 9916 2388 9922 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 10321 2391 10379 2397
rect 10428 2400 11253 2428
rect 8036 2332 8616 2360
rect 8665 2363 8723 2369
rect 8665 2329 8677 2363
rect 8711 2360 8723 2363
rect 10428 2360 10456 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 8711 2332 10456 2360
rect 10781 2363 10839 2369
rect 8711 2329 8723 2332
rect 8665 2323 8723 2329
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11054 2360 11060 2372
rect 10827 2332 11060 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 11348 2360 11376 2468
rect 11793 2465 11805 2499
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12667 2468 13032 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2428 11483 2431
rect 11606 2428 11612 2440
rect 11471 2400 11612 2428
rect 11471 2397 11483 2400
rect 11425 2391 11483 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 11756 2400 12817 2428
rect 11756 2388 11762 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 12894 2360 12900 2372
rect 11348 2332 12900 2360
rect 12894 2320 12900 2332
rect 12952 2320 12958 2372
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 6086 2292 6092 2304
rect 4120 2264 6092 2292
rect 4120 2252 4126 2264
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 11146 2292 11152 2304
rect 9815 2264 11152 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 13004 2292 13032 2468
rect 13078 2456 13084 2508
rect 13136 2496 13142 2508
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 13136 2468 13369 2496
rect 13136 2456 13142 2468
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 13998 2496 14004 2508
rect 13959 2468 14004 2496
rect 13357 2459 13415 2465
rect 13998 2456 14004 2468
rect 14056 2456 14062 2508
rect 14182 2456 14188 2508
rect 14240 2496 14246 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14240 2468 14749 2496
rect 14240 2456 14246 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 14826 2456 14832 2508
rect 14884 2496 14890 2508
rect 15286 2496 15292 2508
rect 14884 2468 15292 2496
rect 14884 2456 14890 2468
rect 15286 2456 15292 2468
rect 15344 2456 15350 2508
rect 15657 2499 15715 2505
rect 15657 2465 15669 2499
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 15672 2428 15700 2459
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 17494 2496 17500 2508
rect 16632 2468 16677 2496
rect 17455 2468 17500 2496
rect 16632 2456 16638 2468
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 13596 2400 15700 2428
rect 13596 2388 13602 2400
rect 14185 2363 14243 2369
rect 14185 2329 14197 2363
rect 14231 2360 14243 2363
rect 15010 2360 15016 2372
rect 14231 2332 15016 2360
rect 14231 2329 14243 2332
rect 14185 2323 14243 2329
rect 15010 2320 15016 2332
rect 15068 2320 15074 2372
rect 14826 2292 14832 2304
rect 13004 2264 14832 2292
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 15562 2292 15568 2304
rect 14967 2264 15568 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 15841 2295 15899 2301
rect 15841 2261 15853 2295
rect 15887 2292 15899 2295
rect 16482 2292 16488 2304
rect 15887 2264 16488 2292
rect 15887 2261 15899 2264
rect 15841 2255 15899 2261
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 17402 2292 17408 2304
rect 16807 2264 17408 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 17402 2252 17408 2264
rect 17460 2252 17466 2304
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17954 2292 17960 2304
rect 17727 2264 17960 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 1118 2048 1124 2100
rect 1176 2088 1182 2100
rect 6454 2088 6460 2100
rect 1176 2060 6460 2088
rect 1176 2048 1182 2060
rect 6454 2048 6460 2060
rect 6512 2088 6518 2100
rect 7282 2088 7288 2100
rect 6512 2060 7288 2088
rect 6512 2048 6518 2060
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 13538 2088 13544 2100
rect 7852 2060 13544 2088
rect 198 1980 204 2032
rect 256 2020 262 2032
rect 5442 2020 5448 2032
rect 256 1992 5448 2020
rect 256 1980 262 1992
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
rect 5810 1980 5816 2032
rect 5868 2020 5874 2032
rect 7852 2020 7880 2060
rect 13538 2048 13544 2060
rect 13596 2048 13602 2100
rect 5868 1992 7880 2020
rect 5868 1980 5874 1992
rect 11330 1980 11336 2032
rect 11388 2020 11394 2032
rect 12158 2020 12164 2032
rect 11388 1992 12164 2020
rect 11388 1980 11394 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 658 1912 664 1964
rect 716 1952 722 1964
rect 7098 1952 7104 1964
rect 716 1924 7104 1952
rect 716 1912 722 1924
rect 7098 1912 7104 1924
rect 7156 1912 7162 1964
rect 2038 1844 2044 1896
rect 2096 1884 2102 1896
rect 5902 1884 5908 1896
rect 2096 1856 5908 1884
rect 2096 1844 2102 1856
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 3326 1776 3332 1828
rect 3384 1816 3390 1828
rect 8846 1816 8852 1828
rect 3384 1788 8852 1816
rect 3384 1776 3390 1788
rect 8846 1776 8852 1788
rect 8904 1776 8910 1828
rect 2498 1708 2504 1760
rect 2556 1748 2562 1760
rect 7742 1748 7748 1760
rect 2556 1720 7748 1748
rect 2556 1708 2562 1720
rect 7742 1708 7748 1720
rect 7800 1708 7806 1760
rect 1578 1640 1584 1692
rect 1636 1680 1642 1692
rect 8018 1680 8024 1692
rect 1636 1652 8024 1680
rect 1636 1640 1642 1652
rect 8018 1640 8024 1652
rect 8076 1640 8082 1692
<< via1 >>
rect 3884 20544 3936 20596
rect 6368 20544 6420 20596
rect 4436 20204 4488 20256
rect 8944 20204 8996 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 4160 20000 4212 20052
rect 4436 20043 4488 20052
rect 4436 20009 4445 20043
rect 4445 20009 4479 20043
rect 4479 20009 4488 20043
rect 4436 20000 4488 20009
rect 5172 20000 5224 20052
rect 12440 20000 12492 20052
rect 12900 20000 12952 20052
rect 13360 20043 13412 20052
rect 13360 20009 13369 20043
rect 13369 20009 13403 20043
rect 13403 20009 13412 20043
rect 13360 20000 13412 20009
rect 14556 20000 14608 20052
rect 15200 20000 15252 20052
rect 15660 20043 15712 20052
rect 15660 20009 15669 20043
rect 15669 20009 15703 20043
rect 15703 20009 15712 20043
rect 15660 20000 15712 20009
rect 16580 20000 16632 20052
rect 17960 20000 18012 20052
rect 2872 19864 2924 19916
rect 3056 19907 3108 19916
rect 3056 19873 3065 19907
rect 3065 19873 3099 19907
rect 3099 19873 3108 19907
rect 3056 19864 3108 19873
rect 5816 19932 5868 19984
rect 6920 19932 6972 19984
rect 5264 19864 5316 19916
rect 6460 19864 6512 19916
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 4988 19796 5040 19848
rect 8760 19864 8812 19916
rect 10600 19907 10652 19916
rect 7196 19796 7248 19848
rect 8300 19839 8352 19848
rect 8300 19805 8309 19839
rect 8309 19805 8343 19839
rect 8343 19805 8352 19839
rect 8300 19796 8352 19805
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 8208 19728 8260 19780
rect 8484 19796 8536 19848
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 11060 19864 11112 19916
rect 12256 19864 12308 19916
rect 13820 19864 13872 19916
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 14464 19864 14516 19916
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 15568 19864 15620 19916
rect 17132 19907 17184 19916
rect 17132 19873 17141 19907
rect 17141 19873 17175 19907
rect 17175 19873 17184 19907
rect 17132 19864 17184 19873
rect 9680 19796 9732 19848
rect 10968 19796 11020 19848
rect 19340 19728 19392 19780
rect 5356 19660 5408 19712
rect 5540 19660 5592 19712
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 2780 19456 2832 19508
rect 3976 19456 4028 19508
rect 2688 19252 2740 19304
rect 4712 19252 4764 19304
rect 4988 19252 5040 19304
rect 6920 19252 6972 19304
rect 11060 19320 11112 19372
rect 11244 19320 11296 19372
rect 7288 19252 7340 19304
rect 2228 19184 2280 19236
rect 1768 19159 1820 19168
rect 1768 19125 1777 19159
rect 1777 19125 1811 19159
rect 1811 19125 1820 19159
rect 1768 19116 1820 19125
rect 3332 19184 3384 19236
rect 5724 19184 5776 19236
rect 6644 19184 6696 19236
rect 9588 19252 9640 19304
rect 11888 19252 11940 19304
rect 9404 19184 9456 19236
rect 10968 19184 11020 19236
rect 14004 19252 14056 19304
rect 16028 19295 16080 19304
rect 3424 19116 3476 19168
rect 3608 19116 3660 19168
rect 6460 19159 6512 19168
rect 6460 19125 6469 19159
rect 6469 19125 6503 19159
rect 6503 19125 6512 19159
rect 6460 19116 6512 19125
rect 8208 19116 8260 19168
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 11060 19116 11112 19168
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 12532 19116 12584 19168
rect 13268 19184 13320 19236
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 16580 19295 16632 19304
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 16856 19252 16908 19304
rect 17224 19252 17276 19304
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 18696 19252 18748 19304
rect 15752 19184 15804 19236
rect 22100 19184 22152 19236
rect 16120 19116 16172 19168
rect 17040 19116 17092 19168
rect 17500 19116 17552 19168
rect 18512 19116 18564 19168
rect 18880 19116 18932 19168
rect 20260 19116 20312 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 2872 18912 2924 18964
rect 3332 18955 3384 18964
rect 3332 18921 3341 18955
rect 3341 18921 3375 18955
rect 3375 18921 3384 18955
rect 3332 18912 3384 18921
rect 4068 18912 4120 18964
rect 5448 18912 5500 18964
rect 5724 18912 5776 18964
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 8208 18844 8260 18896
rect 3608 18751 3660 18760
rect 1584 18683 1636 18692
rect 1584 18649 1593 18683
rect 1593 18649 1627 18683
rect 1627 18649 1636 18683
rect 1584 18640 1636 18649
rect 3608 18717 3617 18751
rect 3617 18717 3651 18751
rect 3651 18717 3660 18751
rect 3608 18708 3660 18717
rect 3792 18776 3844 18828
rect 4896 18776 4948 18828
rect 4988 18776 5040 18828
rect 5448 18819 5500 18828
rect 5448 18785 5482 18819
rect 5482 18785 5500 18819
rect 8760 18912 8812 18964
rect 9312 18912 9364 18964
rect 10416 18912 10468 18964
rect 11980 18912 12032 18964
rect 12808 18912 12860 18964
rect 13268 18955 13320 18964
rect 13268 18921 13277 18955
rect 13277 18921 13311 18955
rect 13311 18921 13320 18955
rect 13268 18912 13320 18921
rect 19340 18912 19392 18964
rect 21180 18912 21232 18964
rect 8852 18844 8904 18896
rect 10876 18844 10928 18896
rect 11612 18844 11664 18896
rect 12900 18844 12952 18896
rect 13820 18887 13872 18896
rect 13820 18853 13829 18887
rect 13829 18853 13863 18887
rect 13863 18853 13872 18887
rect 13820 18844 13872 18853
rect 14188 18844 14240 18896
rect 15568 18887 15620 18896
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 18696 18887 18748 18896
rect 18696 18853 18705 18887
rect 18705 18853 18739 18887
rect 18739 18853 18748 18887
rect 18696 18844 18748 18853
rect 5448 18776 5500 18785
rect 4344 18708 4396 18760
rect 3056 18640 3108 18692
rect 4160 18572 4212 18624
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 7288 18751 7340 18760
rect 4620 18708 4672 18717
rect 7288 18717 7297 18751
rect 7297 18717 7331 18751
rect 7331 18717 7340 18751
rect 7288 18708 7340 18717
rect 5080 18640 5132 18692
rect 4896 18572 4948 18624
rect 11060 18776 11112 18828
rect 11152 18776 11204 18828
rect 11888 18819 11940 18828
rect 9588 18708 9640 18760
rect 11888 18785 11897 18819
rect 11897 18785 11931 18819
rect 11931 18785 11940 18819
rect 11888 18776 11940 18785
rect 12992 18776 13044 18828
rect 13084 18776 13136 18828
rect 15292 18819 15344 18828
rect 11796 18708 11848 18760
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 17960 18776 18012 18828
rect 15568 18708 15620 18760
rect 9404 18572 9456 18624
rect 11152 18572 11204 18624
rect 19800 18572 19852 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 204 18368 256 18420
rect 2596 18368 2648 18420
rect 2780 18368 2832 18420
rect 1676 18343 1728 18352
rect 1676 18309 1685 18343
rect 1685 18309 1719 18343
rect 1719 18309 1728 18343
rect 1676 18300 1728 18309
rect 2320 18300 2372 18352
rect 3056 18300 3108 18352
rect 4712 18368 4764 18420
rect 5080 18368 5132 18420
rect 8484 18368 8536 18420
rect 8576 18368 8628 18420
rect 21640 18368 21692 18420
rect 6368 18343 6420 18352
rect 6368 18309 6377 18343
rect 6377 18309 6411 18343
rect 6411 18309 6420 18343
rect 6368 18300 6420 18309
rect 6460 18300 6512 18352
rect 2688 18232 2740 18284
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 7012 18232 7064 18284
rect 8300 18300 8352 18352
rect 8852 18275 8904 18284
rect 8852 18241 8861 18275
rect 8861 18241 8895 18275
rect 8895 18241 8904 18275
rect 8852 18232 8904 18241
rect 2228 18096 2280 18148
rect 3332 18028 3384 18080
rect 4068 18164 4120 18216
rect 4160 18164 4212 18216
rect 7196 18164 7248 18216
rect 9680 18300 9732 18352
rect 11704 18300 11756 18352
rect 9404 18232 9456 18284
rect 11520 18275 11572 18284
rect 11520 18241 11529 18275
rect 11529 18241 11563 18275
rect 11563 18241 11572 18275
rect 11520 18232 11572 18241
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13820 18232 13872 18284
rect 10692 18164 10744 18216
rect 6644 18096 6696 18148
rect 4896 18028 4948 18080
rect 5080 18028 5132 18080
rect 8300 18096 8352 18148
rect 10232 18096 10284 18148
rect 13176 18164 13228 18216
rect 7196 18071 7248 18080
rect 7196 18037 7205 18071
rect 7205 18037 7239 18071
rect 7239 18037 7248 18071
rect 7196 18028 7248 18037
rect 7748 18028 7800 18080
rect 8760 18028 8812 18080
rect 9220 18028 9272 18080
rect 10784 18028 10836 18080
rect 12348 18028 12400 18080
rect 12532 18028 12584 18080
rect 12900 18071 12952 18080
rect 12900 18037 12909 18071
rect 12909 18037 12943 18071
rect 12943 18037 12952 18071
rect 12900 18028 12952 18037
rect 13728 18028 13780 18080
rect 14096 18028 14148 18080
rect 19432 18028 19484 18080
rect 22560 18028 22612 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 3516 17824 3568 17876
rect 6644 17824 6696 17876
rect 7196 17824 7248 17876
rect 7564 17824 7616 17876
rect 11428 17824 11480 17876
rect 2228 17731 2280 17740
rect 2228 17697 2237 17731
rect 2237 17697 2271 17731
rect 2271 17697 2280 17731
rect 2228 17688 2280 17697
rect 2964 17731 3016 17740
rect 2964 17697 2973 17731
rect 2973 17697 3007 17731
rect 3007 17697 3016 17731
rect 2964 17688 3016 17697
rect 4160 17688 4212 17740
rect 4712 17688 4764 17740
rect 5816 17688 5868 17740
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 8576 17756 8628 17808
rect 13820 17824 13872 17876
rect 20628 17824 20680 17876
rect 7748 17731 7800 17740
rect 7748 17697 7782 17731
rect 7782 17697 7800 17731
rect 7748 17688 7800 17697
rect 1400 17620 1452 17672
rect 2596 17484 2648 17536
rect 3148 17484 3200 17536
rect 3332 17620 3384 17672
rect 7196 17620 7248 17672
rect 7288 17620 7340 17672
rect 3700 17552 3752 17604
rect 4068 17552 4120 17604
rect 5540 17552 5592 17604
rect 5448 17527 5500 17536
rect 5448 17493 5457 17527
rect 5457 17493 5491 17527
rect 5491 17493 5500 17527
rect 5448 17484 5500 17493
rect 7104 17484 7156 17536
rect 10968 17688 11020 17740
rect 11704 17688 11756 17740
rect 8944 17620 8996 17672
rect 9772 17552 9824 17604
rect 10508 17620 10560 17672
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 18512 17620 18564 17672
rect 12164 17552 12216 17604
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 9864 17484 9916 17536
rect 13820 17484 13872 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 1584 17119 1636 17128
rect 1584 17085 1593 17119
rect 1593 17085 1627 17119
rect 1627 17085 1636 17119
rect 1584 17076 1636 17085
rect 2688 17212 2740 17264
rect 4712 17323 4764 17332
rect 4712 17289 4721 17323
rect 4721 17289 4755 17323
rect 4755 17289 4764 17323
rect 4712 17280 4764 17289
rect 5540 17280 5592 17332
rect 6184 17280 6236 17332
rect 2964 17144 3016 17196
rect 6736 17212 6788 17264
rect 9864 17280 9916 17332
rect 10048 17255 10100 17264
rect 10048 17221 10057 17255
rect 10057 17221 10091 17255
rect 10091 17221 10100 17255
rect 10048 17212 10100 17221
rect 10968 17280 11020 17332
rect 11704 17323 11756 17332
rect 11704 17289 11713 17323
rect 11713 17289 11747 17323
rect 11747 17289 11756 17323
rect 11704 17280 11756 17289
rect 11888 17280 11940 17332
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 13912 17280 13964 17332
rect 19340 17280 19392 17332
rect 12624 17212 12676 17264
rect 4252 17076 4304 17128
rect 3608 17008 3660 17060
rect 4160 17008 4212 17060
rect 1676 16940 1728 16992
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5356 16940 5408 16992
rect 6368 17076 6420 17128
rect 6000 16940 6052 16992
rect 6276 16940 6328 16992
rect 7196 17008 7248 17060
rect 7656 17008 7708 17060
rect 9772 17076 9824 17128
rect 11704 17144 11756 17196
rect 9864 17008 9916 17060
rect 7288 16940 7340 16992
rect 7380 16940 7432 16992
rect 7748 16940 7800 16992
rect 8484 16940 8536 16992
rect 11796 17076 11848 17128
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 14280 17144 14332 17196
rect 13452 17119 13504 17128
rect 11152 17008 11204 17060
rect 13452 17085 13461 17119
rect 13461 17085 13495 17119
rect 13495 17085 13504 17119
rect 13452 17076 13504 17085
rect 10968 16940 11020 16992
rect 11244 16940 11296 16992
rect 11888 16940 11940 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 12992 16940 13044 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2228 16736 2280 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 4896 16736 4948 16788
rect 5356 16736 5408 16788
rect 1584 16668 1636 16720
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 5080 16668 5132 16720
rect 6828 16736 6880 16788
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 10140 16736 10192 16788
rect 10876 16736 10928 16788
rect 11244 16736 11296 16788
rect 11612 16736 11664 16788
rect 8484 16711 8536 16720
rect 8484 16677 8493 16711
rect 8493 16677 8527 16711
rect 8527 16677 8536 16711
rect 8484 16668 8536 16677
rect 11152 16668 11204 16720
rect 13452 16668 13504 16720
rect 3424 16600 3476 16652
rect 4160 16600 4212 16652
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 2964 16464 3016 16516
rect 3792 16464 3844 16516
rect 4068 16464 4120 16516
rect 572 16396 624 16448
rect 4160 16396 4212 16448
rect 7564 16600 7616 16652
rect 11244 16600 11296 16652
rect 12348 16600 12400 16652
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 7656 16507 7708 16516
rect 7656 16473 7665 16507
rect 7665 16473 7699 16507
rect 7699 16473 7708 16507
rect 9220 16532 9272 16584
rect 10508 16575 10560 16584
rect 7656 16464 7708 16473
rect 9588 16464 9640 16516
rect 10140 16464 10192 16516
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 11704 16532 11756 16584
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 11796 16464 11848 16516
rect 13636 16464 13688 16516
rect 7748 16396 7800 16448
rect 8208 16396 8260 16448
rect 9128 16396 9180 16448
rect 12256 16396 12308 16448
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 6828 16192 6880 16244
rect 7196 16192 7248 16244
rect 8208 16192 8260 16244
rect 8300 16192 8352 16244
rect 14280 16192 14332 16244
rect 1032 16124 1084 16176
rect 3424 16124 3476 16176
rect 4252 16124 4304 16176
rect 3700 16056 3752 16108
rect 4712 16056 4764 16108
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 2964 15988 3016 16040
rect 3240 15988 3292 16040
rect 7564 16056 7616 16108
rect 9312 16056 9364 16108
rect 6184 16031 6236 16040
rect 1768 15920 1820 15972
rect 1952 15895 2004 15904
rect 1952 15861 1961 15895
rect 1961 15861 1995 15895
rect 1995 15861 2004 15895
rect 1952 15852 2004 15861
rect 2872 15920 2924 15972
rect 3424 15963 3476 15972
rect 3424 15929 3433 15963
rect 3433 15929 3467 15963
rect 3467 15929 3476 15963
rect 3424 15920 3476 15929
rect 3976 15920 4028 15972
rect 6184 15997 6193 16031
rect 6193 15997 6227 16031
rect 6227 15997 6236 16031
rect 6184 15988 6236 15997
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 9588 16056 9640 16108
rect 10048 16056 10100 16108
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 9956 15988 10008 16040
rect 10232 15988 10284 16040
rect 11796 16056 11848 16108
rect 13820 16056 13872 16108
rect 11428 16031 11480 16040
rect 11428 15997 11437 16031
rect 11437 15997 11471 16031
rect 11471 15997 11480 16031
rect 11428 15988 11480 15997
rect 11704 15988 11756 16040
rect 6276 15920 6328 15972
rect 3608 15852 3660 15904
rect 4068 15852 4120 15904
rect 4896 15852 4948 15904
rect 5448 15852 5500 15904
rect 5908 15852 5960 15904
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 9680 15920 9732 15972
rect 13912 15920 13964 15972
rect 9864 15852 9916 15904
rect 10784 15852 10836 15904
rect 11980 15852 12032 15904
rect 12900 15895 12952 15904
rect 12900 15861 12909 15895
rect 12909 15861 12943 15895
rect 12943 15861 12952 15895
rect 12900 15852 12952 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 1952 15648 2004 15700
rect 1676 15512 1728 15564
rect 2412 15555 2464 15564
rect 2412 15521 2421 15555
rect 2421 15521 2455 15555
rect 2455 15521 2464 15555
rect 2412 15512 2464 15521
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 4528 15648 4580 15657
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 6276 15648 6328 15700
rect 6736 15691 6788 15700
rect 6736 15657 6745 15691
rect 6745 15657 6779 15691
rect 6779 15657 6788 15691
rect 6736 15648 6788 15657
rect 7104 15691 7156 15700
rect 7104 15657 7113 15691
rect 7113 15657 7147 15691
rect 7147 15657 7156 15691
rect 7104 15648 7156 15657
rect 7748 15648 7800 15700
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 10692 15648 10744 15700
rect 11704 15648 11756 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 12900 15648 12952 15700
rect 8300 15580 8352 15632
rect 10416 15580 10468 15632
rect 13268 15580 13320 15632
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 8208 15555 8260 15564
rect 3148 15444 3200 15496
rect 3700 15444 3752 15496
rect 8208 15521 8231 15555
rect 8231 15521 8260 15555
rect 9680 15555 9732 15564
rect 8208 15512 8260 15521
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 12716 15512 12768 15564
rect 13820 15512 13872 15564
rect 14556 15512 14608 15564
rect 4896 15444 4948 15496
rect 5356 15444 5408 15496
rect 6828 15444 6880 15496
rect 7380 15487 7432 15496
rect 7380 15453 7389 15487
rect 7389 15453 7423 15487
rect 7423 15453 7432 15487
rect 7380 15444 7432 15453
rect 12624 15487 12676 15496
rect 4160 15308 4212 15360
rect 5448 15308 5500 15360
rect 7288 15376 7340 15428
rect 12624 15453 12633 15487
rect 12633 15453 12667 15487
rect 12667 15453 12676 15487
rect 12624 15444 12676 15453
rect 12348 15376 12400 15428
rect 10784 15308 10836 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 3424 15147 3476 15156
rect 3424 15113 3433 15147
rect 3433 15113 3467 15147
rect 3467 15113 3476 15147
rect 3424 15104 3476 15113
rect 5080 15104 5132 15156
rect 5724 15147 5776 15156
rect 5724 15113 5733 15147
rect 5733 15113 5767 15147
rect 5767 15113 5776 15147
rect 5724 15104 5776 15113
rect 6368 15104 6420 15156
rect 9864 15104 9916 15156
rect 12716 15104 12768 15156
rect 15016 15147 15068 15156
rect 15016 15113 15025 15147
rect 15025 15113 15059 15147
rect 15059 15113 15068 15147
rect 15016 15104 15068 15113
rect 5264 15036 5316 15088
rect 8208 15079 8260 15088
rect 8208 15045 8217 15079
rect 8217 15045 8251 15079
rect 8251 15045 8260 15079
rect 8208 15036 8260 15045
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 1768 14968 1820 15020
rect 3056 14968 3108 15020
rect 3976 14968 4028 15020
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 3700 14900 3752 14952
rect 6276 14900 6328 14952
rect 4160 14832 4212 14884
rect 4896 14832 4948 14884
rect 6736 14900 6788 14952
rect 8208 14900 8260 14952
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 9588 15036 9640 15088
rect 9956 15036 10008 15088
rect 11612 15036 11664 15088
rect 9312 14968 9364 15020
rect 9772 14968 9824 15020
rect 10232 14900 10284 14952
rect 13084 14968 13136 15020
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 13820 14968 13872 15020
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 15936 14968 15988 15020
rect 7288 14832 7340 14884
rect 7380 14832 7432 14884
rect 10692 14832 10744 14884
rect 2688 14807 2740 14816
rect 2688 14773 2697 14807
rect 2697 14773 2731 14807
rect 2731 14773 2740 14807
rect 2688 14764 2740 14773
rect 3148 14764 3200 14816
rect 8484 14764 8536 14816
rect 9312 14764 9364 14816
rect 9680 14764 9732 14816
rect 9772 14764 9824 14816
rect 12256 14900 12308 14952
rect 13636 14900 13688 14952
rect 14372 14943 14424 14952
rect 14372 14909 14381 14943
rect 14381 14909 14415 14943
rect 14415 14909 14424 14943
rect 14372 14900 14424 14909
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 15384 14875 15436 14884
rect 15384 14841 15393 14875
rect 15393 14841 15427 14875
rect 15427 14841 15436 14875
rect 15384 14832 15436 14841
rect 12900 14764 12952 14816
rect 18604 14764 18656 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 9956 14560 10008 14612
rect 15476 14560 15528 14612
rect 4252 14492 4304 14544
rect 5908 14492 5960 14544
rect 6000 14492 6052 14544
rect 7380 14492 7432 14544
rect 10968 14492 11020 14544
rect 11704 14492 11756 14544
rect 13544 14492 13596 14544
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2136 14424 2188 14476
rect 4712 14424 4764 14476
rect 6276 14424 6328 14476
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 3056 14288 3108 14340
rect 5356 14356 5408 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 7840 14424 7892 14476
rect 8300 14424 8352 14476
rect 9772 14424 9824 14476
rect 10876 14467 10928 14476
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 8208 14356 8260 14408
rect 9404 14356 9456 14408
rect 7564 14288 7616 14340
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 10876 14433 10885 14467
rect 10885 14433 10919 14467
rect 10919 14433 10928 14467
rect 10876 14424 10928 14433
rect 12440 14424 12492 14476
rect 12900 14424 12952 14476
rect 13820 14424 13872 14476
rect 19432 14560 19484 14612
rect 11060 14356 11112 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 12256 14288 12308 14340
rect 4068 14263 4120 14272
rect 4068 14229 4077 14263
rect 4077 14229 4111 14263
rect 4111 14229 4120 14263
rect 4068 14220 4120 14229
rect 4712 14220 4764 14272
rect 5172 14220 5224 14272
rect 8392 14220 8444 14272
rect 8484 14220 8536 14272
rect 10416 14220 10468 14272
rect 11060 14220 11112 14272
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 14556 14288 14608 14340
rect 14004 14220 14056 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1768 14016 1820 14068
rect 2044 14016 2096 14068
rect 3700 14016 3752 14068
rect 4896 14016 4948 14068
rect 7656 14016 7708 14068
rect 7840 14059 7892 14068
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 9404 14016 9456 14068
rect 13820 14059 13872 14068
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 4344 13948 4396 14000
rect 3608 13880 3660 13932
rect 4068 13880 4120 13932
rect 6276 13948 6328 14000
rect 8668 13948 8720 14000
rect 10876 13948 10928 14000
rect 11796 13948 11848 14000
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 7656 13880 7708 13932
rect 8944 13880 8996 13932
rect 9864 13880 9916 13932
rect 10232 13880 10284 13932
rect 10416 13880 10468 13932
rect 11704 13880 11756 13932
rect 12072 13880 12124 13932
rect 1400 13812 1452 13864
rect 3056 13812 3108 13864
rect 4160 13812 4212 13864
rect 5448 13812 5500 13864
rect 6368 13855 6420 13864
rect 6368 13821 6377 13855
rect 6377 13821 6411 13855
rect 6411 13821 6420 13855
rect 6368 13812 6420 13821
rect 6920 13812 6972 13864
rect 9404 13812 9456 13864
rect 3424 13744 3476 13796
rect 3792 13744 3844 13796
rect 10876 13812 10928 13864
rect 11060 13812 11112 13864
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 12992 13812 13044 13864
rect 18696 13812 18748 13864
rect 3148 13676 3200 13728
rect 3884 13676 3936 13728
rect 5356 13676 5408 13728
rect 5816 13676 5868 13728
rect 6736 13676 6788 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 7472 13676 7524 13728
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 9864 13676 9916 13728
rect 11520 13676 11572 13728
rect 12440 13676 12492 13728
rect 12808 13676 12860 13728
rect 15936 13744 15988 13796
rect 15016 13676 15068 13728
rect 16028 13676 16080 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 2688 13472 2740 13524
rect 3332 13515 3384 13524
rect 3332 13481 3341 13515
rect 3341 13481 3375 13515
rect 3375 13481 3384 13515
rect 3332 13472 3384 13481
rect 5724 13472 5776 13524
rect 7748 13472 7800 13524
rect 8852 13472 8904 13524
rect 10508 13472 10560 13524
rect 10600 13472 10652 13524
rect 10876 13472 10928 13524
rect 11796 13472 11848 13524
rect 14556 13472 14608 13524
rect 15016 13472 15068 13524
rect 15108 13472 15160 13524
rect 16672 13515 16724 13524
rect 1492 13404 1544 13456
rect 2320 13336 2372 13388
rect 2872 13336 2924 13388
rect 2136 13268 2188 13320
rect 3424 13404 3476 13456
rect 4068 13404 4120 13456
rect 4344 13447 4396 13456
rect 4344 13413 4378 13447
rect 4378 13413 4396 13447
rect 4344 13404 4396 13413
rect 3884 13336 3936 13388
rect 5816 13336 5868 13388
rect 6000 13379 6052 13388
rect 6000 13345 6034 13379
rect 6034 13345 6052 13379
rect 9772 13404 9824 13456
rect 16672 13481 16681 13515
rect 16681 13481 16715 13515
rect 16715 13481 16724 13515
rect 16672 13472 16724 13481
rect 6000 13336 6052 13345
rect 7104 13336 7156 13388
rect 7656 13379 7708 13388
rect 7656 13345 7690 13379
rect 7690 13345 7708 13379
rect 7656 13336 7708 13345
rect 7932 13336 7984 13388
rect 3700 13200 3752 13252
rect 6736 13268 6788 13320
rect 9680 13336 9732 13388
rect 10784 13336 10836 13388
rect 11704 13336 11756 13388
rect 11796 13336 11848 13388
rect 10048 13311 10100 13320
rect 10048 13277 10057 13311
rect 10057 13277 10091 13311
rect 10091 13277 10100 13311
rect 10048 13268 10100 13277
rect 10232 13268 10284 13320
rect 3608 13132 3660 13184
rect 9956 13200 10008 13252
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 12900 13336 12952 13388
rect 13544 13336 13596 13388
rect 14188 13336 14240 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 11244 13268 11296 13277
rect 12532 13268 12584 13320
rect 14556 13268 14608 13320
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 12808 13200 12860 13252
rect 15016 13200 15068 13252
rect 10048 13132 10100 13184
rect 10692 13132 10744 13184
rect 13728 13132 13780 13184
rect 14924 13132 14976 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 3424 12928 3476 12980
rect 3700 12928 3752 12980
rect 3976 12971 4028 12980
rect 3976 12937 3985 12971
rect 3985 12937 4019 12971
rect 4019 12937 4028 12971
rect 3976 12928 4028 12937
rect 3148 12860 3200 12912
rect 5816 12928 5868 12980
rect 6000 12971 6052 12980
rect 6000 12937 6009 12971
rect 6009 12937 6043 12971
rect 6043 12937 6052 12971
rect 6000 12928 6052 12937
rect 7288 12928 7340 12980
rect 7380 12928 7432 12980
rect 9680 12971 9732 12980
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 3700 12792 3752 12844
rect 6736 12860 6788 12912
rect 9680 12937 9689 12971
rect 9689 12937 9723 12971
rect 9723 12937 9732 12971
rect 9680 12928 9732 12937
rect 10232 12928 10284 12980
rect 12072 12971 12124 12980
rect 6276 12792 6328 12844
rect 7656 12792 7708 12844
rect 7748 12792 7800 12844
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 12256 12928 12308 12980
rect 12624 12928 12676 12980
rect 17132 12928 17184 12980
rect 14280 12903 14332 12912
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 5724 12724 5776 12776
rect 6828 12724 6880 12776
rect 11704 12792 11756 12844
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 14280 12869 14289 12903
rect 14289 12869 14323 12903
rect 14323 12869 14332 12903
rect 14280 12860 14332 12869
rect 14188 12792 14240 12844
rect 15108 12835 15160 12844
rect 15108 12801 15117 12835
rect 15117 12801 15151 12835
rect 15151 12801 15160 12835
rect 15108 12792 15160 12801
rect 4988 12656 5040 12708
rect 7012 12656 7064 12708
rect 8944 12656 8996 12708
rect 10232 12656 10284 12708
rect 11244 12656 11296 12708
rect 12440 12656 12492 12708
rect 13820 12656 13872 12708
rect 1584 12588 1636 12640
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 2780 12631 2832 12640
rect 2780 12597 2789 12631
rect 2789 12597 2823 12631
rect 2823 12597 2832 12631
rect 2780 12588 2832 12597
rect 5908 12588 5960 12640
rect 7380 12588 7432 12640
rect 7748 12588 7800 12640
rect 11428 12588 11480 12640
rect 11980 12588 12032 12640
rect 14556 12724 14608 12776
rect 14924 12767 14976 12776
rect 14924 12733 14933 12767
rect 14933 12733 14967 12767
rect 14967 12733 14976 12767
rect 14924 12724 14976 12733
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 15016 12588 15068 12640
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2136 12384 2188 12436
rect 3148 12427 3200 12436
rect 3148 12393 3157 12427
rect 3157 12393 3191 12427
rect 3191 12393 3200 12427
rect 3148 12384 3200 12393
rect 3332 12384 3384 12436
rect 4252 12384 4304 12436
rect 4804 12384 4856 12436
rect 4160 12316 4212 12368
rect 5724 12384 5776 12436
rect 6552 12384 6604 12436
rect 6920 12384 6972 12436
rect 8944 12427 8996 12436
rect 8944 12393 8953 12427
rect 8953 12393 8987 12427
rect 8987 12393 8996 12427
rect 8944 12384 8996 12393
rect 9588 12384 9640 12436
rect 9680 12384 9732 12436
rect 10876 12384 10928 12436
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 12348 12427 12400 12436
rect 12348 12393 12357 12427
rect 12357 12393 12391 12427
rect 12391 12393 12400 12427
rect 12348 12384 12400 12393
rect 14188 12384 14240 12436
rect 14556 12384 14608 12436
rect 9128 12316 9180 12368
rect 10048 12316 10100 12368
rect 2780 12248 2832 12300
rect 3332 12248 3384 12300
rect 3976 12248 4028 12300
rect 2504 12180 2556 12232
rect 3700 12180 3752 12232
rect 1860 12112 1912 12164
rect 5816 12248 5868 12300
rect 6184 12291 6236 12300
rect 6184 12257 6218 12291
rect 6218 12257 6236 12291
rect 6184 12248 6236 12257
rect 7748 12248 7800 12300
rect 8484 12248 8536 12300
rect 10600 12316 10652 12368
rect 10692 12316 10744 12368
rect 11060 12248 11112 12300
rect 13912 12316 13964 12368
rect 12532 12248 12584 12300
rect 7656 12180 7708 12232
rect 9680 12223 9732 12232
rect 9680 12189 9689 12223
rect 9689 12189 9723 12223
rect 9723 12189 9732 12223
rect 9680 12180 9732 12189
rect 9772 12180 9824 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 13084 12223 13136 12232
rect 4896 12044 4948 12096
rect 5448 12044 5500 12096
rect 10140 12112 10192 12164
rect 11244 12112 11296 12164
rect 7380 12044 7432 12096
rect 11152 12044 11204 12096
rect 13084 12189 13093 12223
rect 13093 12189 13127 12223
rect 13127 12189 13136 12223
rect 13084 12180 13136 12189
rect 13912 12044 13964 12096
rect 14464 12044 14516 12096
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2504 11840 2556 11892
rect 4988 11883 5040 11892
rect 4988 11849 4997 11883
rect 4997 11849 5031 11883
rect 5031 11849 5040 11883
rect 4988 11840 5040 11849
rect 5080 11840 5132 11892
rect 12348 11840 12400 11892
rect 13360 11840 13412 11892
rect 14924 11840 14976 11892
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 4896 11704 4948 11756
rect 8668 11772 8720 11824
rect 5908 11704 5960 11756
rect 9312 11704 9364 11756
rect 9404 11704 9456 11756
rect 1584 11679 1636 11688
rect 1584 11645 1593 11679
rect 1593 11645 1627 11679
rect 1627 11645 1636 11679
rect 1584 11636 1636 11645
rect 2044 11636 2096 11688
rect 3700 11636 3752 11688
rect 5448 11568 5500 11620
rect 8208 11636 8260 11688
rect 10968 11636 11020 11688
rect 11060 11636 11112 11688
rect 12348 11704 12400 11756
rect 12440 11747 12492 11756
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 14648 11747 14700 11756
rect 12440 11704 12492 11713
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 17224 11704 17276 11756
rect 11888 11636 11940 11688
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 4436 11543 4488 11552
rect 4436 11509 4445 11543
rect 4445 11509 4479 11543
rect 4479 11509 4488 11543
rect 4436 11500 4488 11509
rect 6920 11500 6972 11552
rect 7288 11500 7340 11552
rect 8208 11500 8260 11552
rect 8484 11568 8536 11620
rect 10876 11568 10928 11620
rect 11244 11611 11296 11620
rect 11244 11577 11253 11611
rect 11253 11577 11287 11611
rect 11287 11577 11296 11611
rect 11244 11568 11296 11577
rect 12808 11568 12860 11620
rect 13084 11636 13136 11688
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 8852 11500 8904 11552
rect 9496 11500 9548 11552
rect 12348 11500 12400 11552
rect 12532 11500 12584 11552
rect 12624 11500 12676 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14280 11500 14332 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2412 11296 2464 11348
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 4436 11296 4488 11348
rect 5264 11296 5316 11348
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 7012 11296 7064 11348
rect 2504 11228 2556 11280
rect 3792 11228 3844 11280
rect 2044 11160 2096 11212
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 5816 11160 5868 11212
rect 4804 11135 4856 11144
rect 4804 11101 4813 11135
rect 4813 11101 4847 11135
rect 4847 11101 4856 11135
rect 4804 11092 4856 11101
rect 4344 11024 4396 11076
rect 6920 11160 6972 11212
rect 7012 11160 7064 11212
rect 7656 11160 7708 11212
rect 6736 11092 6788 11144
rect 10232 11296 10284 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 12440 11296 12492 11348
rect 16672 11296 16724 11348
rect 8484 11228 8536 11280
rect 8576 11228 8628 11280
rect 9312 11228 9364 11280
rect 11152 11228 11204 11280
rect 12532 11228 12584 11280
rect 8944 11160 8996 11212
rect 9128 11160 9180 11212
rect 9404 11160 9456 11212
rect 9772 11160 9824 11212
rect 13176 11203 13228 11212
rect 11060 11092 11112 11144
rect 12348 11092 12400 11144
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 14464 11203 14516 11212
rect 7196 11024 7248 11076
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 12624 11092 12676 11144
rect 6276 10956 6328 11008
rect 9680 10956 9732 11008
rect 11980 10999 12032 11008
rect 11980 10965 11989 10999
rect 11989 10965 12023 10999
rect 12023 10965 12032 10999
rect 11980 10956 12032 10965
rect 12164 10956 12216 11008
rect 12900 11024 12952 11076
rect 14464 11169 14473 11203
rect 14473 11169 14507 11203
rect 14507 11169 14516 11203
rect 14464 11160 14516 11169
rect 14556 11135 14608 11144
rect 14556 11101 14565 11135
rect 14565 11101 14599 11135
rect 14599 11101 14608 11135
rect 14556 11092 14608 11101
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 16856 11024 16908 11076
rect 13084 10956 13136 11008
rect 16580 10956 16632 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 4712 10752 4764 10804
rect 7472 10752 7524 10804
rect 5816 10727 5868 10736
rect 5816 10693 5825 10727
rect 5825 10693 5859 10727
rect 5859 10693 5868 10727
rect 8852 10752 8904 10804
rect 9956 10752 10008 10804
rect 10140 10752 10192 10804
rect 8944 10727 8996 10736
rect 5816 10684 5868 10693
rect 6736 10616 6788 10668
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 6276 10591 6328 10600
rect 2412 10480 2464 10532
rect 4620 10480 4672 10532
rect 4804 10480 4856 10532
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 6276 10548 6328 10557
rect 6368 10548 6420 10600
rect 8668 10548 8720 10600
rect 8944 10693 8953 10727
rect 8953 10693 8987 10727
rect 8987 10693 8996 10727
rect 8944 10684 8996 10693
rect 9312 10684 9364 10736
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 12348 10752 12400 10804
rect 12440 10795 12492 10804
rect 12440 10761 12449 10795
rect 12449 10761 12483 10795
rect 12483 10761 12492 10795
rect 12440 10752 12492 10761
rect 14464 10752 14516 10804
rect 10232 10684 10284 10693
rect 13820 10684 13872 10736
rect 9312 10548 9364 10600
rect 9404 10548 9456 10600
rect 9864 10548 9916 10600
rect 13360 10616 13412 10668
rect 15016 10684 15068 10736
rect 15108 10616 15160 10668
rect 5080 10480 5132 10532
rect 5632 10412 5684 10464
rect 6276 10412 6328 10464
rect 6920 10412 6972 10464
rect 8300 10412 8352 10464
rect 10140 10480 10192 10532
rect 11060 10480 11112 10532
rect 14280 10548 14332 10600
rect 10324 10412 10376 10464
rect 12716 10412 12768 10464
rect 13084 10412 13136 10464
rect 13820 10412 13872 10464
rect 14372 10412 14424 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 3240 10208 3292 10260
rect 3700 10251 3752 10260
rect 3700 10217 3709 10251
rect 3709 10217 3743 10251
rect 3743 10217 3752 10251
rect 3700 10208 3752 10217
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 10324 10208 10376 10260
rect 12900 10208 12952 10260
rect 14372 10208 14424 10260
rect 8852 10140 8904 10192
rect 2872 10072 2924 10124
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 5632 10072 5684 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6460 10072 6512 10124
rect 6644 10115 6696 10124
rect 6644 10081 6678 10115
rect 6678 10081 6696 10115
rect 6644 10072 6696 10081
rect 6920 10072 6972 10124
rect 9404 10072 9456 10124
rect 2044 10004 2096 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5172 10004 5224 10056
rect 5816 10004 5868 10056
rect 8300 10004 8352 10056
rect 8944 10004 8996 10056
rect 5632 9936 5684 9988
rect 7472 9936 7524 9988
rect 9772 10140 9824 10192
rect 9956 10183 10008 10192
rect 9956 10149 9990 10183
rect 9990 10149 10008 10183
rect 9956 10140 10008 10149
rect 10140 10140 10192 10192
rect 10232 10072 10284 10124
rect 12348 10140 12400 10192
rect 12900 10072 12952 10124
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 12440 10004 12492 10056
rect 12716 10004 12768 10056
rect 13176 10004 13228 10056
rect 14096 10004 14148 10056
rect 4068 9911 4120 9920
rect 4068 9877 4077 9911
rect 4077 9877 4111 9911
rect 4111 9877 4120 9911
rect 4068 9868 4120 9877
rect 7656 9868 7708 9920
rect 8668 9868 8720 9920
rect 9404 9868 9456 9920
rect 10324 9868 10376 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 12716 9868 12768 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3976 9664 4028 9716
rect 10416 9664 10468 9716
rect 3056 9596 3108 9648
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 2688 9460 2740 9512
rect 3424 9460 3476 9512
rect 5264 9460 5316 9512
rect 5816 9528 5868 9580
rect 7012 9528 7064 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 2320 9367 2372 9376
rect 2320 9333 2329 9367
rect 2329 9333 2363 9367
rect 2363 9333 2372 9367
rect 2320 9324 2372 9333
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 4160 9392 4212 9444
rect 5172 9392 5224 9444
rect 4712 9324 4764 9376
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 5632 9392 5684 9444
rect 7288 9435 7340 9444
rect 7288 9401 7297 9435
rect 7297 9401 7331 9435
rect 7331 9401 7340 9435
rect 7288 9392 7340 9401
rect 7104 9324 7156 9376
rect 8300 9596 8352 9648
rect 10600 9639 10652 9648
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 11060 9664 11112 9716
rect 16764 9664 16816 9716
rect 10600 9596 10652 9605
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 9956 9528 10008 9580
rect 11704 9596 11756 9648
rect 11888 9596 11940 9648
rect 12532 9596 12584 9648
rect 12716 9596 12768 9648
rect 17960 9596 18012 9648
rect 13636 9528 13688 9580
rect 9496 9460 9548 9512
rect 9680 9460 9732 9512
rect 10600 9460 10652 9512
rect 10876 9392 10928 9444
rect 8300 9324 8352 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 8760 9324 8812 9376
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 10140 9324 10192 9376
rect 11520 9324 11572 9376
rect 14096 9528 14148 9580
rect 14188 9460 14240 9512
rect 15108 9460 15160 9512
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 14556 9324 14608 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 3424 9120 3476 9172
rect 5540 9120 5592 9172
rect 6736 9120 6788 9172
rect 9956 9120 10008 9172
rect 10416 9120 10468 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11612 9120 11664 9172
rect 2504 9052 2556 9104
rect 7104 9052 7156 9104
rect 11520 9052 11572 9104
rect 12348 9120 12400 9172
rect 13912 9120 13964 9172
rect 14372 9120 14424 9172
rect 1584 8959 1636 8968
rect 1584 8925 1593 8959
rect 1593 8925 1627 8959
rect 1627 8925 1636 8959
rect 1584 8916 1636 8925
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 4160 8984 4212 9036
rect 4436 9027 4488 9036
rect 4436 8993 4445 9027
rect 4445 8993 4479 9027
rect 4479 8993 4488 9027
rect 4436 8984 4488 8993
rect 5080 8984 5132 9036
rect 5264 8984 5316 9036
rect 4620 8959 4672 8968
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 4804 8916 4856 8968
rect 7012 8984 7064 9036
rect 8300 8984 8352 9036
rect 9680 8984 9732 9036
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 8668 8916 8720 8968
rect 3424 8823 3476 8832
rect 3424 8789 3433 8823
rect 3433 8789 3467 8823
rect 3467 8789 3476 8823
rect 3424 8780 3476 8789
rect 5080 8780 5132 8832
rect 6644 8780 6696 8832
rect 9864 8848 9916 8900
rect 7656 8780 7708 8832
rect 7932 8780 7984 8832
rect 9772 8780 9824 8832
rect 10048 8848 10100 8900
rect 10508 8916 10560 8968
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 11428 8848 11480 8900
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 13084 8916 13136 8968
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 13820 8916 13872 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 12440 8848 12492 8900
rect 12624 8848 12676 8900
rect 13452 8848 13504 8900
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2044 8576 2096 8628
rect 2320 8576 2372 8628
rect 3976 8576 4028 8628
rect 2596 8508 2648 8560
rect 3424 8440 3476 8492
rect 4160 8440 4212 8492
rect 4896 8440 4948 8492
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 7380 8576 7432 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 14096 8576 14148 8628
rect 14556 8576 14608 8628
rect 12072 8551 12124 8560
rect 12072 8517 12081 8551
rect 12081 8517 12115 8551
rect 12115 8517 12124 8551
rect 12072 8508 12124 8517
rect 12348 8508 12400 8560
rect 4068 8372 4120 8424
rect 11888 8440 11940 8492
rect 13268 8440 13320 8492
rect 14280 8440 14332 8492
rect 5540 8304 5592 8356
rect 7932 8372 7984 8424
rect 7380 8347 7432 8356
rect 3424 8279 3476 8288
rect 3424 8245 3433 8279
rect 3433 8245 3467 8279
rect 3467 8245 3476 8279
rect 3424 8236 3476 8245
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 4160 8236 4212 8288
rect 4712 8236 4764 8288
rect 5172 8236 5224 8288
rect 7380 8313 7414 8347
rect 7414 8313 7432 8347
rect 7380 8304 7432 8313
rect 10232 8372 10284 8424
rect 14188 8372 14240 8424
rect 10876 8304 10928 8356
rect 11152 8304 11204 8356
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 13728 8304 13780 8356
rect 9128 8236 9180 8288
rect 12164 8236 12216 8288
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 13912 8236 13964 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1584 8032 1636 8084
rect 4344 8032 4396 8084
rect 4988 8032 5040 8084
rect 5540 8032 5592 8084
rect 7288 8032 7340 8084
rect 7656 8032 7708 8084
rect 4068 7964 4120 8016
rect 4804 7964 4856 8016
rect 8300 7964 8352 8016
rect 8392 7964 8444 8016
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3976 7896 4028 7948
rect 5356 7896 5408 7948
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6368 7896 6420 7948
rect 6644 7939 6696 7948
rect 6644 7905 6653 7939
rect 6653 7905 6687 7939
rect 6687 7905 6696 7939
rect 6644 7896 6696 7905
rect 7104 7896 7156 7948
rect 7656 7896 7708 7948
rect 3424 7760 3476 7812
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 4344 7828 4396 7880
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 6184 7828 6236 7880
rect 6736 7828 6788 7880
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 9128 7964 9180 8016
rect 10140 7964 10192 8016
rect 10600 8032 10652 8084
rect 10876 8032 10928 8084
rect 11612 8032 11664 8084
rect 14464 8032 14516 8084
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 10232 7896 10284 7948
rect 11612 7896 11664 7948
rect 9312 7828 9364 7880
rect 13820 7964 13872 8016
rect 12072 7939 12124 7948
rect 12072 7905 12106 7939
rect 12106 7905 12124 7939
rect 13728 7939 13780 7948
rect 12072 7896 12124 7905
rect 13728 7905 13762 7939
rect 13762 7905 13780 7939
rect 13728 7896 13780 7905
rect 13452 7871 13504 7880
rect 4068 7760 4120 7812
rect 4712 7692 4764 7744
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 6276 7735 6328 7744
rect 6276 7701 6285 7735
rect 6285 7701 6319 7735
rect 6319 7701 6328 7735
rect 6276 7692 6328 7701
rect 7564 7692 7616 7744
rect 7932 7692 7984 7744
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 11980 7692 12032 7744
rect 13728 7692 13780 7744
rect 14188 7692 14240 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 3240 7488 3292 7540
rect 5816 7488 5868 7540
rect 7196 7488 7248 7540
rect 6276 7420 6328 7472
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2872 7352 2924 7404
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 1400 7284 1452 7336
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 4712 7284 4764 7336
rect 5080 7216 5132 7268
rect 5448 7284 5500 7336
rect 7656 7352 7708 7404
rect 11612 7420 11664 7472
rect 12900 7488 12952 7540
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 7748 7216 7800 7268
rect 9864 7284 9916 7336
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 10324 7216 10376 7268
rect 12440 7284 12492 7336
rect 15752 7420 15804 7472
rect 13544 7352 13596 7404
rect 13728 7352 13780 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 16948 7352 17000 7404
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 3148 7148 3200 7200
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 6000 7191 6052 7200
rect 3424 7148 3476 7157
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 7196 7148 7248 7200
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 8300 7191 8352 7200
rect 7288 7148 7340 7157
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 10140 7148 10192 7200
rect 12716 7216 12768 7268
rect 12992 7216 13044 7268
rect 13820 7259 13872 7268
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 14372 7216 14424 7268
rect 12532 7148 12584 7200
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13360 7148 13412 7200
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 2964 6944 3016 6996
rect 9588 6944 9640 6996
rect 13084 6987 13136 6996
rect 13084 6953 13093 6987
rect 13093 6953 13127 6987
rect 13127 6953 13136 6987
rect 13084 6944 13136 6953
rect 14280 6944 14332 6996
rect 14464 6944 14516 6996
rect 2136 6876 2188 6928
rect 2688 6876 2740 6928
rect 4896 6876 4948 6928
rect 5908 6876 5960 6928
rect 6368 6876 6420 6928
rect 1768 6808 1820 6860
rect 2964 6808 3016 6860
rect 6000 6808 6052 6860
rect 2688 6740 2740 6792
rect 5356 6740 5408 6792
rect 2872 6672 2924 6724
rect 10048 6876 10100 6928
rect 10692 6876 10744 6928
rect 10968 6876 11020 6928
rect 11060 6876 11112 6928
rect 12348 6876 12400 6928
rect 13360 6876 13412 6928
rect 16580 6876 16632 6928
rect 9680 6851 9732 6860
rect 9680 6817 9689 6851
rect 9689 6817 9723 6851
rect 9723 6817 9732 6851
rect 9680 6808 9732 6817
rect 11152 6808 11204 6860
rect 12900 6808 12952 6860
rect 13728 6808 13780 6860
rect 15016 6808 15068 6860
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 7196 6740 7248 6792
rect 4712 6604 4764 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 8576 6647 8628 6656
rect 8576 6613 8585 6647
rect 8585 6613 8619 6647
rect 8619 6613 8628 6647
rect 8576 6604 8628 6613
rect 11612 6740 11664 6792
rect 12992 6740 13044 6792
rect 13268 6740 13320 6792
rect 10692 6672 10744 6724
rect 11060 6715 11112 6724
rect 11060 6681 11069 6715
rect 11069 6681 11103 6715
rect 11103 6681 11112 6715
rect 11060 6672 11112 6681
rect 13820 6672 13872 6724
rect 10600 6604 10652 6656
rect 12348 6604 12400 6656
rect 13268 6604 13320 6656
rect 14556 6740 14608 6792
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 14280 6672 14332 6724
rect 15108 6672 15160 6724
rect 17132 6672 17184 6724
rect 17316 6604 17368 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2228 6400 2280 6452
rect 3424 6400 3476 6452
rect 7288 6400 7340 6452
rect 8576 6400 8628 6452
rect 12808 6400 12860 6452
rect 13820 6400 13872 6452
rect 15752 6400 15804 6452
rect 4068 6332 4120 6384
rect 7748 6332 7800 6384
rect 9312 6375 9364 6384
rect 9312 6341 9321 6375
rect 9321 6341 9355 6375
rect 9355 6341 9364 6375
rect 9312 6332 9364 6341
rect 3976 6264 4028 6316
rect 6276 6307 6328 6316
rect 4988 6196 5040 6248
rect 5264 6196 5316 6248
rect 6276 6273 6285 6307
rect 6285 6273 6319 6307
rect 6319 6273 6328 6307
rect 6276 6264 6328 6273
rect 6920 6264 6972 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 7380 6196 7432 6248
rect 8024 6196 8076 6248
rect 10508 6196 10560 6248
rect 11152 6264 11204 6316
rect 12072 6264 12124 6316
rect 13636 6196 13688 6248
rect 2504 6128 2556 6180
rect 4528 6128 4580 6180
rect 10600 6128 10652 6180
rect 11060 6128 11112 6180
rect 15844 6196 15896 6248
rect 14464 6171 14516 6180
rect 1768 6060 1820 6112
rect 3608 6103 3660 6112
rect 3608 6069 3617 6103
rect 3617 6069 3651 6103
rect 3651 6069 3660 6103
rect 3608 6060 3660 6069
rect 5080 6060 5132 6112
rect 5356 6060 5408 6112
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6920 6060 6972 6112
rect 7380 6060 7432 6112
rect 10048 6060 10100 6112
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 10508 6060 10560 6112
rect 10876 6060 10928 6112
rect 11520 6060 11572 6112
rect 11888 6060 11940 6112
rect 12624 6060 12676 6112
rect 13176 6060 13228 6112
rect 13820 6060 13872 6112
rect 14188 6060 14240 6112
rect 14464 6137 14498 6171
rect 14498 6137 14516 6171
rect 14464 6128 14516 6137
rect 15292 6060 15344 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 16212 6103 16264 6112
rect 16212 6069 16221 6103
rect 16221 6069 16255 6103
rect 16255 6069 16264 6103
rect 16212 6060 16264 6069
rect 16304 6103 16356 6112
rect 16304 6069 16313 6103
rect 16313 6069 16347 6103
rect 16347 6069 16356 6103
rect 16304 6060 16356 6069
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1952 5856 2004 5908
rect 3608 5856 3660 5908
rect 6276 5856 6328 5908
rect 6828 5856 6880 5908
rect 9864 5856 9916 5908
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 11888 5856 11940 5908
rect 11980 5856 12032 5908
rect 7472 5788 7524 5840
rect 9312 5788 9364 5840
rect 10324 5788 10376 5840
rect 2688 5720 2740 5772
rect 2780 5720 2832 5772
rect 4712 5720 4764 5772
rect 5356 5720 5408 5772
rect 6828 5720 6880 5772
rect 2136 5695 2188 5704
rect 2136 5661 2145 5695
rect 2145 5661 2179 5695
rect 2179 5661 2188 5695
rect 2136 5652 2188 5661
rect 3148 5652 3200 5704
rect 3976 5652 4028 5704
rect 9220 5720 9272 5772
rect 11796 5763 11848 5772
rect 11796 5729 11830 5763
rect 11830 5729 11848 5763
rect 11796 5720 11848 5729
rect 13268 5788 13320 5840
rect 15568 5831 15620 5840
rect 13544 5763 13596 5772
rect 3332 5584 3384 5636
rect 5080 5516 5132 5568
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 13820 5763 13872 5772
rect 13820 5729 13854 5763
rect 13854 5729 13872 5763
rect 13820 5720 13872 5729
rect 15568 5797 15602 5831
rect 15602 5797 15620 5831
rect 15568 5788 15620 5797
rect 15844 5856 15896 5908
rect 17316 5831 17368 5840
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 10876 5584 10928 5636
rect 11428 5584 11480 5636
rect 13452 5652 13504 5704
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 17960 5720 18012 5772
rect 19800 5652 19852 5704
rect 12900 5627 12952 5636
rect 12900 5593 12909 5627
rect 12909 5593 12943 5627
rect 12943 5593 12952 5627
rect 12900 5584 12952 5593
rect 6552 5516 6604 5568
rect 6736 5516 6788 5568
rect 8024 5516 8076 5568
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 13268 5516 13320 5568
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 15292 5516 15344 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 4068 5312 4120 5364
rect 4804 5312 4856 5364
rect 5540 5312 5592 5364
rect 7472 5312 7524 5364
rect 5724 5244 5776 5296
rect 6184 5244 6236 5296
rect 8300 5312 8352 5364
rect 11060 5312 11112 5364
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 8024 5176 8076 5228
rect 1768 5108 1820 5160
rect 2596 5108 2648 5160
rect 4160 5108 4212 5160
rect 4712 5108 4764 5160
rect 3976 5040 4028 5092
rect 6460 5108 6512 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 8760 5108 8812 5160
rect 10232 5176 10284 5228
rect 14188 5312 14240 5364
rect 16212 5312 16264 5364
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 14464 5176 14516 5228
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 9680 5108 9732 5160
rect 5540 5040 5592 5092
rect 6368 5040 6420 5092
rect 3240 4972 3292 5024
rect 7380 4972 7432 5024
rect 14556 5108 14608 5160
rect 14832 5151 14884 5160
rect 14832 5117 14841 5151
rect 14841 5117 14875 5151
rect 14875 5117 14884 5151
rect 15568 5176 15620 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 14832 5108 14884 5117
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 15936 5040 15988 5092
rect 10140 4972 10192 5024
rect 10416 4972 10468 5024
rect 11060 4972 11112 5024
rect 12900 4972 12952 5024
rect 13636 4972 13688 5024
rect 14188 4972 14240 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 20628 4972 20680 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4712 4768 4764 4820
rect 5632 4768 5684 4820
rect 6092 4768 6144 4820
rect 10692 4768 10744 4820
rect 11704 4768 11756 4820
rect 11980 4768 12032 4820
rect 12900 4811 12952 4820
rect 12900 4777 12909 4811
rect 12909 4777 12943 4811
rect 12943 4777 12952 4811
rect 12900 4768 12952 4777
rect 14188 4811 14240 4820
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 16304 4768 16356 4820
rect 7748 4743 7800 4752
rect 7748 4709 7757 4743
rect 7757 4709 7791 4743
rect 7791 4709 7800 4743
rect 7748 4700 7800 4709
rect 7932 4700 7984 4752
rect 13912 4700 13964 4752
rect 14004 4700 14056 4752
rect 15108 4700 15160 4752
rect 15384 4700 15436 4752
rect 2228 4675 2280 4684
rect 2228 4641 2237 4675
rect 2237 4641 2271 4675
rect 2271 4641 2280 4675
rect 2228 4632 2280 4641
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 4068 4632 4120 4684
rect 4804 4632 4856 4684
rect 4988 4632 5040 4684
rect 6276 4632 6328 4684
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 5448 4564 5500 4616
rect 7380 4632 7432 4684
rect 7104 4564 7156 4616
rect 8208 4564 8260 4616
rect 8852 4675 8904 4684
rect 8852 4641 8861 4675
rect 8861 4641 8895 4675
rect 8895 4641 8904 4675
rect 8852 4632 8904 4641
rect 9312 4632 9364 4684
rect 11796 4632 11848 4684
rect 12072 4632 12124 4684
rect 13268 4675 13320 4684
rect 5540 4539 5592 4548
rect 5540 4505 5549 4539
rect 5549 4505 5583 4539
rect 5583 4505 5592 4539
rect 5540 4496 5592 4505
rect 7656 4496 7708 4548
rect 7932 4496 7984 4548
rect 10232 4607 10284 4616
rect 8392 4539 8444 4548
rect 8392 4505 8401 4539
rect 8401 4505 8435 4539
rect 8435 4505 8444 4539
rect 8392 4496 8444 4505
rect 5080 4428 5132 4480
rect 6184 4428 6236 4480
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 10324 4564 10376 4616
rect 10876 4564 10928 4616
rect 11152 4428 11204 4480
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 12440 4496 12492 4548
rect 14280 4564 14332 4616
rect 15200 4632 15252 4684
rect 15752 4675 15804 4684
rect 15752 4641 15761 4675
rect 15761 4641 15795 4675
rect 15795 4641 15804 4675
rect 15752 4632 15804 4641
rect 16948 4564 17000 4616
rect 17040 4496 17092 4548
rect 13544 4428 13596 4480
rect 18788 4428 18840 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2412 4224 2464 4276
rect 6368 4224 6420 4276
rect 7104 4267 7156 4276
rect 7104 4233 7113 4267
rect 7113 4233 7147 4267
rect 7147 4233 7156 4267
rect 7104 4224 7156 4233
rect 7748 4224 7800 4276
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 6460 4156 6512 4208
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 7288 4088 7340 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 4804 4020 4856 4072
rect 6736 4020 6788 4072
rect 11060 4156 11112 4208
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 10508 4088 10560 4140
rect 11244 4088 11296 4140
rect 11796 4156 11848 4208
rect 13544 4224 13596 4276
rect 13452 4156 13504 4208
rect 9496 4020 9548 4072
rect 10324 4020 10376 4072
rect 11704 4020 11756 4072
rect 12072 4020 12124 4072
rect 14464 4063 14516 4072
rect 3240 3952 3292 4004
rect 3884 3952 3936 4004
rect 4252 3952 4304 4004
rect 10140 3952 10192 4004
rect 10600 3952 10652 4004
rect 3976 3884 4028 3936
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 5264 3884 5316 3936
rect 5540 3884 5592 3936
rect 7104 3884 7156 3936
rect 7748 3884 7800 3936
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 11336 3927 11388 3936
rect 8576 3884 8628 3893
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 11612 3884 11664 3936
rect 11796 3884 11848 3936
rect 12808 3952 12860 4004
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 15936 4088 15988 4140
rect 14648 3952 14700 4004
rect 15016 3952 15068 4004
rect 13176 3884 13228 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3516 3680 3568 3732
rect 2412 3612 2464 3664
rect 4804 3612 4856 3664
rect 5172 3680 5224 3732
rect 7104 3680 7156 3732
rect 10416 3680 10468 3732
rect 11060 3680 11112 3732
rect 8576 3612 8628 3664
rect 9680 3612 9732 3664
rect 10232 3612 10284 3664
rect 13360 3680 13412 3732
rect 11612 3612 11664 3664
rect 11796 3612 11848 3664
rect 16764 3680 16816 3732
rect 13820 3612 13872 3664
rect 6828 3544 6880 3596
rect 7288 3587 7340 3596
rect 7288 3553 7322 3587
rect 7322 3553 7340 3587
rect 7288 3544 7340 3553
rect 7564 3544 7616 3596
rect 1768 3519 1820 3528
rect 1768 3485 1777 3519
rect 1777 3485 1811 3519
rect 1811 3485 1820 3519
rect 1768 3476 1820 3485
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 5172 3476 5224 3528
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 8944 3476 8996 3528
rect 11244 3544 11296 3596
rect 12072 3544 12124 3596
rect 12256 3544 12308 3596
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 11428 3519 11480 3528
rect 9772 3476 9824 3485
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 12532 3544 12584 3596
rect 13912 3544 13964 3596
rect 12900 3476 12952 3528
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 6644 3408 6696 3460
rect 8208 3408 8260 3460
rect 12808 3451 12860 3460
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 14004 3476 14056 3528
rect 15384 3544 15436 3596
rect 16120 3476 16172 3528
rect 12808 3408 12860 3417
rect 3976 3340 4028 3392
rect 5264 3340 5316 3392
rect 5632 3340 5684 3392
rect 6552 3340 6604 3392
rect 8300 3340 8352 3392
rect 10508 3340 10560 3392
rect 11796 3340 11848 3392
rect 12532 3340 12584 3392
rect 12624 3340 12676 3392
rect 14096 3340 14148 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 3332 3136 3384 3188
rect 4160 3136 4212 3188
rect 4804 3136 4856 3188
rect 5356 3136 5408 3188
rect 8392 3136 8444 3188
rect 9312 3136 9364 3188
rect 10232 3136 10284 3188
rect 21088 3136 21140 3188
rect 7288 3068 7340 3120
rect 2872 3000 2924 3052
rect 3240 3000 3292 3052
rect 3976 3000 4028 3052
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 3056 2932 3108 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7104 3000 7156 3052
rect 11060 3068 11112 3120
rect 9220 3000 9272 3052
rect 9864 3000 9916 3052
rect 10508 3000 10560 3052
rect 12716 3068 12768 3120
rect 14280 3068 14332 3120
rect 16028 3068 16080 3120
rect 19248 3068 19300 3120
rect 8208 2975 8260 2984
rect 4252 2864 4304 2916
rect 4712 2864 4764 2916
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 3608 2796 3660 2848
rect 5816 2864 5868 2916
rect 7564 2864 7616 2916
rect 8208 2941 8217 2975
rect 8217 2941 8251 2975
rect 8251 2941 8260 2975
rect 8208 2932 8260 2941
rect 10784 2932 10836 2984
rect 11060 2932 11112 2984
rect 13360 3000 13412 3052
rect 15384 3000 15436 3052
rect 8300 2864 8352 2916
rect 7288 2796 7340 2848
rect 8208 2796 8260 2848
rect 8760 2796 8812 2848
rect 13912 2932 13964 2984
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 15108 2932 15160 2984
rect 22468 3000 22520 3052
rect 16120 2975 16172 2984
rect 15200 2864 15252 2916
rect 10324 2839 10376 2848
rect 10324 2805 10333 2839
rect 10333 2805 10367 2839
rect 10367 2805 10376 2839
rect 10324 2796 10376 2805
rect 10416 2796 10468 2848
rect 11244 2839 11296 2848
rect 11244 2805 11253 2839
rect 11253 2805 11287 2839
rect 11287 2805 11296 2839
rect 11244 2796 11296 2805
rect 12900 2839 12952 2848
rect 12900 2805 12909 2839
rect 12909 2805 12943 2839
rect 12943 2805 12952 2839
rect 12900 2796 12952 2805
rect 13268 2796 13320 2848
rect 16120 2941 16129 2975
rect 16129 2941 16163 2975
rect 16163 2941 16172 2975
rect 16120 2932 16172 2941
rect 17040 2975 17092 2984
rect 17040 2941 17049 2975
rect 17049 2941 17083 2975
rect 17083 2941 17092 2975
rect 17040 2932 17092 2941
rect 17132 2932 17184 2984
rect 18880 2975 18932 2984
rect 18880 2941 18889 2975
rect 18889 2941 18923 2975
rect 18923 2941 18932 2975
rect 18880 2932 18932 2941
rect 22008 2864 22060 2916
rect 16948 2796 17000 2848
rect 17868 2796 17920 2848
rect 19708 2796 19760 2848
rect 19800 2796 19852 2848
rect 21548 2796 21600 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 3424 2592 3476 2644
rect 4068 2635 4120 2644
rect 4068 2601 4077 2635
rect 4077 2601 4111 2635
rect 4111 2601 4120 2635
rect 4068 2592 4120 2601
rect 7380 2592 7432 2644
rect 7564 2635 7616 2644
rect 7564 2601 7573 2635
rect 7573 2601 7607 2635
rect 7607 2601 7616 2635
rect 7564 2592 7616 2601
rect 8392 2592 8444 2644
rect 10416 2592 10468 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 2964 2524 3016 2576
rect 3976 2524 4028 2576
rect 3792 2456 3844 2508
rect 4160 2456 4212 2508
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 2872 2388 2924 2397
rect 5264 2456 5316 2508
rect 6000 2524 6052 2576
rect 8116 2524 8168 2576
rect 9588 2524 9640 2576
rect 10784 2524 10836 2576
rect 19800 2592 19852 2644
rect 5908 2456 5960 2508
rect 20168 2524 20220 2576
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6368 2388 6420 2440
rect 7012 2388 7064 2440
rect 7564 2388 7616 2440
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 6184 2320 6236 2372
rect 8944 2388 8996 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 9864 2388 9916 2440
rect 11060 2320 11112 2372
rect 11612 2388 11664 2440
rect 11704 2388 11756 2440
rect 12900 2320 12952 2372
rect 4068 2252 4120 2304
rect 6092 2252 6144 2304
rect 11152 2252 11204 2304
rect 13084 2456 13136 2508
rect 14004 2499 14056 2508
rect 14004 2465 14013 2499
rect 14013 2465 14047 2499
rect 14047 2465 14056 2499
rect 14004 2456 14056 2465
rect 14188 2456 14240 2508
rect 14832 2456 14884 2508
rect 15292 2456 15344 2508
rect 13544 2388 13596 2440
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 17500 2499 17552 2508
rect 16580 2456 16632 2465
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 15016 2320 15068 2372
rect 14832 2252 14884 2304
rect 15568 2252 15620 2304
rect 16488 2252 16540 2304
rect 17408 2252 17460 2304
rect 17960 2252 18012 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 1124 2048 1176 2100
rect 6460 2048 6512 2100
rect 7288 2048 7340 2100
rect 204 1980 256 2032
rect 5448 1980 5500 2032
rect 5816 1980 5868 2032
rect 13544 2048 13596 2100
rect 11336 1980 11388 2032
rect 12164 1980 12216 2032
rect 664 1912 716 1964
rect 7104 1912 7156 1964
rect 2044 1844 2096 1896
rect 5908 1844 5960 1896
rect 3332 1776 3384 1828
rect 8852 1776 8904 1828
rect 2504 1708 2556 1760
rect 7748 1708 7800 1760
rect 1584 1640 1636 1692
rect 8024 1640 8076 1692
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 1030 22320 1086 22800
rect 1490 22320 1546 22800
rect 1950 22320 2006 22800
rect 2410 22320 2466 22800
rect 2870 22320 2926 22800
rect 3238 22536 3294 22545
rect 3238 22471 3294 22480
rect 216 18426 244 22320
rect 204 18420 256 18426
rect 204 18362 256 18368
rect 584 16454 612 22320
rect 572 16448 624 16454
rect 572 16390 624 16396
rect 1044 16182 1072 22320
rect 1504 19394 1532 22320
rect 1860 19712 1912 19718
rect 1858 19680 1860 19689
rect 1912 19680 1914 19689
rect 1858 19615 1914 19624
rect 1504 19366 1900 19394
rect 1766 19272 1822 19281
rect 1766 19207 1822 19216
rect 1780 19174 1808 19207
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17678 1440 18770
rect 1582 18728 1638 18737
rect 1582 18663 1584 18672
rect 1636 18663 1638 18672
rect 1584 18634 1636 18640
rect 1676 18352 1728 18358
rect 1674 18320 1676 18329
rect 1728 18320 1730 18329
rect 1674 18255 1730 18264
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1766 17368 1822 17377
rect 1766 17303 1768 17312
rect 1820 17303 1822 17312
rect 1768 17274 1820 17280
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1596 16726 1624 17070
rect 1676 16992 1728 16998
rect 1872 16946 1900 19366
rect 1676 16934 1728 16940
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1688 16658 1716 16934
rect 1780 16918 1900 16946
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1582 16416 1638 16425
rect 1582 16351 1638 16360
rect 1596 16250 1624 16351
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1032 16176 1084 16182
rect 1032 16118 1084 16124
rect 1398 16144 1454 16153
rect 1398 16079 1454 16088
rect 1412 16046 1440 16079
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1780 15978 1808 16918
rect 1858 16824 1914 16833
rect 1858 16759 1860 16768
rect 1912 16759 1914 16768
rect 1860 16730 1912 16736
rect 1964 16017 1992 22320
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2240 18154 2268 19178
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 18358 2360 18770
rect 2320 18352 2372 18358
rect 2424 18329 2452 22320
rect 2884 20040 2912 22320
rect 2884 20012 3004 20040
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2320 18294 2372 18300
rect 2410 18320 2466 18329
rect 2410 18255 2466 18264
rect 2228 18148 2280 18154
rect 2228 18090 2280 18096
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 16794 2268 17682
rect 2608 17542 2636 18362
rect 2700 18290 2728 19246
rect 2792 18426 2820 19450
rect 2884 18970 2912 19858
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2700 17270 2728 18226
rect 2976 17864 3004 20012
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 3068 18698 3096 19858
rect 3056 18692 3108 18698
rect 3056 18634 3108 18640
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 2884 17836 3004 17864
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 1950 16008 2006 16017
rect 1768 15972 1820 15978
rect 2884 15978 2912 17836
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2976 17202 3004 17682
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2976 16046 3004 16458
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 1950 15943 2006 15952
rect 2872 15972 2924 15978
rect 1768 15914 1820 15920
rect 2872 15914 2924 15920
rect 1952 15904 2004 15910
rect 1582 15872 1638 15881
rect 2884 15881 2912 15914
rect 1952 15846 2004 15852
rect 2870 15872 2926 15881
rect 1582 15807 1638 15816
rect 1596 15706 1624 15807
rect 1964 15706 1992 15846
rect 2870 15807 2926 15816
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2410 15600 2466 15609
rect 1676 15564 1728 15570
rect 2410 15535 2412 15544
rect 1676 15506 1728 15512
rect 2464 15535 2466 15544
rect 2412 15506 2464 15512
rect 1688 15026 1716 15506
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1674 14920 1730 14929
rect 1674 14855 1730 14864
rect 1688 14618 1716 14855
rect 1676 14612 1728 14618
rect 1676 14554 1728 14560
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 10713 1440 13806
rect 1504 13462 1532 14418
rect 1780 14074 1808 14962
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 14074 2084 14350
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2148 13938 2176 14418
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 2148 13326 2176 13874
rect 2700 13530 2728 14758
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1596 11694 1624 12582
rect 2148 12442 2176 12582
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 1872 11762 1900 12106
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 2056 11218 2084 11630
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1398 10704 1454 10713
rect 1398 10639 1454 10648
rect 1412 7342 1440 10639
rect 2056 10606 2084 11154
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2056 10062 2084 10542
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2056 8974 2084 9998
rect 2332 9466 2360 13330
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2424 11354 2452 12786
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 12306 2820 12582
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11898 2544 12174
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2424 10538 2452 11290
rect 2516 11286 2544 11834
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2412 10532 2464 10538
rect 2412 10474 2464 10480
rect 2884 10282 2912 13330
rect 2976 12481 3004 15982
rect 3068 15745 3096 18294
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3160 17785 3188 17818
rect 3146 17776 3202 17785
rect 3146 17711 3202 17720
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3054 15736 3110 15745
rect 3054 15671 3110 15680
rect 3160 15502 3188 17478
rect 3252 16046 3280 22471
rect 3330 22320 3386 22800
rect 3790 22320 3846 22800
rect 4250 22320 4306 22800
rect 4710 22320 4766 22800
rect 5170 22320 5226 22800
rect 5630 22320 5686 22800
rect 6090 22320 6146 22800
rect 6550 22320 6606 22800
rect 7010 22320 7066 22800
rect 7470 22320 7526 22800
rect 7930 22320 7986 22800
rect 8390 22320 8446 22800
rect 8850 22320 8906 22800
rect 9310 22320 9366 22800
rect 9770 22320 9826 22800
rect 10230 22320 10286 22800
rect 10690 22320 10746 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12438 22320 12494 22800
rect 12898 22320 12954 22800
rect 13358 22320 13414 22800
rect 13818 22320 13874 22800
rect 14278 22320 14334 22800
rect 14738 22320 14794 22800
rect 15198 22320 15254 22800
rect 15658 22320 15714 22800
rect 16118 22320 16174 22800
rect 16578 22320 16634 22800
rect 17038 22320 17094 22800
rect 17498 22320 17554 22800
rect 17958 22320 18014 22800
rect 18418 22320 18474 22800
rect 18878 22320 18934 22800
rect 19338 22320 19394 22800
rect 19798 22320 19854 22800
rect 20258 22320 20314 22800
rect 20718 22320 20774 22800
rect 21178 22320 21234 22800
rect 21638 22320 21694 22800
rect 22098 22320 22154 22800
rect 22558 22320 22614 22800
rect 3344 19394 3372 22320
rect 3514 21584 3570 21593
rect 3514 21519 3570 21528
rect 3344 19366 3464 19394
rect 3436 19281 3464 19366
rect 3422 19272 3478 19281
rect 3332 19236 3384 19242
rect 3422 19207 3478 19216
rect 3332 19178 3384 19184
rect 3344 18970 3372 19178
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3332 18080 3384 18086
rect 3330 18048 3332 18057
rect 3384 18048 3386 18057
rect 3330 17983 3386 17992
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3344 16794 3372 17614
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3436 16658 3464 19110
rect 3528 17882 3556 21519
rect 3698 21176 3754 21185
rect 3698 21111 3754 21120
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3620 18766 3648 19110
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3620 17066 3648 18702
rect 3712 17610 3740 21111
rect 3804 18834 3832 22320
rect 3974 22128 4030 22137
rect 3974 22063 4030 22072
rect 3882 20632 3938 20641
rect 3882 20567 3884 20576
rect 3936 20567 3938 20576
rect 3884 20538 3936 20544
rect 3988 20482 4016 22063
rect 3896 20454 4016 20482
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3790 18728 3846 18737
rect 3790 18663 3846 18672
rect 3700 17604 3752 17610
rect 3700 17546 3752 17552
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3608 16584 3660 16590
rect 3606 16552 3608 16561
rect 3660 16552 3662 16561
rect 3804 16522 3832 18663
rect 3896 17105 3924 20454
rect 3974 20224 4030 20233
rect 3974 20159 4030 20168
rect 3988 19514 4016 20159
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4080 18970 4108 19654
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4172 18714 4200 19994
rect 3988 18686 4200 18714
rect 3882 17096 3938 17105
rect 3882 17031 3938 17040
rect 3606 16487 3662 16496
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3436 15978 3464 16118
rect 3700 16108 3752 16114
rect 3988 16096 4016 18686
rect 4160 18624 4212 18630
rect 4066 18592 4122 18601
rect 4160 18566 4212 18572
rect 4066 18527 4122 18536
rect 4080 18222 4108 18527
rect 4172 18222 4200 18566
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 16522 4108 17546
rect 4172 17066 4200 17682
rect 4264 17134 4292 22320
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4448 20058 4476 20198
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 4724 19938 4752 22320
rect 5184 20058 5212 22320
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 4724 19910 4844 19938
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4724 19310 4752 19790
rect 4712 19304 4764 19310
rect 4342 19272 4398 19281
rect 4712 19246 4764 19252
rect 4342 19207 4398 19216
rect 4356 18766 4384 19207
rect 4618 18864 4674 18873
rect 4618 18799 4674 18808
rect 4632 18766 4660 18799
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4724 18426 4752 19246
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 17338 4752 17682
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4172 16658 4200 17002
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 3700 16050 3752 16056
rect 3896 16068 4016 16096
rect 3424 15972 3476 15978
rect 3424 15914 3476 15920
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3514 15736 3570 15745
rect 3514 15671 3570 15680
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3422 15464 3478 15473
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3068 14346 3096 14962
rect 3160 14822 3188 15438
rect 3422 15399 3478 15408
rect 3436 15162 3464 15399
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3068 13870 3096 14282
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 12918 3188 13670
rect 3148 12912 3200 12918
rect 3148 12854 3200 12860
rect 2962 12472 3018 12481
rect 2962 12407 3018 12416
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2792 10254 2912 10282
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2332 9438 2452 9466
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 1596 8090 1624 8910
rect 2056 8634 2084 8910
rect 2332 8634 2360 9318
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 2424 7342 2452 9438
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2516 7886 2544 9046
rect 2608 8566 2636 9522
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 1400 7336 1452 7342
rect 2412 7336 2464 7342
rect 1400 7278 1452 7284
rect 2410 7304 2412 7313
rect 2464 7304 2466 7313
rect 2410 7239 2466 7248
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6118 1808 6802
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5166 1808 6054
rect 1964 5914 1992 7142
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 2148 6440 2176 6870
rect 2228 6452 2280 6458
rect 2148 6412 2228 6440
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2148 5710 2176 6412
rect 2228 6394 2280 6400
rect 2516 6186 2544 7346
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2608 5166 2636 8502
rect 2700 6934 2728 9454
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 2700 5778 2728 6734
rect 2792 5778 2820 10254
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2884 7410 2912 10066
rect 3068 9654 3096 11154
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 6730 2912 7346
rect 2976 7002 3004 7686
rect 3160 7290 3188 12378
rect 3252 10266 3280 14894
rect 3330 14512 3386 14521
rect 3330 14447 3386 14456
rect 3344 13530 3372 14447
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3436 13462 3464 13738
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3528 13308 3556 15671
rect 3620 13938 3648 15846
rect 3712 15502 3740 16050
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 15065 3740 15438
rect 3698 15056 3754 15065
rect 3698 14991 3754 15000
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14074 3740 14894
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3344 13280 3556 13308
rect 3344 12442 3372 13280
rect 3712 13258 3740 14010
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3068 7262 3188 7290
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 1780 4078 1808 5102
rect 2228 4684 2280 4690
rect 2228 4626 2280 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1780 3534 1808 4014
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2240 2650 2268 4626
rect 2332 3194 2360 4626
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2424 4282 2452 4558
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2424 3670 2452 4218
rect 2792 4049 2820 5714
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2976 3097 3004 6802
rect 2962 3088 3018 3097
rect 2872 3052 2924 3058
rect 2962 3023 3018 3032
rect 2872 2994 2924 3000
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1124 2100 1176 2106
rect 1124 2042 1176 2048
rect 204 2032 256 2038
rect 204 1974 256 1980
rect 216 480 244 1974
rect 664 1964 716 1970
rect 664 1906 716 1912
rect 676 480 704 1906
rect 1136 480 1164 2042
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 1584 1692 1636 1698
rect 1584 1634 1636 1640
rect 1596 480 1624 1634
rect 2056 480 2084 1838
rect 2504 1760 2556 1766
rect 2504 1702 2556 1708
rect 2516 480 2544 1702
rect 2792 1193 2820 2790
rect 2884 2446 2912 2994
rect 2976 2582 3004 3023
rect 3068 2990 3096 7262
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 5817 3188 7142
rect 3146 5808 3202 5817
rect 3146 5743 3202 5752
rect 3148 5704 3200 5710
rect 3252 5692 3280 7482
rect 3344 7290 3372 12242
rect 3436 9518 3464 12922
rect 3620 12617 3648 13126
rect 3712 12986 3740 13194
rect 3804 13025 3832 13738
rect 3896 13734 3924 16068
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3988 15026 4016 15914
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15706 4108 15846
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4172 15366 4200 16390
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3974 13968 4030 13977
rect 4080 13938 4108 14214
rect 3974 13903 4030 13912
rect 4068 13932 4120 13938
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3790 13016 3846 13025
rect 3700 12980 3752 12986
rect 3790 12951 3846 12960
rect 3700 12922 3752 12928
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 3712 12238 3740 12786
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3712 11694 3740 12174
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3712 10266 3740 11630
rect 3804 11286 3832 12718
rect 3792 11280 3844 11286
rect 3792 11222 3844 11228
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3424 8832 3476 8838
rect 3528 8820 3556 9522
rect 3790 9344 3846 9353
rect 3790 9279 3846 9288
rect 3476 8792 3556 8820
rect 3424 8774 3476 8780
rect 3436 8498 3464 8774
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7818 3464 8230
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3344 7262 3556 7290
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3200 5664 3280 5692
rect 3148 5646 3200 5652
rect 3160 3913 3188 5646
rect 3344 5642 3372 7142
rect 3436 6458 3464 7142
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3252 4010 3280 4966
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3146 3904 3202 3913
rect 3146 3839 3202 3848
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3068 2145 3096 2926
rect 3054 2136 3110 2145
rect 3054 2071 3110 2080
rect 3160 2020 3188 3839
rect 3252 3058 3280 3946
rect 3344 3194 3372 4558
rect 3528 3890 3556 7262
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 5914 3648 6054
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3528 3862 3648 3890
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3436 2650 3464 3470
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 2976 1992 3188 2020
rect 2778 1184 2834 1193
rect 2778 1119 2834 1128
rect 2976 480 3004 1992
rect 3332 1828 3384 1834
rect 3332 1770 3384 1776
rect 3344 1601 3372 1770
rect 3330 1592 3386 1601
rect 3330 1527 3386 1536
rect 3528 1442 3556 3674
rect 3620 2854 3648 3862
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3804 2514 3832 9279
rect 3896 5234 3924 13330
rect 3988 12986 4016 13903
rect 4068 13874 4120 13880
rect 4172 13870 4200 14826
rect 4264 14550 4292 16118
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4526 16008 4582 16017
rect 4526 15943 4582 15952
rect 4434 15872 4490 15881
rect 4434 15807 4490 15816
rect 4448 15570 4476 15807
rect 4540 15706 4568 15943
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4540 15473 4568 15642
rect 4526 15464 4582 15473
rect 4526 15399 4582 15408
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4724 14482 4752 16050
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4816 14385 4844 19910
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5000 19310 5028 19790
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5000 18834 5028 19246
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4908 18714 4936 18770
rect 5276 18714 5304 19858
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 4908 18686 5028 18714
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4908 18086 4936 18566
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16794 4936 16934
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4896 15904 4948 15910
rect 4894 15872 4896 15881
rect 4948 15872 4950 15881
rect 4894 15807 4950 15816
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4908 14890 4936 15438
rect 4896 14884 4948 14890
rect 4896 14826 4948 14832
rect 4250 14376 4306 14385
rect 4250 14311 4306 14320
rect 4802 14376 4858 14385
rect 4802 14311 4858 14320
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4066 13560 4122 13569
rect 4122 13518 4200 13546
rect 4066 13495 4122 13504
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3974 12336 4030 12345
rect 3974 12271 3976 12280
rect 4028 12271 4030 12280
rect 3976 12242 4028 12248
rect 4080 11354 4108 13398
rect 4172 12374 4200 13518
rect 4264 12753 4292 14311
rect 4712 14272 4764 14278
rect 5000 14260 5028 18686
rect 5080 18692 5132 18698
rect 5080 18634 5132 18640
rect 5184 18686 5304 18714
rect 5092 18426 5120 18634
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5080 18080 5132 18086
rect 5078 18048 5080 18057
rect 5132 18048 5134 18057
rect 5078 17983 5134 17992
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 5092 15706 5120 16662
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 4712 14214 4764 14220
rect 4816 14232 5028 14260
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4356 13462 4384 13942
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4250 12744 4306 12753
rect 4250 12679 4306 12688
rect 4264 12442 4292 12679
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4250 11656 4306 11665
rect 4250 11591 4306 11600
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4264 10033 4292 11591
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4356 11082 4384 11494
rect 4448 11354 4476 11494
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4724 11234 4752 14214
rect 4816 12442 4844 14232
rect 4894 14104 4950 14113
rect 4894 14039 4896 14048
rect 4948 14039 4950 14048
rect 4896 14010 4948 14016
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4908 11762 4936 12038
rect 5000 11898 5028 12650
rect 5092 11898 5120 15098
rect 5184 14278 5212 18686
rect 5368 16998 5396 19654
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5460 18834 5488 18906
rect 5552 18873 5580 19654
rect 5538 18864 5594 18873
rect 5448 18828 5500 18834
rect 5538 18799 5594 18808
rect 5448 18770 5500 18776
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5264 16992 5316 16998
rect 5262 16960 5264 16969
rect 5356 16992 5408 16998
rect 5316 16960 5318 16969
rect 5356 16934 5408 16940
rect 5262 16895 5318 16904
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5368 15502 5396 16730
rect 5460 16561 5488 17478
rect 5552 17338 5580 17546
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5644 17218 5672 22320
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5736 18970 5764 19178
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5736 18290 5764 18906
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5828 17746 5856 19926
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 6104 17592 6132 22320
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6380 18358 6408 20538
rect 6460 19916 6512 19922
rect 6460 19858 6512 19864
rect 6472 19174 6500 19858
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6472 18358 6500 19110
rect 6368 18352 6420 18358
rect 6368 18294 6420 18300
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 5552 17190 5672 17218
rect 5828 17564 6132 17592
rect 5446 16552 5502 16561
rect 5446 16487 5502 16496
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15706 5488 15846
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5276 14770 5304 15030
rect 5276 14742 5396 14770
rect 5368 14414 5396 14742
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5460 13870 5488 15302
rect 5448 13864 5500 13870
rect 5354 13832 5410 13841
rect 5448 13806 5500 13812
rect 5354 13767 5410 13776
rect 5368 13734 5396 13767
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5460 12102 5488 13806
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4986 11792 5042 11801
rect 4896 11756 4948 11762
rect 4986 11727 5042 11736
rect 4896 11698 4948 11704
rect 4724 11206 4936 11234
rect 4804 11144 4856 11150
rect 4804 11086 4856 11092
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4632 10305 4660 10474
rect 4618 10296 4674 10305
rect 4618 10231 4674 10240
rect 4526 10160 4582 10169
rect 4526 10095 4528 10104
rect 4580 10095 4582 10104
rect 4528 10066 4580 10072
rect 4724 10062 4752 10746
rect 4816 10538 4844 11086
rect 4908 10577 4936 11206
rect 4894 10568 4950 10577
rect 4804 10532 4856 10538
rect 4894 10503 4950 10512
rect 4804 10474 4856 10480
rect 4712 10056 4764 10062
rect 4250 10024 4306 10033
rect 4712 9998 4764 10004
rect 4250 9959 4306 9968
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3974 9752 4030 9761
rect 3974 9687 3976 9696
rect 4028 9687 4030 9696
rect 3976 9658 4028 9664
rect 3974 8800 4030 8809
rect 3974 8735 4030 8744
rect 3988 8634 4016 8735
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4080 8430 4108 9862
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4172 9042 4200 9386
rect 4264 9194 4292 9959
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4620 9580 4672 9586
rect 4724 9568 4752 9998
rect 4672 9540 4752 9568
rect 4620 9522 4672 9528
rect 4264 9166 4384 9194
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4356 8888 4384 9166
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4172 8860 4384 8888
rect 4172 8498 4200 8860
rect 4448 8820 4476 8978
rect 4632 8974 4660 9522
rect 4712 9376 4764 9382
rect 4908 9364 4936 10503
rect 4764 9336 4936 9364
rect 4712 9318 4764 9324
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4264 8792 4476 8820
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4068 8288 4120 8294
rect 3974 8256 4030 8265
rect 4068 8230 4120 8236
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3974 8191 4030 8200
rect 3988 7954 4016 8191
rect 4080 8022 4108 8230
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 4066 7848 4122 7857
rect 4066 7783 4068 7792
rect 4120 7783 4122 7792
rect 4068 7754 4120 7760
rect 4172 7410 4200 8230
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6390 4108 6831
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3988 5710 4016 6258
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3974 5400 4030 5409
rect 3974 5335 4030 5344
rect 4068 5364 4120 5370
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3988 5098 4016 5335
rect 4068 5306 4120 5312
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 4080 5001 4108 5306
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4066 4992 4122 5001
rect 4066 4927 4122 4936
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3436 1414 3556 1442
rect 3436 480 3464 1414
rect 3896 480 3924 3946
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3988 3398 4016 3878
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3988 2582 4016 2994
rect 4080 2650 4108 4626
rect 4172 3194 4200 5102
rect 4264 4010 4292 8792
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8294 4752 9318
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4356 7886 4384 8026
rect 4816 8022 4844 8910
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4724 7342 4752 7686
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4724 6662 4752 7278
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4528 6180 4580 6186
rect 4528 6122 4580 6128
rect 4540 5953 4568 6122
rect 4526 5944 4582 5953
rect 4526 5879 4582 5888
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5166 4752 5714
rect 4816 5370 4844 7958
rect 4908 7886 4936 8434
rect 5000 8090 5028 11727
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5460 11506 5488 11562
rect 5276 11478 5488 11506
rect 5276 11354 5304 11478
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 9042 5120 10474
rect 5172 10056 5224 10062
rect 5170 10024 5172 10033
rect 5224 10024 5226 10033
rect 5276 10010 5304 11290
rect 5276 9982 5488 10010
rect 5170 9959 5226 9968
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5092 8838 5120 8978
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 8498 5120 8774
rect 5080 8492 5132 8498
rect 5184 8480 5212 9386
rect 5276 9042 5304 9454
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5184 8452 5304 8480
rect 5080 8434 5132 8440
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4908 6934 4936 7822
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 5000 6338 5028 8026
rect 5092 7274 5120 8434
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4908 6310 5028 6338
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4712 5160 4764 5166
rect 4764 5120 4844 5148
rect 4712 5102 4764 5108
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4724 2922 4752 4762
rect 4816 4690 4844 5120
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4816 4078 4844 4626
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3670 4844 4014
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4908 3505 4936 6310
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5000 4690 5028 6190
rect 5080 6112 5132 6118
rect 5184 6100 5212 8230
rect 5276 6254 5304 8452
rect 5368 7954 5396 9318
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5460 7834 5488 9982
rect 5552 9178 5580 17190
rect 5722 15872 5778 15881
rect 5722 15807 5778 15816
rect 5736 15162 5764 15807
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5736 13530 5764 13874
rect 5828 13818 5856 17564
rect 6564 17490 6592 22320
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 6932 19310 6960 19926
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6656 18154 6684 19178
rect 6918 18320 6974 18329
rect 7024 18290 7052 22320
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 6918 18255 6974 18264
rect 7012 18284 7064 18290
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6104 17462 6592 17490
rect 5998 17096 6054 17105
rect 5998 17031 6054 17040
rect 6012 16998 6040 17031
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5998 16008 6054 16017
rect 5998 15943 6054 15952
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5920 15745 5948 15846
rect 5906 15736 5962 15745
rect 5906 15671 5962 15680
rect 5906 14920 5962 14929
rect 5906 14855 5962 14864
rect 5920 14550 5948 14855
rect 6012 14550 6040 15943
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 5828 13790 5948 13818
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5736 12782 5764 13466
rect 5828 13394 5856 13670
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5828 12986 5856 13330
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 10130 5672 10406
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5632 9988 5684 9994
rect 5736 9976 5764 12378
rect 5828 12306 5856 12922
rect 5920 12866 5948 13790
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6012 12986 6040 13330
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5920 12838 6040 12866
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5920 11762 5948 12582
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 10742 5856 11154
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5814 10296 5870 10305
rect 5814 10231 5870 10240
rect 5828 10062 5856 10231
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5684 9948 5764 9976
rect 5632 9930 5684 9936
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5552 8090 5580 8298
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5368 7806 5488 7834
rect 5368 6882 5396 7806
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7342 5488 7686
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5368 6854 5488 6882
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5368 6118 5396 6734
rect 5356 6112 5408 6118
rect 5184 6072 5304 6100
rect 5080 6054 5132 6060
rect 5092 5574 5120 6054
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4894 3496 4950 3505
rect 4894 3431 4950 3440
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4712 2916 4764 2922
rect 4712 2858 4764 2864
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 4066 2544 4122 2553
rect 4066 2479 4122 2488
rect 4160 2508 4212 2514
rect 4080 2310 4108 2479
rect 4160 2450 4212 2456
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2502 0 2558 480
rect 2962 0 3018 480
rect 3422 0 3478 480
rect 3882 0 3938 480
rect 4172 241 4200 2450
rect 4264 1442 4292 2858
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1414 4384 1442
rect 4356 480 4384 1414
rect 4816 480 4844 3130
rect 5092 2972 5120 4422
rect 5276 3942 5304 6072
rect 5356 6054 5408 6060
rect 5368 5778 5396 6054
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5460 4706 5488 6854
rect 5552 5370 5580 8026
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5644 5148 5672 9386
rect 5736 5302 5764 9948
rect 5828 9586 5856 9998
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7546 5856 7890
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 6012 7290 6040 12838
rect 5828 7262 6040 7290
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5644 5120 5764 5148
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5368 4678 5488 4706
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5184 3738 5212 3878
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5172 3528 5224 3534
rect 5170 3496 5172 3505
rect 5224 3496 5226 3505
rect 5170 3431 5226 3440
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5276 3058 5304 3334
rect 5368 3194 5396 4678
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5172 2984 5224 2990
rect 5092 2944 5172 2972
rect 5172 2926 5224 2932
rect 5460 2553 5488 4558
rect 5552 4554 5580 5034
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5446 2544 5502 2553
rect 5264 2508 5316 2514
rect 5446 2479 5502 2488
rect 5264 2450 5316 2456
rect 5276 480 5304 2450
rect 5460 2038 5488 2479
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 5552 649 5580 3878
rect 5644 3398 5672 4762
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5538 640 5594 649
rect 5538 575 5594 584
rect 5736 480 5764 5120
rect 5828 2961 5856 7262
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5814 2952 5870 2961
rect 5814 2887 5816 2896
rect 5868 2887 5870 2896
rect 5816 2858 5868 2864
rect 5828 2827 5856 2858
rect 5920 2514 5948 6870
rect 6012 6866 6040 7142
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6104 6746 6132 17462
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6196 16046 6224 17274
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6288 16590 6316 16934
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6288 15706 6316 15914
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6380 15162 6408 17070
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14482 6316 14894
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6288 12850 6316 13942
rect 6380 13870 6408 15098
rect 6656 14498 6684 17818
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6748 15706 6776 17206
rect 6840 16794 6868 17682
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6840 16153 6868 16186
rect 6826 16144 6882 16153
rect 6826 16079 6882 16088
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6840 15502 6868 15846
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6564 14470 6684 14498
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6564 12442 6592 14470
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11354 6224 12242
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6288 10606 6316 10950
rect 6656 10713 6684 14350
rect 6748 13734 6776 14894
rect 6932 13954 6960 18255
rect 7012 18226 7064 18232
rect 7208 18222 7236 19790
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7300 18766 7328 19246
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7208 17882 7236 18022
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7300 17678 7328 18702
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 15706 7144 17478
rect 7208 17066 7236 17614
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7300 16998 7328 17614
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7208 16046 7236 16186
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7300 15434 7328 16934
rect 7392 15502 7420 16934
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7286 15056 7342 15065
rect 7286 14991 7342 15000
rect 7300 14890 7328 14991
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7300 14396 7328 14826
rect 7392 14550 7420 14826
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7300 14368 7420 14396
rect 6932 13926 7052 13954
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6748 13326 6776 13670
rect 6736 13320 6788 13326
rect 6788 13280 6868 13308
rect 6736 13262 6788 13268
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6748 11150 6776 12854
rect 6840 12782 6868 13280
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6932 12442 6960 13806
rect 7024 12714 7052 13926
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 7010 12472 7066 12481
rect 6920 12436 6972 12442
rect 7010 12407 7066 12416
rect 6920 12378 6972 12384
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11218 6960 11494
rect 7024 11354 7052 12407
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6642 10704 6698 10713
rect 6748 10674 6776 11086
rect 6642 10639 6698 10648
rect 6736 10668 6788 10674
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10464 6328 10470
rect 6274 10432 6276 10441
rect 6328 10432 6330 10441
rect 6274 10367 6330 10376
rect 6380 10130 6408 10542
rect 6656 10248 6684 10639
rect 6736 10610 6788 10616
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6472 10220 6684 10248
rect 6472 10130 6500 10220
rect 6932 10130 6960 10406
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6656 8838 6684 10066
rect 7024 9586 7052 11154
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7116 9466 7144 13330
rect 7208 11082 7236 13670
rect 7300 12986 7328 13670
rect 7392 12986 7420 14368
rect 7484 13818 7512 22320
rect 7944 20346 7972 22320
rect 7760 20318 7972 20346
rect 7760 18086 7788 20318
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 8220 19174 8248 19722
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18902 8248 19110
rect 8208 18896 8260 18902
rect 8208 18838 8260 18844
rect 8312 18358 8340 19790
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7564 17876 7616 17882
rect 7564 17818 7616 17824
rect 7576 16969 7604 17818
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7562 16960 7618 16969
rect 7562 16895 7618 16904
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7576 16114 7604 16594
rect 7668 16522 7696 17002
rect 7760 16998 7788 17682
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7760 15706 7788 16390
rect 8220 16250 8248 16390
rect 8312 16250 8340 18090
rect 8404 17354 8432 22320
rect 8864 20040 8892 22320
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8588 20012 8892 20040
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8496 18426 8524 19790
rect 8588 19281 8616 20012
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8574 19272 8630 19281
rect 8574 19207 8630 19216
rect 8772 18970 8800 19858
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8588 17814 8616 18362
rect 8864 18290 8892 18838
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8404 17326 8616 17354
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16726 8524 16934
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8312 15638 8340 15846
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8220 15094 8248 15506
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 14113 7604 14282
rect 7562 14104 7618 14113
rect 7668 14074 7696 14350
rect 7562 14039 7618 14048
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7484 13790 7604 13818
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12481 7420 12582
rect 7378 12472 7434 12481
rect 7378 12407 7434 12416
rect 7286 12200 7342 12209
rect 7286 12135 7342 12144
rect 7300 11558 7328 12135
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7116 9438 7236 9466
rect 7300 9450 7328 11494
rect 7392 10656 7420 12038
rect 7484 10810 7512 13670
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7392 10628 7512 10656
rect 7484 9994 7512 10628
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6748 8922 6776 9114
rect 7116 9110 7144 9318
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6748 8894 6960 8922
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6196 7290 6224 7822
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7478 6316 7686
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6196 7262 6316 7290
rect 6012 6718 6132 6746
rect 6012 2582 6040 6718
rect 6288 6322 6316 7262
rect 6380 6934 6408 7890
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 4826 6132 6054
rect 6288 5914 6316 6258
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6184 5296 6236 5302
rect 6184 5238 6236 5244
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6090 4584 6146 4593
rect 6196 4570 6224 5238
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6146 4542 6224 4570
rect 6090 4519 6146 4528
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5828 2038 5856 2382
rect 5816 2032 5868 2038
rect 5816 1974 5868 1980
rect 5920 1902 5948 2450
rect 6104 2310 6132 4519
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6196 4146 6224 4422
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6196 3754 6224 4082
rect 6288 4060 6316 4626
rect 6380 4282 6408 5034
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6472 4214 6500 5102
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6288 4032 6500 4060
rect 6196 3726 6408 3754
rect 6182 3632 6238 3641
rect 6182 3567 6238 3576
rect 6196 2378 6224 3567
rect 6380 3534 6408 3726
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6380 2446 6408 3470
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6196 480 6224 2314
rect 6472 2106 6500 4032
rect 6564 3398 6592 5510
rect 6656 3466 6684 7890
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 5574 6776 7822
rect 6932 6322 6960 8894
rect 7024 8673 7052 8978
rect 7010 8664 7066 8673
rect 7010 8599 7066 8608
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6932 6225 6960 6258
rect 6918 6216 6974 6225
rect 6918 6151 6974 6160
rect 6920 6112 6972 6118
rect 6840 6072 6920 6100
rect 6840 5914 6868 6072
rect 6920 6054 6972 6060
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6840 5166 6868 5714
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6736 4072 6788 4078
rect 6734 4040 6736 4049
rect 6788 4040 6790 4049
rect 6734 3975 6790 3984
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6748 2836 6776 3975
rect 6840 3602 6868 5102
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6748 2808 6868 2836
rect 6840 2666 6868 2808
rect 6656 2638 6868 2666
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6656 480 6684 2638
rect 7024 2446 7052 8599
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7116 5386 7144 7890
rect 7208 7546 7236 9438
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 9353 7328 9386
rect 7286 9344 7342 9353
rect 7286 9279 7342 9288
rect 7392 8974 7420 9522
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7300 8090 7328 8910
rect 7392 8634 7420 8910
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7484 8514 7512 9930
rect 7392 8486 7512 8514
rect 7392 8362 7420 8486
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7576 7750 7604 13790
rect 7668 13394 7696 13874
rect 7760 13530 7788 14350
rect 7852 14074 7880 14418
rect 8220 14414 8248 14894
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7760 12850 7788 13466
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7668 12238 7696 12786
rect 7944 12730 7972 13330
rect 7760 12702 7972 12730
rect 7760 12646 7788 12702
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7654 11656 7710 11665
rect 7654 11591 7710 11600
rect 7668 11218 7696 11591
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7668 8838 7696 9862
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7668 7954 7696 8026
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7208 6798 7236 7142
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7300 6458 7328 7142
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7392 6338 7420 6598
rect 7300 6310 7420 6338
rect 7472 6316 7524 6322
rect 7116 5358 7236 5386
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 4282 7144 4558
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7104 3936 7156 3942
rect 7102 3904 7104 3913
rect 7156 3904 7158 3913
rect 7102 3839 7158 3848
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7116 3058 7144 3674
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7116 1970 7144 2994
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7208 1442 7236 5358
rect 7300 4146 7328 6310
rect 7472 6258 7524 6264
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 6118 7420 6190
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7484 5846 7512 6258
rect 7472 5840 7524 5846
rect 7392 5800 7472 5828
rect 7392 5030 7420 5800
rect 7472 5782 7524 5788
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4690 7420 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3602 7328 4082
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7300 3126 7328 3538
rect 7288 3120 7340 3126
rect 7286 3088 7288 3097
rect 7340 3088 7342 3097
rect 7286 3023 7342 3032
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7300 2106 7328 2790
rect 7484 2666 7512 5306
rect 7576 3602 7604 6598
rect 7668 4554 7696 7346
rect 7760 7274 7788 12242
rect 8312 11778 8340 14418
rect 8496 14278 8524 14758
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8220 11750 8340 11778
rect 8220 11694 8248 11750
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10266 8248 11494
rect 8298 10704 8354 10713
rect 8298 10639 8354 10648
rect 8312 10470 8340 10639
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9654 8340 9998
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8312 9042 8340 9318
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7944 8430 7972 8774
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8404 8022 8432 14214
rect 8482 12744 8538 12753
rect 8482 12679 8538 12688
rect 8496 12306 8524 12679
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 11286 8524 11562
rect 8588 11286 8616 17326
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8680 14006 8708 14894
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8680 11121 8708 11766
rect 8666 11112 8722 11121
rect 8666 11047 8722 11056
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8574 10160 8630 10169
rect 8574 10095 8630 10104
rect 8482 9480 8538 9489
rect 8482 9415 8538 9424
rect 8496 9382 8524 9415
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7750 7972 7822
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 7449 7972 7686
rect 7930 7440 7986 7449
rect 7930 7375 7986 7384
rect 8312 7290 8340 7958
rect 7748 7268 7800 7274
rect 8312 7262 8432 7290
rect 7748 7210 7800 7216
rect 7760 6390 7788 7210
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 8024 6248 8076 6254
rect 8076 6208 8248 6236
rect 8024 6190 8076 6196
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5234 8064 5510
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7748 4752 7800 4758
rect 7932 4752 7984 4758
rect 7748 4694 7800 4700
rect 7930 4720 7932 4729
rect 7984 4720 7986 4729
rect 8220 4706 8248 6208
rect 8312 5370 8340 7142
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7760 4282 7788 4694
rect 7930 4655 7986 4664
rect 8128 4678 8248 4706
rect 7930 4584 7986 4593
rect 7930 4519 7932 4528
rect 7984 4519 7986 4528
rect 7932 4490 7984 4496
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7748 3936 7800 3942
rect 8128 3924 8156 4678
rect 8208 4616 8260 4622
rect 8260 4576 8340 4604
rect 8208 4558 8260 4564
rect 8128 3896 8248 3924
rect 7748 3878 7800 3884
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7392 2650 7512 2666
rect 7576 2650 7604 2858
rect 7380 2644 7512 2650
rect 7432 2638 7512 2644
rect 7564 2644 7616 2650
rect 7380 2586 7432 2592
rect 7564 2586 7616 2592
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7116 1414 7236 1442
rect 7116 480 7144 1414
rect 7576 480 7604 2382
rect 7760 1766 7788 3878
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8220 3466 8248 3896
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 2990 8248 3402
rect 8312 3398 8340 4576
rect 8404 4554 8432 7262
rect 8496 7188 8524 9318
rect 8588 7256 8616 10095
rect 8680 9926 8708 10542
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8680 9586 8708 9862
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8772 9382 8800 18022
rect 8956 17678 8984 20198
rect 9324 18970 9352 22320
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9404 19236 9456 19242
rect 9404 19178 9456 19184
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9416 18630 9444 19178
rect 9600 18766 9628 19246
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9416 18290 9444 18566
rect 9692 18358 9720 19790
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 9232 16590 9260 18022
rect 9784 17728 9812 22320
rect 10244 19802 10272 22320
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 9692 17700 9812 17728
rect 10152 19774 10272 19802
rect 9692 17626 9720 17700
rect 9600 17598 9720 17626
rect 9772 17604 9824 17610
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 8942 15464 8998 15473
rect 8942 15399 8998 15408
rect 8956 13938 8984 15399
rect 9034 14784 9090 14793
rect 9034 14719 9090 14728
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8850 13832 8906 13841
rect 8850 13767 8906 13776
rect 8864 13530 8892 13767
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8956 12442 8984 12650
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 10810 8892 11494
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8956 10742 8984 11154
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 8968 8720 8974
rect 8666 8936 8668 8945
rect 8720 8936 8722 8945
rect 8666 8871 8722 8880
rect 8772 8401 8800 9318
rect 8758 8392 8814 8401
rect 8758 8327 8814 8336
rect 8588 7228 8800 7256
rect 8496 7160 8708 7188
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6458 8616 6598
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8680 4978 8708 7160
rect 8772 6338 8800 7228
rect 8864 6474 8892 10134
rect 8956 10062 8984 10678
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9048 6610 9076 14719
rect 9140 12374 9168 16390
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9140 10044 9168 11154
rect 9232 10169 9260 16526
rect 9600 16522 9628 17598
rect 9772 17546 9824 17552
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9600 16114 9628 16458
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9324 15706 9352 16050
rect 9692 15978 9720 17478
rect 9784 17134 9812 17546
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9876 17338 9904 17478
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9876 15994 9904 17002
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9968 16046 9996 16730
rect 10060 16114 10088 17206
rect 10152 16810 10180 19774
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10244 18154 10272 19654
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10152 16794 10364 16810
rect 10140 16788 10364 16794
rect 10192 16782 10364 16788
rect 10140 16730 10192 16736
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9784 15966 9904 15994
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10046 16008 10102 16017
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9324 15026 9352 15642
rect 9680 15564 9732 15570
rect 9784 15552 9812 15966
rect 10046 15943 10102 15952
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9732 15524 9812 15552
rect 9680 15506 9732 15512
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9324 14074 9352 14758
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 14074 9444 14350
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9404 13864 9456 13870
rect 9456 13824 9536 13852
rect 9404 13806 9456 13812
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9324 11286 9352 11698
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9324 11082 9352 11222
rect 9416 11218 9444 11698
rect 9508 11558 9536 13824
rect 9600 12442 9628 15030
rect 9784 15026 9812 15524
rect 9876 15162 9904 15846
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9956 15088 10008 15094
rect 9954 15056 9956 15065
rect 10008 15056 10010 15065
rect 9772 15020 9824 15026
rect 9954 14991 10010 15000
rect 9772 14962 9824 14968
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9692 14618 9720 14758
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9784 14482 9812 14758
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9968 13977 9996 14554
rect 9954 13968 10010 13977
rect 9864 13932 9916 13938
rect 9954 13903 10010 13912
rect 9864 13874 9916 13880
rect 9876 13734 9904 13874
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9784 13462 9812 13670
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 12986 9720 13330
rect 10060 13326 10088 15943
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9692 12345 9720 12378
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9586 12064 9642 12073
rect 9586 11999 9642 12008
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9324 10606 9352 10678
rect 9312 10600 9364 10606
rect 9404 10600 9456 10606
rect 9312 10542 9364 10548
rect 9402 10568 9404 10577
rect 9456 10568 9458 10577
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9140 10016 9260 10044
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 8022 9168 8230
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9232 6905 9260 10016
rect 9324 7886 9352 10542
rect 9402 10503 9458 10512
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9416 9926 9444 10066
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9508 9518 9536 11494
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9600 9466 9628 11999
rect 9692 11014 9720 12174
rect 9784 11218 9812 12174
rect 9968 11529 9996 13194
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12782 10088 13126
rect 10152 12866 10180 16458
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10244 14958 10272 15982
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10244 14414 10272 14894
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 13938 10272 14350
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10244 12986 10272 13262
rect 10336 13002 10364 16782
rect 10428 15638 10456 18906
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10520 16590 10548 17614
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10428 13938 10456 14214
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10612 13530 10640 19858
rect 10704 18222 10732 22320
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10980 19242 11008 19790
rect 11072 19378 11100 19858
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10888 18902 10916 19110
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 11072 18834 11100 19110
rect 11164 18834 11192 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11256 18714 11284 19314
rect 11624 18902 11652 22320
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 11072 18686 11284 18714
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 16833 10824 18022
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10980 17338 11008 17682
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10782 16824 10838 16833
rect 10980 16810 11008 16934
rect 10888 16794 11008 16810
rect 10782 16759 10838 16768
rect 10876 16788 11008 16794
rect 10928 16782 11008 16788
rect 10876 16730 10928 16736
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10704 15706 10732 16050
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10704 14890 10732 15642
rect 10796 15366 10824 15846
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10968 14544 11020 14550
rect 10966 14512 10968 14521
rect 11020 14512 11022 14521
rect 10876 14476 10928 14482
rect 10966 14447 11022 14456
rect 10876 14418 10928 14424
rect 10888 14006 10916 14418
rect 11072 14414 11100 18686
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 17218 11192 18566
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11716 18358 11744 19110
rect 11900 18834 11928 19246
rect 11992 18970 12020 22320
rect 12452 20058 12480 22320
rect 12912 20058 12940 22320
rect 13372 20058 13400 22320
rect 13832 20074 13860 22320
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13360 20052 13412 20058
rect 13832 20046 13952 20074
rect 13360 19994 13412 20000
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17921 11560 18226
rect 11518 17912 11574 17921
rect 11428 17876 11480 17882
rect 11518 17847 11574 17856
rect 11428 17818 11480 17824
rect 11440 17762 11468 17818
rect 11440 17734 11652 17762
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11164 17190 11284 17218
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11164 16726 11192 17002
rect 11256 16998 11284 17190
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11242 16824 11298 16833
rect 11624 16794 11652 17734
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17338 11744 17682
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11716 17202 11744 17274
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11242 16759 11244 16768
rect 11296 16759 11298 16768
rect 11612 16788 11664 16794
rect 11244 16730 11296 16736
rect 11612 16730 11664 16736
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 16561 11284 16594
rect 11716 16590 11744 17138
rect 11808 17134 11836 18702
rect 11900 17338 11928 18770
rect 12162 17912 12218 17921
rect 12162 17847 12218 17856
rect 12176 17610 12204 17847
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11796 17128 11848 17134
rect 12164 17128 12216 17134
rect 11848 17076 12112 17082
rect 11796 17070 12112 17076
rect 12164 17070 12216 17076
rect 11808 17054 12112 17070
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11704 16584 11756 16590
rect 11242 16552 11298 16561
rect 11704 16526 11756 16532
rect 11242 16487 11298 16496
rect 11796 16516 11848 16522
rect 11796 16458 11848 16464
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11426 16144 11482 16153
rect 11808 16114 11836 16458
rect 11426 16079 11482 16088
rect 11796 16108 11848 16114
rect 11440 16046 11468 16079
rect 11796 16050 11848 16056
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11716 15706 11744 15982
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11060 14408 11112 14414
rect 10966 14376 11022 14385
rect 11060 14350 11112 14356
rect 10966 14311 11022 14320
rect 10876 14000 10928 14006
rect 10876 13942 10928 13948
rect 10876 13864 10928 13870
rect 10874 13832 10876 13841
rect 10928 13832 10930 13841
rect 10874 13767 10930 13776
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10520 13410 10548 13466
rect 10782 13424 10838 13433
rect 10520 13382 10732 13410
rect 10704 13190 10732 13382
rect 10782 13359 10784 13368
rect 10836 13359 10838 13368
rect 10784 13330 10836 13336
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10232 12980 10284 12986
rect 10336 12974 10824 13002
rect 10232 12922 10284 12928
rect 10152 12838 10456 12866
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9954 11520 10010 11529
rect 9954 11455 10010 11464
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9770 10296 9826 10305
rect 9770 10231 9826 10240
rect 9784 10198 9812 10231
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9692 9518 9720 9549
rect 9680 9512 9732 9518
rect 9600 9460 9680 9466
rect 9600 9454 9732 9460
rect 9600 9438 9720 9454
rect 9494 9344 9550 9353
rect 9494 9279 9550 9288
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9218 6896 9274 6905
rect 9218 6831 9274 6840
rect 9048 6582 9168 6610
rect 8864 6446 9076 6474
rect 8772 6310 8892 6338
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 5166 8800 5510
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8680 4950 8800 4978
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8666 3904 8722 3913
rect 8588 3670 8616 3878
rect 8666 3839 8722 3848
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8312 2922 8340 3334
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8116 2576 8168 2582
rect 8114 2544 8116 2553
rect 8168 2544 8170 2553
rect 8114 2479 8170 2488
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 8036 1698 8064 2382
rect 8024 1692 8076 1698
rect 8024 1634 8076 1640
rect 8220 1034 8248 2790
rect 8404 2650 8432 3130
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8680 1986 8708 3839
rect 8772 2854 8800 4950
rect 8864 4690 8892 6310
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8128 1006 8248 1034
rect 8588 1958 8708 1986
rect 8128 480 8156 1006
rect 8588 480 8616 1958
rect 8864 1834 8892 4626
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8956 2446 8984 3470
rect 8944 2440 8996 2446
rect 8944 2382 8996 2388
rect 8852 1828 8904 1834
rect 8852 1770 8904 1776
rect 9048 480 9076 6446
rect 9140 3754 9168 6582
rect 9232 5778 9260 6831
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9324 5846 9352 6326
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9324 4282 9352 4626
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9508 4078 9536 9279
rect 9586 9072 9642 9081
rect 9692 9042 9720 9438
rect 9586 9007 9642 9016
rect 9680 9036 9732 9042
rect 9600 8673 9628 9007
rect 9680 8978 9732 8984
rect 9876 8906 9904 10542
rect 9968 10198 9996 10746
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 9586 9996 10134
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9968 9178 9996 9318
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10060 9058 10088 12310
rect 10244 12238 10272 12650
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 10810 10180 12106
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10244 10742 10272 11290
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10140 10532 10192 10538
rect 10140 10474 10192 10480
rect 10152 10198 10180 10474
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10244 10130 10272 10678
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10266 10364 10406
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10428 10146 10456 12838
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10612 10169 10640 12310
rect 10598 10160 10654 10169
rect 10232 10124 10284 10130
rect 10428 10118 10548 10146
rect 10232 10066 10284 10072
rect 10140 9376 10192 9382
rect 10138 9344 10140 9353
rect 10192 9344 10194 9353
rect 10138 9279 10194 9288
rect 9968 9030 10088 9058
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9586 8664 9642 8673
rect 9586 8599 9642 8608
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9140 3726 9536 3754
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9218 3088 9274 3097
rect 9218 3023 9220 3032
rect 9272 3023 9274 3032
rect 9220 2994 9272 3000
rect 9324 2446 9352 3130
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9508 480 9536 3726
rect 9600 2582 9628 6938
rect 9692 6866 9720 7890
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9692 3670 9720 5102
rect 9784 4146 9812 8774
rect 9876 7342 9904 8842
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9876 5681 9904 5850
rect 9862 5672 9918 5681
rect 9862 5607 9918 5616
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9772 3528 9824 3534
rect 9770 3496 9772 3505
rect 9824 3496 9826 3505
rect 9770 3431 9826 3440
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9588 2576 9640 2582
rect 9588 2518 9640 2524
rect 9876 2446 9904 2994
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9968 480 9996 9030
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 10060 6934 10088 8842
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8022 10180 8570
rect 10244 8430 10272 10066
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10244 7954 10272 8366
rect 10232 7948 10284 7954
rect 10232 7890 10284 7896
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10048 6112 10100 6118
rect 10046 6080 10048 6089
rect 10100 6080 10102 6089
rect 10046 6015 10102 6024
rect 10152 5273 10180 7142
rect 10138 5264 10194 5273
rect 10244 5234 10272 7346
rect 10336 7274 10364 9862
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10428 9178 10456 9658
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10520 9058 10548 10118
rect 10598 10095 10654 10104
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10612 9518 10640 9590
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10428 9030 10548 9058
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5846 10364 6054
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10428 5681 10456 9030
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8537 10548 8910
rect 10506 8528 10562 8537
rect 10506 8463 10562 8472
rect 10520 6769 10548 8463
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 10612 6662 10640 8026
rect 10704 6934 10732 12310
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10704 6440 10732 6666
rect 10520 6412 10732 6440
rect 10520 6254 10548 6412
rect 10598 6352 10654 6361
rect 10598 6287 10654 6296
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10612 6186 10640 6287
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5914 10548 6054
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10414 5672 10470 5681
rect 10414 5607 10470 5616
rect 10138 5199 10194 5208
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10152 4010 10180 4966
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10244 3670 10272 4558
rect 10336 4078 10364 4558
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10428 3738 10456 4966
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10598 4176 10654 4185
rect 10508 4140 10560 4146
rect 10598 4111 10654 4120
rect 10508 4082 10560 4088
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10244 3194 10272 3606
rect 10520 3398 10548 4082
rect 10612 4010 10640 4111
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10520 3058 10548 3334
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10322 2952 10378 2961
rect 10322 2887 10378 2896
rect 10336 2854 10364 2887
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10428 2650 10456 2790
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10704 2530 10732 4762
rect 10796 2990 10824 12974
rect 10888 12442 10916 13466
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10980 11694 11008 14311
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11072 13870 11100 14214
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 13920 11652 15030
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11716 14550 11744 14758
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11716 13938 11744 14486
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11532 13892 11652 13920
rect 11704 13932 11756 13938
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11532 13734 11560 13892
rect 11704 13874 11756 13880
rect 11610 13832 11666 13841
rect 11610 13767 11666 13776
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11244 13320 11296 13326
rect 11164 13280 11244 13308
rect 11164 12696 11192 13280
rect 11244 13262 11296 13268
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11624 12832 11652 13767
rect 11808 13530 11836 13942
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11794 13424 11850 13433
rect 11704 13388 11756 13394
rect 11794 13359 11796 13368
rect 11704 13330 11756 13336
rect 11848 13359 11850 13368
rect 11796 13330 11848 13336
rect 11716 12850 11744 13330
rect 11532 12804 11652 12832
rect 11704 12844 11756 12850
rect 11244 12708 11296 12714
rect 11164 12668 11244 12696
rect 11244 12650 11296 12656
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11072 11694 11100 12242
rect 11256 12170 11284 12650
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12481 11468 12582
rect 11426 12472 11482 12481
rect 11426 12407 11482 12416
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11152 12096 11204 12102
rect 11532 12084 11560 12804
rect 11704 12786 11756 12792
rect 11900 12730 11928 16934
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15706 12020 15846
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12084 14090 12112 17054
rect 11716 12702 11928 12730
rect 11992 14062 12112 14090
rect 11716 12209 11744 12702
rect 11992 12646 12020 14062
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12084 12986 12112 13874
rect 12176 13870 12204 17070
rect 12268 16454 12296 19858
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18086 12572 19110
rect 13280 18970 13308 19178
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 12348 18080 12400 18086
rect 12532 18080 12584 18086
rect 12400 18040 12480 18068
rect 12348 18022 12400 18028
rect 12452 17338 12480 18040
rect 12820 18068 12848 18906
rect 13832 18902 13860 19858
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 12912 18170 12940 18838
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13004 18290 13032 18770
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12912 18142 13032 18170
rect 12900 18080 12952 18086
rect 12820 18040 12900 18068
rect 12532 18022 12584 18028
rect 12900 18022 12952 18028
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 12544 17354 12572 17614
rect 12440 17332 12492 17338
rect 12544 17326 12664 17354
rect 12440 17274 12492 17280
rect 12636 17270 12664 17326
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12360 15434 12388 16594
rect 12636 16590 12664 17206
rect 13004 16998 13032 18142
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12636 15502 12664 16526
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12728 15162 12756 15506
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12820 15042 12848 16934
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12912 15706 12940 15846
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12728 15014 12848 15042
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12268 14346 12296 14894
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12452 13870 12480 14418
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12452 13734 12480 13806
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 11980 12640 12032 12646
rect 11808 12588 11980 12594
rect 11808 12582 12032 12588
rect 11808 12566 12020 12582
rect 11702 12200 11758 12209
rect 11702 12135 11758 12144
rect 11532 12056 11652 12084
rect 11152 12038 11204 12044
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10888 11121 10916 11562
rect 11072 11354 11100 11630
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11286 11192 12038
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11060 11144 11112 11150
rect 10874 11112 10930 11121
rect 11256 11132 11284 11562
rect 11060 11086 11112 11092
rect 11164 11104 11284 11132
rect 10874 11047 10930 11056
rect 11072 10538 11100 11086
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 9926 11100 10474
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10874 9616 10930 9625
rect 10874 9551 10930 9560
rect 10888 9450 10916 9551
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 11072 9178 11100 9658
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11164 8945 11192 11104
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11520 9376 11572 9382
rect 11624 9353 11652 12056
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11520 9318 11572 9324
rect 11610 9344 11666 9353
rect 11532 9110 11560 9318
rect 11610 9279 11666 9288
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11520 9104 11572 9110
rect 11426 9072 11482 9081
rect 11520 9046 11572 9052
rect 11426 9007 11482 9016
rect 11244 8968 11296 8974
rect 11150 8936 11206 8945
rect 11244 8910 11296 8916
rect 11150 8871 11206 8880
rect 11256 8820 11284 8910
rect 11440 8906 11468 9007
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11164 8792 11284 8820
rect 11164 8362 11192 8792
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10888 8090 10916 8298
rect 11624 8090 11652 9114
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11624 7857 11652 7890
rect 11610 7848 11666 7857
rect 11610 7783 11666 7792
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 6934 11100 7686
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7478 11652 7783
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5914 10916 6054
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10888 4622 10916 5578
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 3505 10916 4558
rect 10874 3496 10930 3505
rect 10874 3431 10930 3440
rect 10980 3380 11008 6870
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11058 6760 11114 6769
rect 11058 6695 11060 6704
rect 11112 6695 11114 6704
rect 11060 6666 11112 6672
rect 11164 6322 11192 6802
rect 11624 6798 11652 7414
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11624 6440 11652 6734
rect 11440 6412 11652 6440
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5370 11100 6122
rect 11440 5642 11468 6412
rect 11716 6338 11744 9590
rect 11532 6310 11744 6338
rect 11532 6118 11560 6310
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11808 5896 11836 12566
rect 11992 12517 12020 12566
rect 11886 12472 11942 12481
rect 11886 12407 11888 12416
rect 11940 12407 11942 12416
rect 11888 12378 11940 12384
rect 12162 12200 12218 12209
rect 12162 12135 12218 12144
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11900 11529 11928 11630
rect 11886 11520 11942 11529
rect 11886 11455 11942 11464
rect 11900 9654 11928 11455
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 11992 11014 12020 11183
rect 12176 11132 12204 12135
rect 12084 11104 12204 11132
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 12084 10044 12112 11104
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 11992 10016 12112 10044
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11886 8936 11942 8945
rect 11886 8871 11942 8880
rect 11900 8498 11928 8871
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11992 7834 12020 10016
rect 12070 8800 12126 8809
rect 12070 8735 12126 8744
rect 12084 8566 12112 8735
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 12084 7954 12112 8502
rect 12176 8294 12204 10950
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 11992 7806 12112 7834
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11992 7410 12020 7686
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12084 7041 12112 7806
rect 12268 7154 12296 12922
rect 12452 12714 12480 13670
rect 12544 13326 12572 14214
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 13161 12572 13262
rect 12530 13152 12586 13161
rect 12530 13087 12586 13096
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12440 12708 12492 12714
rect 12440 12650 12492 12656
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12360 11898 12388 12378
rect 12452 12288 12480 12650
rect 12532 12300 12584 12306
rect 12452 12260 12532 12288
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12452 11762 12480 12260
rect 12532 12242 12584 12248
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12360 11558 12388 11698
rect 12636 11558 12664 12922
rect 12348 11552 12400 11558
rect 12532 11552 12584 11558
rect 12348 11494 12400 11500
rect 12530 11520 12532 11529
rect 12624 11552 12676 11558
rect 12584 11520 12586 11529
rect 12624 11494 12676 11500
rect 12530 11455 12586 11464
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12360 10810 12388 11086
rect 12452 10810 12480 11290
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12360 10198 12388 10746
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9466 12480 9998
rect 12544 9654 12572 11222
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12636 9489 12664 11086
rect 12728 10470 12756 15014
rect 13004 14906 13032 16934
rect 13096 15026 13124 18770
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13004 14878 13124 14906
rect 12900 14816 12952 14822
rect 12898 14784 12900 14793
rect 12952 14784 12954 14793
rect 12898 14719 12954 14728
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12912 13852 12940 14418
rect 12992 13864 13044 13870
rect 12912 13824 12992 13852
rect 12992 13806 13044 13812
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13258 12848 13670
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12806 11792 12862 11801
rect 12806 11727 12862 11736
rect 12820 11626 12848 11727
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12912 11506 12940 13330
rect 13096 12594 13124 14878
rect 12820 11478 12940 11506
rect 13004 12566 13124 12594
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10062 12756 10406
rect 12820 10305 12848 11478
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 12806 10296 12862 10305
rect 12912 10266 12940 11018
rect 12806 10231 12862 10240
rect 12900 10260 12952 10266
rect 12900 10202 12952 10208
rect 12912 10130 12940 10202
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9654 12756 9862
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12622 9480 12678 9489
rect 12452 9438 12572 9466
rect 12438 9344 12494 9353
rect 12438 9279 12494 9288
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12360 9081 12388 9114
rect 12346 9072 12402 9081
rect 12346 9007 12402 9016
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 8566 12388 8910
rect 12452 8906 12480 9279
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12346 8392 12402 8401
rect 12346 8327 12402 8336
rect 12176 7126 12296 7154
rect 12070 7032 12126 7041
rect 12070 6967 12126 6976
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11978 6080 12034 6089
rect 11900 5914 11928 6054
rect 11978 6015 12034 6024
rect 11992 5914 12020 6015
rect 11716 5868 11836 5896
rect 11888 5908 11940 5914
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4214 11100 4966
rect 11716 4826 11744 5868
rect 11888 5850 11940 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11808 5658 11836 5714
rect 11808 5630 12020 5658
rect 11992 5234 12020 5630
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11992 4826 12020 5170
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12084 4690 12112 6258
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10888 3352 11008 3380
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10796 2582 10824 2926
rect 10428 2502 10732 2530
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10428 480 10456 2502
rect 10888 480 10916 3352
rect 11072 3126 11100 3674
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2378 11100 2926
rect 11164 2650 11192 4422
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11808 4214 11836 4626
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11256 3602 11284 4082
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11336 3936 11388 3942
rect 11612 3936 11664 3942
rect 11388 3896 11612 3924
rect 11336 3878 11388 3884
rect 11612 3878 11664 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11428 3528 11480 3534
rect 11426 3496 11428 3505
rect 11480 3496 11482 3505
rect 11426 3431 11482 3440
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11244 2848 11296 2854
rect 11244 2790 11296 2796
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11256 2394 11284 2790
rect 11624 2446 11652 3606
rect 11716 2446 11744 4014
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3670 11836 3878
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 12084 3602 12112 4014
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11164 2366 11284 2394
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11164 2310 11192 2366
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11348 480 11376 1974
rect 11808 480 11836 3334
rect 12176 2038 12204 7126
rect 12254 7032 12310 7041
rect 12360 7018 12388 8327
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7342 12480 8230
rect 12440 7336 12492 7342
rect 12544 7313 12572 9438
rect 12622 9415 12678 9424
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12440 7278 12492 7284
rect 12530 7304 12586 7313
rect 12530 7239 12586 7248
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12360 6990 12480 7018
rect 12254 6967 12310 6976
rect 12268 6440 12296 6967
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12360 6662 12388 6870
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12268 6412 12388 6440
rect 12256 3596 12308 3602
rect 12360 3584 12388 6412
rect 12452 4554 12480 6990
rect 12544 5930 12572 7142
rect 12636 6118 12664 8842
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 7274 12756 8774
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12714 7168 12770 7177
rect 12714 7103 12770 7112
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12544 5902 12664 5930
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12532 3596 12584 3602
rect 12360 3556 12532 3584
rect 12256 3538 12308 3544
rect 12532 3538 12584 3544
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 12268 480 12296 3538
rect 12636 3398 12664 5902
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12544 3210 12572 3334
rect 12728 3210 12756 7103
rect 12820 6458 12848 8298
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 7546 12940 8230
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12898 7440 12954 7449
rect 12898 7375 12954 7384
rect 12912 7206 12940 7375
rect 13004 7274 13032 12566
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 13096 11694 13124 12174
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13188 11218 13216 18158
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13464 16726 13492 17070
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13634 16552 13690 16561
rect 13634 16487 13636 16496
rect 13688 16487 13690 16496
rect 13636 16458 13688 16464
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13280 15026 13308 15574
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13544 14544 13596 14550
rect 13542 14512 13544 14521
rect 13596 14512 13598 14521
rect 13542 14447 13598 14456
rect 13556 13394 13584 14447
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 13096 10470 13124 10950
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 9217 13124 10406
rect 13188 10146 13216 11154
rect 13372 10674 13400 11834
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13542 10160 13598 10169
rect 13188 10118 13400 10146
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13082 9208 13138 9217
rect 13082 9143 13138 9152
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 7410 13124 8910
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 13004 6882 13032 7210
rect 13096 7002 13124 7346
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12900 6860 12952 6866
rect 13004 6854 13124 6882
rect 12900 6802 12952 6808
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12912 5642 12940 6802
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4826 12940 4966
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13004 4706 13032 6734
rect 12912 4678 13032 4706
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12820 3466 12848 3946
rect 12912 3534 12940 4678
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 12544 3182 12756 3210
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12728 480 12756 3062
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 12912 2378 12940 2790
rect 13096 2514 13124 6854
rect 13188 6361 13216 9998
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13280 8809 13308 8910
rect 13266 8800 13322 8809
rect 13266 8735 13322 8744
rect 13280 8498 13308 8735
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13372 8378 13400 10118
rect 13452 10124 13504 10130
rect 13542 10095 13598 10104
rect 13452 10066 13504 10072
rect 13464 8906 13492 10066
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13280 8350 13400 8378
rect 13280 6798 13308 8350
rect 13452 7880 13504 7886
rect 13450 7848 13452 7857
rect 13504 7848 13506 7857
rect 13450 7783 13506 7792
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6934 13400 7142
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13268 6656 13320 6662
rect 13320 6616 13400 6644
rect 13268 6598 13320 6604
rect 13174 6352 13230 6361
rect 13174 6287 13230 6296
rect 13188 6118 13216 6287
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13280 5574 13308 5782
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13372 4706 13400 6616
rect 13464 6236 13492 7783
rect 13556 7410 13584 10095
rect 13648 9586 13676 14894
rect 13740 13954 13768 18022
rect 13832 17882 13860 18226
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13832 17218 13860 17478
rect 13924 17338 13952 20046
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14004 19304 14056 19310
rect 14004 19246 14056 19252
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 13832 17190 13952 17218
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13832 15570 13860 16050
rect 13924 15978 13952 17190
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14482 13860 14962
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 14074 13860 14418
rect 14016 14278 14044 19246
rect 14200 18902 14228 19858
rect 14292 19174 14320 22320
rect 14752 20754 14780 22320
rect 14568 20726 14780 20754
rect 14568 20058 14596 20726
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15212 20058 15240 22320
rect 15672 20058 15700 22320
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13740 13926 14044 13954
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13740 9466 13768 13126
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13832 11558 13860 12650
rect 13912 12368 13964 12374
rect 13910 12336 13912 12345
rect 13964 12336 13966 12345
rect 13910 12271 13966 12280
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11665 13952 12038
rect 13910 11656 13966 11665
rect 13910 11591 13966 11600
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 10742 13860 11494
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 9636 13860 10406
rect 13832 9608 13952 9636
rect 13924 9489 13952 9608
rect 13910 9480 13966 9489
rect 13740 9438 13860 9466
rect 13832 9058 13860 9438
rect 13910 9415 13966 9424
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9178 13952 9318
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13740 9030 13860 9058
rect 13740 8362 13768 9030
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13832 8022 13860 8910
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13740 7750 13768 7890
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 13740 6866 13768 7346
rect 13832 7274 13860 7958
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13924 7206 13952 8230
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 6458 13860 6666
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13636 6248 13688 6254
rect 13464 6208 13636 6236
rect 13464 5794 13492 6208
rect 13636 6190 13688 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13464 5778 13584 5794
rect 13832 5778 13860 6054
rect 13464 5772 13596 5778
rect 13464 5766 13544 5772
rect 13544 5714 13596 5720
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13452 5704 13504 5710
rect 13504 5652 13860 5658
rect 13452 5646 13860 5652
rect 13464 5630 13860 5646
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13268 4684 13320 4690
rect 13372 4678 13492 4706
rect 13268 4626 13320 4632
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 13188 480 13216 3878
rect 13280 2854 13308 4626
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13372 3738 13400 4558
rect 13464 4214 13492 4678
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 4486 13584 4558
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13556 4282 13584 4422
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13464 3074 13492 4150
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13372 3058 13492 3074
rect 13360 3052 13492 3058
rect 13412 3046 13492 3052
rect 13360 2994 13412 3000
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13556 2446 13584 3470
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13556 2106 13584 2382
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13648 480 13676 4966
rect 13832 3670 13860 5630
rect 13924 4758 13952 7142
rect 14016 4758 14044 13926
rect 14108 12481 14136 18022
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14292 17202 14320 17682
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14292 17082 14320 17138
rect 14200 17054 14320 17082
rect 14200 13394 14228 17054
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14292 16250 14320 16594
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14188 13388 14240 13394
rect 14188 13330 14240 13336
rect 14200 12850 14228 13330
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14094 12472 14150 12481
rect 14094 12407 14150 12416
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14094 11792 14150 11801
rect 14094 11727 14150 11736
rect 14108 10062 14136 11727
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14200 9625 14228 12378
rect 14292 12345 14320 12854
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14384 11914 14412 14894
rect 14476 12102 14504 19858
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15014 15600 15070 15609
rect 14556 15564 14608 15570
rect 15014 15535 15070 15544
rect 14556 15506 14608 15512
rect 14568 15026 14596 15506
rect 15028 15162 15056 15535
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14568 14346 14596 14962
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 15106 13968 15162 13977
rect 15106 13903 15162 13912
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15028 13530 15056 13670
rect 15120 13530 15148 13903
rect 14556 13524 14608 13530
rect 15016 13524 15068 13530
rect 14608 13484 14688 13512
rect 14556 13466 14608 13472
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14568 12782 14596 13262
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14660 12628 14688 13484
rect 15016 13466 15068 13472
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12782 14964 13126
rect 15028 12782 15056 13194
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14924 12776 14976 12782
rect 14924 12718 14976 12724
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14568 12600 14688 12628
rect 15016 12640 15068 12646
rect 14568 12442 14596 12600
rect 15016 12582 15068 12588
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14384 11886 14504 11914
rect 14936 11898 14964 12038
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14370 11520 14426 11529
rect 14292 10606 14320 11494
rect 14370 11455 14426 11464
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 14384 10554 14412 11455
rect 14476 11336 14504 11886
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14646 11792 14702 11801
rect 14646 11727 14648 11736
rect 14700 11727 14702 11736
rect 14648 11698 14700 11704
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14476 11308 14964 11336
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14476 10810 14504 11154
rect 14556 11144 14608 11150
rect 14648 11144 14700 11150
rect 14556 11086 14608 11092
rect 14646 11112 14648 11121
rect 14700 11112 14702 11121
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14384 10526 14504 10554
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14278 10296 14334 10305
rect 14384 10266 14412 10406
rect 14278 10231 14334 10240
rect 14372 10260 14424 10266
rect 14186 9616 14242 9625
rect 14096 9580 14148 9586
rect 14186 9551 14242 9560
rect 14096 9522 14148 9528
rect 14108 8634 14136 9522
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14200 8430 14228 9454
rect 14292 8974 14320 10231
rect 14372 10202 14424 10208
rect 14476 9602 14504 10526
rect 14384 9574 14504 9602
rect 14384 9178 14412 9574
rect 14568 9466 14596 11086
rect 14646 11047 14702 11056
rect 14936 10588 14964 11308
rect 15028 10742 15056 12582
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15120 10674 15148 12786
rect 15304 11257 15332 18770
rect 15382 15056 15438 15065
rect 15382 14991 15438 15000
rect 15396 14890 15424 14991
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 15488 14618 15516 19858
rect 15580 18902 15608 19858
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 14936 10560 15056 10588
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14476 9438 14596 9466
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8498 14320 8910
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14108 6769 14136 7346
rect 14094 6760 14150 6769
rect 14094 6695 14150 6704
rect 14094 6216 14150 6225
rect 14094 6151 14150 6160
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 14108 4706 14136 6151
rect 14200 6118 14228 7686
rect 14384 7274 14412 9114
rect 14476 8090 14504 9438
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8634 14596 9318
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 15028 7562 15056 10560
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14568 7534 15056 7562
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 7002 14504 7142
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14292 6730 14320 6938
rect 14568 6882 14596 7534
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14384 6854 14596 6882
rect 15016 6860 15068 6866
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5370 14228 6054
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14200 5114 14228 5306
rect 14200 5086 14320 5114
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4826 14228 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14108 4678 14228 4706
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 2990 13952 3538
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14016 2514 14044 3470
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14004 2508 14056 2514
rect 14004 2450 14056 2456
rect 14108 480 14136 3334
rect 14200 2514 14228 4678
rect 14292 4622 14320 5086
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14384 3210 14412 6854
rect 15016 6802 15068 6808
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14476 5234 14504 6122
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 14568 5166 14596 6734
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14830 5264 14886 5273
rect 14936 5234 14964 5510
rect 14830 5199 14886 5208
rect 14924 5228 14976 5234
rect 14844 5166 14872 5199
rect 14924 5170 14976 5176
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14462 4176 14518 4185
rect 14462 4111 14518 4120
rect 14476 4078 14504 4111
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14292 3182 14412 3210
rect 14568 4010 14688 4026
rect 15028 4010 15056 6802
rect 15120 6730 15148 9454
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5710 15332 6054
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 14568 4004 14700 4010
rect 14568 3998 14648 4004
rect 14292 3126 14320 3182
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14568 480 14596 3998
rect 14648 3946 14700 3952
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15120 2990 15148 4694
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14740 2984 14792 2990
rect 14738 2952 14740 2961
rect 15108 2984 15160 2990
rect 14792 2952 14794 2961
rect 15108 2926 15160 2932
rect 15212 2922 15240 4626
rect 14738 2887 14794 2896
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15304 2514 15332 5510
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4758 15424 4966
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15488 3641 15516 14554
rect 15580 12646 15608 18702
rect 15764 14385 15792 19178
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15948 14414 15976 14962
rect 15936 14408 15988 14414
rect 15750 14376 15806 14385
rect 15936 14350 15988 14356
rect 15750 14311 15806 14320
rect 15948 13802 15976 14350
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15672 8537 15700 13330
rect 15948 13326 15976 13738
rect 16040 13734 16068 19246
rect 16132 19174 16160 22320
rect 16592 20058 16620 22320
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 16592 11014 16620 19246
rect 16670 13832 16726 13841
rect 16670 13767 16726 13776
rect 16684 13530 16712 13767
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11354 16712 11630
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16776 9722 16804 13262
rect 16868 11082 16896 19246
rect 17052 19174 17080 22320
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17144 12986 17172 19858
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17236 11762 17264 19246
rect 17512 19174 17540 22320
rect 17972 20058 18000 22320
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18432 19802 18460 22320
rect 18432 19774 18552 19802
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19174 18552 19774
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 17972 9654 18000 18770
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18524 17241 18552 17614
rect 18510 17232 18566 17241
rect 18510 17167 18566 17176
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18616 14822 18644 19246
rect 18708 18902 18736 19246
rect 18892 19174 18920 22320
rect 19352 19786 19380 22320
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 19352 17338 19380 18906
rect 19812 18630 19840 22320
rect 20272 19174 20300 22320
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19432 18080 19484 18086
rect 20732 18068 20760 22320
rect 21192 18970 21220 22320
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21652 18426 21680 22320
rect 22112 19242 22140 22320
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 22572 18086 22600 22320
rect 19432 18022 19484 18028
rect 20640 18040 20760 18068
rect 22560 18080 22612 18086
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 19444 14618 19472 18022
rect 20640 17882 20668 18040
rect 22560 18022 22612 18028
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 15658 8528 15714 8537
rect 15658 8463 15714 8472
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15764 6866 15792 7414
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5846 15608 6054
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15580 5234 15608 5782
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15764 4690 15792 6394
rect 15856 6254 15884 6734
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 15856 5914 15884 6054
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16224 5370 16252 6054
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 15936 5092 15988 5098
rect 15936 5034 15988 5040
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15948 4146 15976 5034
rect 16316 4826 16344 6054
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15474 3632 15530 3641
rect 15384 3596 15436 3602
rect 15474 3567 15530 3576
rect 15384 3538 15436 3544
rect 15396 3058 15424 3538
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14844 2310 14872 2450
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 15028 480 15056 2314
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15580 480 15608 2246
rect 16040 480 16068 3062
rect 16132 2990 16160 3470
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16592 2514 16620 6870
rect 16960 5234 16988 7346
rect 17498 6896 17554 6905
rect 17498 6831 17554 6840
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 3738 16804 4966
rect 16960 4622 16988 5170
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 17052 2990 17080 4490
rect 17144 2990 17172 6666
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 5846 17356 6598
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16500 480 16528 2246
rect 16960 480 16988 2790
rect 17512 2514 17540 6831
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18708 5817 18736 13806
rect 17958 5808 18014 5817
rect 17958 5743 17960 5752
rect 18012 5743 18014 5752
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 17960 5714 18012 5720
rect 19800 5704 19852 5710
rect 18878 5672 18934 5681
rect 19800 5646 19852 5652
rect 18878 5607 18934 5616
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17420 480 17448 2246
rect 17880 480 17908 2790
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 1170 18000 2246
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18368 1170
rect 18340 480 18368 1142
rect 18800 480 18828 4422
rect 18892 2990 18920 5607
rect 19812 5166 19840 5646
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 19248 3120 19300 3126
rect 19248 3062 19300 3068
rect 18880 2984 18932 2990
rect 18880 2926 18932 2932
rect 19260 480 19288 3062
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19720 480 19748 2790
rect 19812 2650 19840 2790
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 20168 2576 20220 2582
rect 20168 2518 20220 2524
rect 20180 480 20208 2518
rect 20640 480 20668 4966
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21100 480 21128 3130
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21560 480 21588 2790
rect 22020 480 22048 2858
rect 22480 480 22508 2994
rect 4158 232 4214 241
rect 4158 167 4214 176
rect 4342 0 4398 480
rect 4802 0 4858 480
rect 5262 0 5318 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6642 0 6698 480
rect 7102 0 7158 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8574 0 8630 480
rect 9034 0 9090 480
rect 9494 0 9550 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13634 0 13690 480
rect 14094 0 14150 480
rect 14554 0 14610 480
rect 15014 0 15070 480
rect 15566 0 15622 480
rect 16026 0 16082 480
rect 16486 0 16542 480
rect 16946 0 17002 480
rect 17406 0 17462 480
rect 17866 0 17922 480
rect 18326 0 18382 480
rect 18786 0 18842 480
rect 19246 0 19302 480
rect 19706 0 19762 480
rect 20166 0 20222 480
rect 20626 0 20682 480
rect 21086 0 21142 480
rect 21546 0 21602 480
rect 22006 0 22062 480
rect 22466 0 22522 480
<< via2 >>
rect 3238 22480 3294 22536
rect 1858 19660 1860 19680
rect 1860 19660 1912 19680
rect 1912 19660 1914 19680
rect 1858 19624 1914 19660
rect 1766 19216 1822 19272
rect 1582 18692 1638 18728
rect 1582 18672 1584 18692
rect 1584 18672 1636 18692
rect 1636 18672 1638 18692
rect 1674 18300 1676 18320
rect 1676 18300 1728 18320
rect 1728 18300 1730 18320
rect 1674 18264 1730 18300
rect 1766 17332 1822 17368
rect 1766 17312 1768 17332
rect 1768 17312 1820 17332
rect 1820 17312 1822 17332
rect 1582 16360 1638 16416
rect 1398 16088 1454 16144
rect 1858 16788 1914 16824
rect 1858 16768 1860 16788
rect 1860 16768 1912 16788
rect 1912 16768 1914 16788
rect 2410 18264 2466 18320
rect 1950 15952 2006 16008
rect 1582 15816 1638 15872
rect 2870 15816 2926 15872
rect 2410 15564 2466 15600
rect 2410 15544 2412 15564
rect 2412 15544 2464 15564
rect 2464 15544 2466 15564
rect 1674 14864 1730 14920
rect 1398 10648 1454 10704
rect 3146 17720 3202 17776
rect 3054 15680 3110 15736
rect 3514 21528 3570 21584
rect 3422 19216 3478 19272
rect 3330 18028 3332 18048
rect 3332 18028 3384 18048
rect 3384 18028 3386 18048
rect 3330 17992 3386 18028
rect 3698 21120 3754 21176
rect 3974 22072 4030 22128
rect 3882 20596 3938 20632
rect 3882 20576 3884 20596
rect 3884 20576 3936 20596
rect 3936 20576 3938 20596
rect 3790 18672 3846 18728
rect 3606 16532 3608 16552
rect 3608 16532 3660 16552
rect 3660 16532 3662 16552
rect 3606 16496 3662 16532
rect 3974 20168 4030 20224
rect 3882 17040 3938 17096
rect 4066 18536 4122 18592
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4342 19216 4398 19272
rect 4618 18808 4674 18864
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3514 15680 3570 15736
rect 3422 15408 3478 15464
rect 2962 12416 3018 12472
rect 2410 7284 2412 7304
rect 2412 7284 2464 7304
rect 2464 7284 2466 7304
rect 2410 7248 2466 7284
rect 3330 14456 3386 14512
rect 3698 15000 3754 15056
rect 2778 3984 2834 4040
rect 2962 3032 3018 3088
rect 3146 5752 3202 5808
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 3974 13912 4030 13968
rect 3790 12960 3846 13016
rect 3606 12552 3662 12608
rect 3790 9288 3846 9344
rect 3146 3848 3202 3904
rect 3054 2080 3110 2136
rect 2778 1128 2834 1184
rect 3330 1536 3386 1592
rect 4526 15952 4582 16008
rect 4434 15816 4490 15872
rect 4526 15408 4582 15464
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4894 15852 4896 15872
rect 4896 15852 4948 15872
rect 4948 15852 4950 15872
rect 4894 15816 4950 15852
rect 4250 14320 4306 14376
rect 4802 14320 4858 14376
rect 4066 13504 4122 13560
rect 3974 12300 4030 12336
rect 3974 12280 3976 12300
rect 3976 12280 4028 12300
rect 4028 12280 4030 12300
rect 5078 18028 5080 18048
rect 5080 18028 5132 18048
rect 5132 18028 5134 18048
rect 5078 17992 5134 18028
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4250 12688 4306 12744
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4250 11600 4306 11656
rect 4894 14068 4950 14104
rect 4894 14048 4896 14068
rect 4896 14048 4948 14068
rect 4948 14048 4950 14068
rect 5538 18808 5594 18864
rect 5262 16940 5264 16960
rect 5264 16940 5316 16960
rect 5316 16940 5318 16960
rect 5262 16904 5318 16940
rect 5446 16496 5502 16552
rect 5354 13776 5410 13832
rect 4986 11736 5042 11792
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4618 10240 4674 10296
rect 4526 10124 4582 10160
rect 4526 10104 4528 10124
rect 4528 10104 4580 10124
rect 4580 10104 4582 10124
rect 4894 10512 4950 10568
rect 4250 9968 4306 10024
rect 3974 9716 4030 9752
rect 3974 9696 3976 9716
rect 3976 9696 4028 9716
rect 4028 9696 4030 9716
rect 3974 8744 4030 8800
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 3974 8200 4030 8256
rect 4066 7812 4122 7848
rect 4066 7792 4068 7812
rect 4068 7792 4120 7812
rect 4120 7792 4122 7812
rect 4066 6840 4122 6896
rect 3974 5344 4030 5400
rect 4066 4936 4122 4992
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4526 5888 4582 5944
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 5170 10004 5172 10024
rect 5172 10004 5224 10024
rect 5224 10004 5226 10024
rect 5170 9968 5226 10004
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 5722 15816 5778 15872
rect 6918 18264 6974 18320
rect 5998 17040 6054 17096
rect 5998 15952 6054 16008
rect 5906 15680 5962 15736
rect 5906 14864 5962 14920
rect 5814 10240 5870 10296
rect 4894 3440 4950 3496
rect 4066 2488 4122 2544
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5170 3476 5172 3496
rect 5172 3476 5224 3496
rect 5224 3476 5226 3496
rect 5170 3440 5226 3476
rect 5446 2488 5502 2544
rect 5538 584 5594 640
rect 5814 2916 5870 2952
rect 5814 2896 5816 2916
rect 5816 2896 5868 2916
rect 5868 2896 5870 2916
rect 6826 16088 6882 16144
rect 7286 15000 7342 15056
rect 7010 12416 7066 12472
rect 6642 10648 6698 10704
rect 6274 10412 6276 10432
rect 6276 10412 6328 10432
rect 6328 10412 6330 10432
rect 6274 10376 6330 10412
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7562 16904 7618 16960
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 8574 19216 8630 19272
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7562 14048 7618 14104
rect 7378 12416 7434 12472
rect 7286 12144 7342 12200
rect 6090 4528 6146 4584
rect 6182 3576 6238 3632
rect 7010 8608 7066 8664
rect 6918 6160 6974 6216
rect 6734 4020 6736 4040
rect 6736 4020 6788 4040
rect 6788 4020 6790 4040
rect 6734 3984 6790 4020
rect 7286 9288 7342 9344
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7654 11600 7710 11656
rect 7102 3884 7104 3904
rect 7104 3884 7156 3904
rect 7156 3884 7158 3904
rect 7102 3848 7158 3884
rect 7286 3068 7288 3088
rect 7288 3068 7340 3088
rect 7340 3068 7342 3088
rect 7286 3032 7342 3068
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8298 10648 8354 10704
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 8482 12688 8538 12744
rect 8666 11056 8722 11112
rect 8574 10104 8630 10160
rect 8482 9424 8538 9480
rect 7930 7384 7986 7440
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7930 4700 7932 4720
rect 7932 4700 7984 4720
rect 7984 4700 7986 4720
rect 7930 4664 7986 4700
rect 7930 4548 7986 4584
rect 7930 4528 7932 4548
rect 7932 4528 7984 4548
rect 7984 4528 7986 4548
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 8942 15408 8998 15464
rect 9034 14728 9090 14784
rect 8850 13776 8906 13832
rect 8666 8916 8668 8936
rect 8668 8916 8720 8936
rect 8720 8916 8722 8936
rect 8666 8880 8722 8916
rect 8758 8336 8814 8392
rect 10046 15952 10102 16008
rect 9954 15036 9956 15056
rect 9956 15036 10008 15056
rect 10008 15036 10010 15056
rect 9954 15000 10010 15036
rect 9954 13912 10010 13968
rect 9678 12280 9734 12336
rect 9586 12008 9642 12064
rect 9402 10548 9404 10568
rect 9404 10548 9456 10568
rect 9456 10548 9458 10568
rect 9218 10104 9274 10160
rect 9402 10512 9458 10548
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 10782 16768 10838 16824
rect 10966 14492 10968 14512
rect 10968 14492 11020 14512
rect 11020 14492 11022 14512
rect 10966 14456 11022 14492
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11518 17856 11574 17912
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11242 16788 11298 16824
rect 11242 16768 11244 16788
rect 11244 16768 11296 16788
rect 11296 16768 11298 16788
rect 12162 17856 12218 17912
rect 11242 16496 11298 16552
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11426 16088 11482 16144
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 10966 14320 11022 14376
rect 10874 13812 10876 13832
rect 10876 13812 10928 13832
rect 10928 13812 10930 13832
rect 10874 13776 10930 13812
rect 10782 13388 10838 13424
rect 10782 13368 10784 13388
rect 10784 13368 10836 13388
rect 10836 13368 10838 13388
rect 9954 11464 10010 11520
rect 9770 10240 9826 10296
rect 9494 9288 9550 9344
rect 9218 6840 9274 6896
rect 8666 3848 8722 3904
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8114 2524 8116 2544
rect 8116 2524 8168 2544
rect 8168 2524 8170 2544
rect 8114 2488 8170 2524
rect 9586 9016 9642 9072
rect 10138 9324 10140 9344
rect 10140 9324 10192 9344
rect 10192 9324 10194 9344
rect 10138 9288 10194 9324
rect 9586 8608 9642 8664
rect 9218 3052 9274 3088
rect 9218 3032 9220 3052
rect 9220 3032 9272 3052
rect 9272 3032 9274 3052
rect 9862 5616 9918 5672
rect 9770 3476 9772 3496
rect 9772 3476 9824 3496
rect 9824 3476 9826 3496
rect 9770 3440 9826 3476
rect 10046 6060 10048 6080
rect 10048 6060 10100 6080
rect 10100 6060 10102 6080
rect 10046 6024 10102 6060
rect 10138 5208 10194 5264
rect 10598 10104 10654 10160
rect 10506 8472 10562 8528
rect 10506 6704 10562 6760
rect 10598 6296 10654 6352
rect 10414 5616 10470 5672
rect 10598 4120 10654 4176
rect 10322 2896 10378 2952
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11610 13776 11666 13832
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11794 13388 11850 13424
rect 11794 13368 11796 13388
rect 11796 13368 11848 13388
rect 11848 13368 11850 13388
rect 11426 12416 11482 12472
rect 11702 12144 11758 12200
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 10874 11056 10930 11112
rect 10874 9560 10930 9616
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11610 9288 11666 9344
rect 11426 9016 11482 9072
rect 11150 8880 11206 8936
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11610 7792 11666 7848
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 10874 3440 10930 3496
rect 11058 6724 11114 6760
rect 11058 6704 11060 6724
rect 11060 6704 11112 6724
rect 11112 6704 11114 6724
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11886 12436 11942 12472
rect 11886 12416 11888 12436
rect 11888 12416 11940 12436
rect 11940 12416 11942 12436
rect 12162 12144 12218 12200
rect 11886 11464 11942 11520
rect 11978 11192 12034 11248
rect 11886 8880 11942 8936
rect 12070 8744 12126 8800
rect 12530 13096 12586 13152
rect 12530 11500 12532 11520
rect 12532 11500 12584 11520
rect 12584 11500 12586 11520
rect 12530 11464 12586 11500
rect 12898 14764 12900 14784
rect 12900 14764 12952 14784
rect 12952 14764 12954 14784
rect 12898 14728 12954 14764
rect 12806 11736 12862 11792
rect 12806 10240 12862 10296
rect 12438 9288 12494 9344
rect 12346 9016 12402 9072
rect 12346 8336 12402 8392
rect 12070 6976 12126 7032
rect 11978 6024 12034 6080
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11426 3476 11428 3496
rect 11428 3476 11480 3496
rect 11480 3476 11482 3496
rect 11426 3440 11482 3476
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12254 6976 12310 7032
rect 12622 9424 12678 9480
rect 12530 7248 12586 7304
rect 12714 7112 12770 7168
rect 12898 7384 12954 7440
rect 13634 16516 13690 16552
rect 13634 16496 13636 16516
rect 13636 16496 13688 16516
rect 13688 16496 13690 16516
rect 13542 14492 13544 14512
rect 13544 14492 13596 14512
rect 13596 14492 13598 14512
rect 13542 14456 13598 14492
rect 13082 9152 13138 9208
rect 13266 8744 13322 8800
rect 13542 10104 13598 10160
rect 13450 7828 13452 7848
rect 13452 7828 13504 7848
rect 13504 7828 13506 7848
rect 13450 7792 13506 7828
rect 13174 6296 13230 6352
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13910 12316 13912 12336
rect 13912 12316 13964 12336
rect 13964 12316 13966 12336
rect 13910 12280 13966 12316
rect 13910 11600 13966 11656
rect 13910 9424 13966 9480
rect 14094 12416 14150 12472
rect 14094 11736 14150 11792
rect 14278 12280 14334 12336
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 15014 15544 15070 15600
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 15106 13912 15162 13968
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14370 11464 14426 11520
rect 14646 11756 14702 11792
rect 14646 11736 14648 11756
rect 14648 11736 14700 11756
rect 14700 11736 14702 11756
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14646 11092 14648 11112
rect 14648 11092 14700 11112
rect 14700 11092 14702 11112
rect 14278 10240 14334 10296
rect 14186 9560 14242 9616
rect 14646 11056 14702 11092
rect 15382 15000 15438 15056
rect 15290 11192 15346 11248
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14094 6704 14150 6760
rect 14094 6160 14150 6216
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14830 5208 14886 5264
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14462 4120 14518 4176
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14738 2932 14740 2952
rect 14740 2932 14792 2952
rect 14792 2932 14794 2952
rect 14738 2896 14794 2932
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15750 14320 15806 14376
rect 16670 13776 16726 13832
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18510 17176 18566 17232
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 15658 8472 15714 8528
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 15474 3576 15530 3632
rect 17498 6840 17554 6896
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 5772 18014 5808
rect 17958 5752 17960 5772
rect 17960 5752 18012 5772
rect 18012 5752 18014 5772
rect 18694 5752 18750 5808
rect 18878 5616 18934 5672
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 4158 176 4214 232
<< metal3 >>
rect 0 22538 480 22568
rect 3233 22538 3299 22541
rect 0 22536 3299 22538
rect 0 22480 3238 22536
rect 3294 22480 3299 22536
rect 0 22478 3299 22480
rect 0 22448 480 22478
rect 3233 22475 3299 22478
rect 0 22130 480 22160
rect 3969 22130 4035 22133
rect 0 22128 4035 22130
rect 0 22072 3974 22128
rect 4030 22072 4035 22128
rect 0 22070 4035 22072
rect 0 22040 480 22070
rect 3969 22067 4035 22070
rect 0 21586 480 21616
rect 3509 21586 3575 21589
rect 0 21584 3575 21586
rect 0 21528 3514 21584
rect 3570 21528 3575 21584
rect 0 21526 3575 21528
rect 0 21496 480 21526
rect 3509 21523 3575 21526
rect 0 21178 480 21208
rect 3693 21178 3759 21181
rect 0 21176 3759 21178
rect 0 21120 3698 21176
rect 3754 21120 3759 21176
rect 0 21118 3759 21120
rect 0 21088 480 21118
rect 3693 21115 3759 21118
rect 0 20634 480 20664
rect 3877 20634 3943 20637
rect 0 20632 3943 20634
rect 0 20576 3882 20632
rect 3938 20576 3943 20632
rect 0 20574 3943 20576
rect 0 20544 480 20574
rect 3877 20571 3943 20574
rect 0 20226 480 20256
rect 3969 20226 4035 20229
rect 0 20224 4035 20226
rect 0 20168 3974 20224
rect 4030 20168 4035 20224
rect 0 20166 4035 20168
rect 0 20136 480 20166
rect 3969 20163 4035 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19682 480 19712
rect 1853 19682 1919 19685
rect 0 19680 1919 19682
rect 0 19624 1858 19680
rect 1914 19624 1919 19680
rect 0 19622 1919 19624
rect 0 19592 480 19622
rect 1853 19619 1919 19622
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 1761 19274 1827 19277
rect 0 19272 1827 19274
rect 0 19216 1766 19272
rect 1822 19216 1827 19272
rect 0 19214 1827 19216
rect 0 19184 480 19214
rect 1761 19211 1827 19214
rect 3417 19274 3483 19277
rect 4337 19274 4403 19277
rect 8569 19274 8635 19277
rect 3417 19272 3618 19274
rect 3417 19216 3422 19272
rect 3478 19216 3618 19272
rect 3417 19214 3618 19216
rect 3417 19211 3483 19214
rect 0 18730 480 18760
rect 1577 18730 1643 18733
rect 0 18728 1643 18730
rect 0 18672 1582 18728
rect 1638 18672 1643 18728
rect 0 18670 1643 18672
rect 3558 18730 3618 19214
rect 4337 19272 8635 19274
rect 4337 19216 4342 19272
rect 4398 19216 8574 19272
rect 8630 19216 8635 19272
rect 4337 19214 8635 19216
rect 4337 19211 4403 19214
rect 8569 19211 8635 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 4613 18866 4679 18869
rect 5533 18866 5599 18869
rect 4064 18864 5599 18866
rect 4064 18808 4618 18864
rect 4674 18808 5538 18864
rect 5594 18808 5599 18864
rect 4064 18806 5599 18808
rect 3785 18730 3851 18733
rect 3558 18728 3851 18730
rect 3558 18672 3790 18728
rect 3846 18672 3851 18728
rect 3558 18670 3851 18672
rect 0 18640 480 18670
rect 1577 18667 1643 18670
rect 3785 18667 3851 18670
rect 4064 18597 4124 18806
rect 4613 18803 4679 18806
rect 5533 18803 5599 18806
rect 4061 18592 4127 18597
rect 4061 18536 4066 18592
rect 4122 18536 4127 18592
rect 4061 18531 4127 18536
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1669 18322 1735 18325
rect 0 18320 1735 18322
rect 0 18264 1674 18320
rect 1730 18264 1735 18320
rect 0 18262 1735 18264
rect 0 18232 480 18262
rect 1669 18259 1735 18262
rect 2405 18322 2471 18325
rect 6913 18322 6979 18325
rect 2405 18320 6979 18322
rect 2405 18264 2410 18320
rect 2466 18264 6918 18320
rect 6974 18264 6979 18320
rect 2405 18262 6979 18264
rect 2405 18259 2471 18262
rect 6913 18259 6979 18262
rect 3325 18050 3391 18053
rect 5073 18050 5139 18053
rect 3325 18048 5139 18050
rect 3325 17992 3330 18048
rect 3386 17992 5078 18048
rect 5134 17992 5139 18048
rect 3325 17990 5139 17992
rect 3325 17987 3391 17990
rect 5073 17987 5139 17990
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 11513 17914 11579 17917
rect 12157 17914 12223 17917
rect 11513 17912 12223 17914
rect 11513 17856 11518 17912
rect 11574 17856 12162 17912
rect 12218 17856 12223 17912
rect 11513 17854 12223 17856
rect 11513 17851 11579 17854
rect 12157 17851 12223 17854
rect 0 17778 480 17808
rect 3141 17778 3207 17781
rect 0 17776 3207 17778
rect 0 17720 3146 17776
rect 3202 17720 3207 17776
rect 0 17718 3207 17720
rect 0 17688 480 17718
rect 3141 17715 3207 17718
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1761 17370 1827 17373
rect 0 17368 1827 17370
rect 0 17312 1766 17368
rect 1822 17312 1827 17368
rect 0 17310 1827 17312
rect 0 17280 480 17310
rect 1761 17307 1827 17310
rect 18505 17234 18571 17237
rect 22320 17234 22800 17264
rect 18505 17232 22800 17234
rect 18505 17176 18510 17232
rect 18566 17176 22800 17232
rect 18505 17174 22800 17176
rect 18505 17171 18571 17174
rect 22320 17144 22800 17174
rect 3877 17098 3943 17101
rect 5993 17098 6059 17101
rect 3877 17096 6059 17098
rect 3877 17040 3882 17096
rect 3938 17040 5998 17096
rect 6054 17040 6059 17096
rect 3877 17038 6059 17040
rect 3877 17035 3943 17038
rect 5993 17035 6059 17038
rect 5257 16964 5323 16965
rect 5206 16900 5212 16964
rect 5276 16962 5323 16964
rect 7557 16962 7623 16965
rect 5276 16960 7623 16962
rect 5318 16904 7562 16960
rect 7618 16904 7623 16960
rect 5276 16902 7623 16904
rect 5276 16900 5323 16902
rect 5257 16899 5323 16900
rect 7557 16899 7623 16902
rect 7808 16896 8128 16897
rect 0 16826 480 16856
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 1853 16826 1919 16829
rect 0 16824 1919 16826
rect 0 16768 1858 16824
rect 1914 16768 1919 16824
rect 0 16766 1919 16768
rect 0 16736 480 16766
rect 1853 16763 1919 16766
rect 10777 16826 10843 16829
rect 11237 16826 11303 16829
rect 10777 16824 11303 16826
rect 10777 16768 10782 16824
rect 10838 16768 11242 16824
rect 11298 16768 11303 16824
rect 10777 16766 11303 16768
rect 10777 16763 10843 16766
rect 11237 16763 11303 16766
rect 3601 16554 3667 16557
rect 5441 16554 5507 16557
rect 3601 16552 5507 16554
rect 3601 16496 3606 16552
rect 3662 16496 5446 16552
rect 5502 16496 5507 16552
rect 3601 16494 5507 16496
rect 3601 16491 3667 16494
rect 5441 16491 5507 16494
rect 11237 16554 11303 16557
rect 13629 16554 13695 16557
rect 11237 16552 13695 16554
rect 11237 16496 11242 16552
rect 11298 16496 13634 16552
rect 13690 16496 13695 16552
rect 11237 16494 13695 16496
rect 11237 16491 11303 16494
rect 13629 16491 13695 16494
rect 0 16418 480 16448
rect 1577 16418 1643 16421
rect 0 16416 1643 16418
rect 0 16360 1582 16416
rect 1638 16360 1643 16416
rect 0 16358 1643 16360
rect 0 16328 480 16358
rect 1577 16355 1643 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 1393 16146 1459 16149
rect 6821 16146 6887 16149
rect 11421 16146 11487 16149
rect 1393 16144 6378 16146
rect 1393 16088 1398 16144
rect 1454 16088 6378 16144
rect 1393 16086 6378 16088
rect 1393 16083 1459 16086
rect 1945 16010 2011 16013
rect 4521 16010 4587 16013
rect 5993 16010 6059 16013
rect 1945 16008 4587 16010
rect 1945 15952 1950 16008
rect 2006 15952 4526 16008
rect 4582 15952 4587 16008
rect 1945 15950 4587 15952
rect 1945 15947 2011 15950
rect 4521 15947 4587 15950
rect 4662 16008 6059 16010
rect 4662 15952 5998 16008
rect 6054 15952 6059 16008
rect 4662 15950 6059 15952
rect 6318 16010 6378 16086
rect 6821 16144 11487 16146
rect 6821 16088 6826 16144
rect 6882 16088 11426 16144
rect 11482 16088 11487 16144
rect 6821 16086 11487 16088
rect 6821 16083 6887 16086
rect 11421 16083 11487 16086
rect 10041 16010 10107 16013
rect 6318 16008 10107 16010
rect 6318 15952 10046 16008
rect 10102 15952 10107 16008
rect 6318 15950 10107 15952
rect 0 15874 480 15904
rect 1577 15874 1643 15877
rect 0 15872 1643 15874
rect 0 15816 1582 15872
rect 1638 15816 1643 15872
rect 0 15814 1643 15816
rect 0 15784 480 15814
rect 1577 15811 1643 15814
rect 2865 15874 2931 15877
rect 4429 15874 4495 15877
rect 4662 15874 4722 15950
rect 5993 15947 6059 15950
rect 10041 15947 10107 15950
rect 2865 15872 4722 15874
rect 2865 15816 2870 15872
rect 2926 15816 4434 15872
rect 4490 15816 4722 15872
rect 2865 15814 4722 15816
rect 4889 15874 4955 15877
rect 5717 15874 5783 15877
rect 4889 15872 5783 15874
rect 4889 15816 4894 15872
rect 4950 15816 5722 15872
rect 5778 15816 5783 15872
rect 4889 15814 5783 15816
rect 2865 15811 2931 15814
rect 4429 15811 4495 15814
rect 4889 15811 4955 15814
rect 5717 15811 5783 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 3049 15738 3115 15741
rect 3509 15738 3575 15741
rect 5901 15738 5967 15741
rect 3049 15736 5967 15738
rect 3049 15680 3054 15736
rect 3110 15680 3514 15736
rect 3570 15680 5906 15736
rect 5962 15680 5967 15736
rect 3049 15678 5967 15680
rect 3049 15675 3115 15678
rect 3509 15675 3575 15678
rect 5901 15675 5967 15678
rect 2405 15602 2471 15605
rect 15009 15602 15075 15605
rect 2405 15600 15075 15602
rect 2405 15544 2410 15600
rect 2466 15544 15014 15600
rect 15070 15544 15075 15600
rect 2405 15542 15075 15544
rect 2405 15539 2471 15542
rect 15009 15539 15075 15542
rect 0 15466 480 15496
rect 3417 15466 3483 15469
rect 0 15464 3483 15466
rect 0 15408 3422 15464
rect 3478 15408 3483 15464
rect 0 15406 3483 15408
rect 0 15376 480 15406
rect 3417 15403 3483 15406
rect 4521 15466 4587 15469
rect 8937 15466 9003 15469
rect 4521 15464 9003 15466
rect 4521 15408 4526 15464
rect 4582 15408 8942 15464
rect 8998 15408 9003 15464
rect 4521 15406 9003 15408
rect 4521 15403 4587 15406
rect 8937 15403 9003 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 3693 15058 3759 15061
rect 7281 15058 7347 15061
rect 3693 15056 7347 15058
rect 3693 15000 3698 15056
rect 3754 15000 7286 15056
rect 7342 15000 7347 15056
rect 3693 14998 7347 15000
rect 3693 14995 3759 14998
rect 7281 14995 7347 14998
rect 9949 15058 10015 15061
rect 15377 15058 15443 15061
rect 9949 15056 15443 15058
rect 9949 15000 9954 15056
rect 10010 15000 15382 15056
rect 15438 15000 15443 15056
rect 9949 14998 15443 15000
rect 9949 14995 10015 14998
rect 15377 14995 15443 14998
rect 0 14922 480 14952
rect 1669 14922 1735 14925
rect 0 14920 1735 14922
rect 0 14864 1674 14920
rect 1730 14864 1735 14920
rect 0 14862 1735 14864
rect 0 14832 480 14862
rect 1669 14859 1735 14862
rect 5901 14922 5967 14925
rect 5901 14920 8402 14922
rect 5901 14864 5906 14920
rect 5962 14864 8402 14920
rect 5901 14862 8402 14864
rect 5901 14859 5967 14862
rect 8342 14786 8402 14862
rect 9029 14786 9095 14789
rect 12893 14786 12959 14789
rect 8342 14784 12959 14786
rect 8342 14728 9034 14784
rect 9090 14728 12898 14784
rect 12954 14728 12959 14784
rect 8342 14726 12959 14728
rect 9029 14723 9095 14726
rect 12893 14723 12959 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 0 14514 480 14544
rect 3325 14514 3391 14517
rect 0 14512 3391 14514
rect 0 14456 3330 14512
rect 3386 14456 3391 14512
rect 0 14454 3391 14456
rect 0 14424 480 14454
rect 3325 14451 3391 14454
rect 10961 14514 11027 14517
rect 13537 14514 13603 14517
rect 10961 14512 13603 14514
rect 10961 14456 10966 14512
rect 11022 14456 13542 14512
rect 13598 14456 13603 14512
rect 10961 14454 13603 14456
rect 10961 14451 11027 14454
rect 13537 14451 13603 14454
rect 4245 14378 4311 14381
rect 4797 14378 4863 14381
rect 4245 14376 4863 14378
rect 4245 14320 4250 14376
rect 4306 14320 4802 14376
rect 4858 14320 4863 14376
rect 4245 14318 4863 14320
rect 4245 14315 4311 14318
rect 4797 14315 4863 14318
rect 10961 14378 11027 14381
rect 15745 14378 15811 14381
rect 10961 14376 15811 14378
rect 10961 14320 10966 14376
rect 11022 14320 15750 14376
rect 15806 14320 15811 14376
rect 10961 14318 15811 14320
rect 10961 14315 11027 14318
rect 15745 14315 15811 14318
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 4889 14106 4955 14109
rect 7557 14106 7623 14109
rect 4889 14104 7623 14106
rect 4889 14048 4894 14104
rect 4950 14048 7562 14104
rect 7618 14048 7623 14104
rect 4889 14046 7623 14048
rect 4889 14043 4955 14046
rect 7557 14043 7623 14046
rect 0 13970 480 14000
rect 3969 13970 4035 13973
rect 0 13968 4035 13970
rect 0 13912 3974 13968
rect 4030 13912 4035 13968
rect 0 13910 4035 13912
rect 0 13880 480 13910
rect 3969 13907 4035 13910
rect 9949 13970 10015 13973
rect 15101 13970 15167 13973
rect 9949 13968 15167 13970
rect 9949 13912 9954 13968
rect 10010 13912 15106 13968
rect 15162 13912 15167 13968
rect 9949 13910 15167 13912
rect 9949 13907 10015 13910
rect 15101 13907 15167 13910
rect 5349 13834 5415 13837
rect 8845 13834 8911 13837
rect 5349 13832 8911 13834
rect 5349 13776 5354 13832
rect 5410 13776 8850 13832
rect 8906 13776 8911 13832
rect 5349 13774 8911 13776
rect 5349 13771 5415 13774
rect 8845 13771 8911 13774
rect 10869 13834 10935 13837
rect 11605 13834 11671 13837
rect 16665 13834 16731 13837
rect 10869 13832 16731 13834
rect 10869 13776 10874 13832
rect 10930 13776 11610 13832
rect 11666 13776 16670 13832
rect 16726 13776 16731 13832
rect 10869 13774 16731 13776
rect 10869 13771 10935 13774
rect 11605 13771 11671 13774
rect 16665 13771 16731 13774
rect 7808 13632 8128 13633
rect 0 13562 480 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 4061 13562 4127 13565
rect 0 13560 4127 13562
rect 0 13504 4066 13560
rect 4122 13504 4127 13560
rect 0 13502 4127 13504
rect 0 13472 480 13502
rect 4061 13499 4127 13502
rect 10777 13426 10843 13429
rect 11789 13426 11855 13429
rect 10777 13424 11855 13426
rect 10777 13368 10782 13424
rect 10838 13368 11794 13424
rect 11850 13368 11855 13424
rect 10777 13366 11855 13368
rect 10777 13363 10843 13366
rect 11789 13363 11855 13366
rect 12525 13156 12591 13157
rect 12525 13152 12572 13156
rect 12636 13154 12642 13156
rect 12525 13096 12530 13152
rect 12525 13092 12572 13096
rect 12636 13094 12682 13154
rect 12636 13092 12642 13094
rect 12525 13091 12591 13092
rect 4376 13088 4696 13089
rect 0 13018 480 13048
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 3785 13018 3851 13021
rect 0 13016 3851 13018
rect 0 12960 3790 13016
rect 3846 12960 3851 13016
rect 0 12958 3851 12960
rect 0 12928 480 12958
rect 3785 12955 3851 12958
rect 4245 12746 4311 12749
rect 8477 12746 8543 12749
rect 4245 12744 8543 12746
rect 4245 12688 4250 12744
rect 4306 12688 8482 12744
rect 8538 12688 8543 12744
rect 4245 12686 8543 12688
rect 4245 12683 4311 12686
rect 8477 12683 8543 12686
rect 0 12610 480 12640
rect 3601 12610 3667 12613
rect 0 12608 3667 12610
rect 0 12552 3606 12608
rect 3662 12552 3667 12608
rect 0 12550 3667 12552
rect 0 12520 480 12550
rect 3601 12547 3667 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 2957 12474 3023 12477
rect 7005 12474 7071 12477
rect 7373 12474 7439 12477
rect 2957 12472 7439 12474
rect 2957 12416 2962 12472
rect 3018 12416 7010 12472
rect 7066 12416 7378 12472
rect 7434 12416 7439 12472
rect 2957 12414 7439 12416
rect 2957 12411 3023 12414
rect 7005 12411 7071 12414
rect 7373 12411 7439 12414
rect 11421 12474 11487 12477
rect 11881 12474 11947 12477
rect 14089 12474 14155 12477
rect 11421 12472 11947 12474
rect 11421 12416 11426 12472
rect 11482 12416 11886 12472
rect 11942 12416 11947 12472
rect 11421 12414 11947 12416
rect 11421 12411 11487 12414
rect 11881 12411 11947 12414
rect 12022 12472 14155 12474
rect 12022 12416 14094 12472
rect 14150 12416 14155 12472
rect 12022 12414 14155 12416
rect 3969 12338 4035 12341
rect 9673 12338 9739 12341
rect 12022 12338 12082 12414
rect 14089 12411 14155 12414
rect 3969 12336 9739 12338
rect 3969 12280 3974 12336
rect 4030 12280 9678 12336
rect 9734 12280 9739 12336
rect 3969 12278 9739 12280
rect 3969 12275 4035 12278
rect 9673 12275 9739 12278
rect 11470 12278 12082 12338
rect 13905 12338 13971 12341
rect 14273 12338 14339 12341
rect 13905 12336 14339 12338
rect 13905 12280 13910 12336
rect 13966 12280 14278 12336
rect 14334 12280 14339 12336
rect 13905 12278 14339 12280
rect 7281 12202 7347 12205
rect 11470 12202 11530 12278
rect 13905 12275 13971 12278
rect 14273 12275 14339 12278
rect 4248 12142 7114 12202
rect 0 12066 480 12096
rect 4248 12066 4308 12142
rect 0 12006 4308 12066
rect 7054 12066 7114 12142
rect 7281 12200 11530 12202
rect 7281 12144 7286 12200
rect 7342 12144 11530 12200
rect 7281 12142 11530 12144
rect 11697 12202 11763 12205
rect 12157 12202 12223 12205
rect 11697 12200 12223 12202
rect 11697 12144 11702 12200
rect 11758 12144 12162 12200
rect 12218 12144 12223 12200
rect 11697 12142 12223 12144
rect 7281 12139 7347 12142
rect 11697 12139 11763 12142
rect 12157 12139 12223 12142
rect 9581 12066 9647 12069
rect 7054 12064 9647 12066
rect 7054 12008 9586 12064
rect 9642 12008 9647 12064
rect 7054 12006 9647 12008
rect 0 11976 480 12006
rect 9581 12003 9647 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 4981 11794 5047 11797
rect 5206 11794 5212 11796
rect 4981 11792 5212 11794
rect 4981 11736 4986 11792
rect 5042 11736 5212 11792
rect 4981 11734 5212 11736
rect 4981 11731 5047 11734
rect 5206 11732 5212 11734
rect 5276 11732 5282 11796
rect 12566 11732 12572 11796
rect 12636 11794 12642 11796
rect 12801 11794 12867 11797
rect 14089 11794 14155 11797
rect 14641 11794 14707 11797
rect 12636 11792 14707 11794
rect 12636 11736 12806 11792
rect 12862 11736 14094 11792
rect 14150 11736 14646 11792
rect 14702 11736 14707 11792
rect 12636 11734 14707 11736
rect 12636 11732 12642 11734
rect 12801 11731 12867 11734
rect 14089 11731 14155 11734
rect 14641 11731 14707 11734
rect 0 11658 480 11688
rect 4245 11658 4311 11661
rect 0 11656 4311 11658
rect 0 11600 4250 11656
rect 4306 11600 4311 11656
rect 0 11598 4311 11600
rect 0 11568 480 11598
rect 4245 11595 4311 11598
rect 7649 11658 7715 11661
rect 13905 11658 13971 11661
rect 7649 11656 13971 11658
rect 7649 11600 7654 11656
rect 7710 11600 13910 11656
rect 13966 11600 13971 11656
rect 7649 11598 13971 11600
rect 7649 11595 7715 11598
rect 13905 11595 13971 11598
rect 9949 11522 10015 11525
rect 11881 11522 11947 11525
rect 9949 11520 11947 11522
rect 9949 11464 9954 11520
rect 10010 11464 11886 11520
rect 11942 11464 11947 11520
rect 9949 11462 11947 11464
rect 9949 11459 10015 11462
rect 11881 11459 11947 11462
rect 12525 11522 12591 11525
rect 14365 11522 14431 11525
rect 12525 11520 14431 11522
rect 12525 11464 12530 11520
rect 12586 11464 14370 11520
rect 14426 11464 14431 11520
rect 12525 11462 14431 11464
rect 12525 11459 12591 11462
rect 14365 11459 14431 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 11973 11250 12039 11253
rect 15285 11250 15351 11253
rect 11973 11248 15351 11250
rect 11973 11192 11978 11248
rect 12034 11192 15290 11248
rect 15346 11192 15351 11248
rect 11973 11190 15351 11192
rect 11973 11187 12039 11190
rect 15285 11187 15351 11190
rect 0 11114 480 11144
rect 8661 11114 8727 11117
rect 0 11112 8727 11114
rect 0 11056 8666 11112
rect 8722 11056 8727 11112
rect 0 11054 8727 11056
rect 0 11024 480 11054
rect 8661 11051 8727 11054
rect 10869 11114 10935 11117
rect 14641 11114 14707 11117
rect 10869 11112 14707 11114
rect 10869 11056 10874 11112
rect 10930 11056 14646 11112
rect 14702 11056 14707 11112
rect 10869 11054 14707 11056
rect 10869 11051 10935 11054
rect 14641 11051 14707 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 0 10706 480 10736
rect 1393 10706 1459 10709
rect 0 10704 1459 10706
rect 0 10648 1398 10704
rect 1454 10648 1459 10704
rect 0 10646 1459 10648
rect 0 10616 480 10646
rect 1393 10643 1459 10646
rect 6637 10706 6703 10709
rect 8293 10706 8359 10709
rect 6637 10704 8359 10706
rect 6637 10648 6642 10704
rect 6698 10648 8298 10704
rect 8354 10648 8359 10704
rect 6637 10646 8359 10648
rect 6637 10643 6703 10646
rect 8293 10643 8359 10646
rect 4889 10570 4955 10573
rect 9397 10570 9463 10573
rect 4889 10568 9463 10570
rect 4889 10512 4894 10568
rect 4950 10512 9402 10568
rect 9458 10512 9463 10568
rect 4889 10510 9463 10512
rect 4889 10507 4955 10510
rect 9397 10507 9463 10510
rect 6269 10434 6335 10437
rect 4340 10432 6335 10434
rect 4340 10376 6274 10432
rect 6330 10376 6335 10432
rect 4340 10374 6335 10376
rect 0 10162 480 10192
rect 4340 10162 4400 10374
rect 6269 10371 6335 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 4613 10298 4679 10301
rect 5809 10298 5875 10301
rect 4613 10296 5875 10298
rect 4613 10240 4618 10296
rect 4674 10240 5814 10296
rect 5870 10240 5875 10296
rect 4613 10238 5875 10240
rect 4613 10235 4679 10238
rect 5809 10235 5875 10238
rect 9765 10298 9831 10301
rect 12801 10298 12867 10301
rect 14273 10298 14339 10301
rect 9765 10296 14339 10298
rect 9765 10240 9770 10296
rect 9826 10240 12806 10296
rect 12862 10240 14278 10296
rect 14334 10240 14339 10296
rect 9765 10238 14339 10240
rect 9765 10235 9831 10238
rect 12801 10235 12867 10238
rect 14273 10235 14339 10238
rect 0 10102 4400 10162
rect 4521 10162 4587 10165
rect 8569 10162 8635 10165
rect 9213 10162 9279 10165
rect 4521 10160 9279 10162
rect 4521 10104 4526 10160
rect 4582 10104 8574 10160
rect 8630 10104 9218 10160
rect 9274 10104 9279 10160
rect 4521 10102 9279 10104
rect 0 10072 480 10102
rect 4521 10099 4587 10102
rect 8569 10099 8635 10102
rect 9213 10099 9279 10102
rect 10593 10162 10659 10165
rect 13537 10162 13603 10165
rect 10593 10160 13603 10162
rect 10593 10104 10598 10160
rect 10654 10104 13542 10160
rect 13598 10104 13603 10160
rect 10593 10102 13603 10104
rect 10593 10099 10659 10102
rect 13537 10099 13603 10102
rect 4245 10026 4311 10029
rect 5165 10026 5231 10029
rect 4245 10024 5231 10026
rect 4245 9968 4250 10024
rect 4306 9968 5170 10024
rect 5226 9968 5231 10024
rect 4245 9966 5231 9968
rect 4245 9963 4311 9966
rect 5165 9963 5231 9966
rect 4376 9824 4696 9825
rect 0 9754 480 9784
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 3969 9754 4035 9757
rect 0 9752 4035 9754
rect 0 9696 3974 9752
rect 4030 9696 4035 9752
rect 0 9694 4035 9696
rect 0 9664 480 9694
rect 3969 9691 4035 9694
rect 10869 9618 10935 9621
rect 10869 9616 12818 9618
rect 10869 9560 10874 9616
rect 10930 9560 12818 9616
rect 10869 9558 12818 9560
rect 10869 9555 10935 9558
rect 8477 9482 8543 9485
rect 12617 9482 12683 9485
rect 8477 9480 12683 9482
rect 8477 9424 8482 9480
rect 8538 9424 12622 9480
rect 12678 9424 12683 9480
rect 8477 9422 12683 9424
rect 12758 9482 12818 9558
rect 14038 9556 14044 9620
rect 14108 9618 14114 9620
rect 14181 9618 14247 9621
rect 14108 9616 14247 9618
rect 14108 9560 14186 9616
rect 14242 9560 14247 9616
rect 14108 9558 14247 9560
rect 14108 9556 14114 9558
rect 14181 9555 14247 9558
rect 13905 9482 13971 9485
rect 12758 9480 13971 9482
rect 12758 9424 13910 9480
rect 13966 9424 13971 9480
rect 12758 9422 13971 9424
rect 8477 9419 8543 9422
rect 12617 9419 12683 9422
rect 13905 9419 13971 9422
rect 3785 9346 3851 9349
rect 7281 9346 7347 9349
rect 3785 9344 7347 9346
rect 3785 9288 3790 9344
rect 3846 9288 7286 9344
rect 7342 9288 7347 9344
rect 3785 9286 7347 9288
rect 3785 9283 3851 9286
rect 7281 9283 7347 9286
rect 9489 9346 9555 9349
rect 10133 9346 10199 9349
rect 9489 9344 10199 9346
rect 9489 9288 9494 9344
rect 9550 9288 10138 9344
rect 10194 9288 10199 9344
rect 9489 9286 10199 9288
rect 9489 9283 9555 9286
rect 10133 9283 10199 9286
rect 11605 9346 11671 9349
rect 12433 9346 12499 9349
rect 11605 9344 12499 9346
rect 11605 9288 11610 9344
rect 11666 9288 12438 9344
rect 12494 9288 12499 9344
rect 11605 9286 12499 9288
rect 11605 9283 11671 9286
rect 12433 9283 12499 9286
rect 7808 9280 8128 9281
rect 0 9210 480 9240
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 13077 9210 13143 9213
rect 0 9150 4906 9210
rect 0 9120 480 9150
rect 4846 8938 4906 9150
rect 11286 9208 13143 9210
rect 11286 9152 13082 9208
rect 13138 9152 13143 9208
rect 11286 9150 13143 9152
rect 9581 9074 9647 9077
rect 11286 9074 11346 9150
rect 13077 9147 13143 9150
rect 9581 9072 11346 9074
rect 9581 9016 9586 9072
rect 9642 9016 11346 9072
rect 9581 9014 11346 9016
rect 11421 9074 11487 9077
rect 12341 9074 12407 9077
rect 11421 9072 12407 9074
rect 11421 9016 11426 9072
rect 11482 9016 12346 9072
rect 12402 9016 12407 9072
rect 11421 9014 12407 9016
rect 9581 9011 9647 9014
rect 11421 9011 11487 9014
rect 12341 9011 12407 9014
rect 8661 8938 8727 8941
rect 11145 8940 11211 8941
rect 4846 8936 8727 8938
rect 4846 8880 8666 8936
rect 8722 8880 8727 8936
rect 4846 8878 8727 8880
rect 8661 8875 8727 8878
rect 11094 8876 11100 8940
rect 11164 8938 11211 8940
rect 11881 8938 11947 8941
rect 11164 8936 11947 8938
rect 11206 8880 11886 8936
rect 11942 8880 11947 8936
rect 11164 8878 11947 8880
rect 11164 8876 11211 8878
rect 11145 8875 11211 8876
rect 11881 8875 11947 8878
rect 0 8802 480 8832
rect 3969 8802 4035 8805
rect 0 8800 4035 8802
rect 0 8744 3974 8800
rect 4030 8744 4035 8800
rect 0 8742 4035 8744
rect 0 8712 480 8742
rect 3969 8739 4035 8742
rect 12065 8802 12131 8805
rect 13261 8802 13327 8805
rect 12065 8800 13327 8802
rect 12065 8744 12070 8800
rect 12126 8744 13266 8800
rect 13322 8744 13327 8800
rect 12065 8742 13327 8744
rect 12065 8739 12131 8742
rect 13261 8739 13327 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 7005 8666 7071 8669
rect 9581 8666 9647 8669
rect 7005 8664 9647 8666
rect 7005 8608 7010 8664
rect 7066 8608 9586 8664
rect 9642 8608 9647 8664
rect 7005 8606 9647 8608
rect 7005 8603 7071 8606
rect 9581 8603 9647 8606
rect 10501 8530 10567 8533
rect 15653 8530 15719 8533
rect 10501 8528 15719 8530
rect 10501 8472 10506 8528
rect 10562 8472 15658 8528
rect 15714 8472 15719 8528
rect 10501 8470 15719 8472
rect 10501 8467 10567 8470
rect 15653 8467 15719 8470
rect 8753 8394 8819 8397
rect 12341 8394 12407 8397
rect 8753 8392 12407 8394
rect 8753 8336 8758 8392
rect 8814 8336 12346 8392
rect 12402 8336 12407 8392
rect 8753 8334 12407 8336
rect 8753 8331 8819 8334
rect 12341 8331 12407 8334
rect 0 8258 480 8288
rect 3969 8258 4035 8261
rect 0 8256 4035 8258
rect 0 8200 3974 8256
rect 4030 8200 4035 8256
rect 0 8198 4035 8200
rect 0 8168 480 8198
rect 3969 8195 4035 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 0 7850 480 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 480 7790
rect 4061 7787 4127 7790
rect 11605 7850 11671 7853
rect 13445 7850 13511 7853
rect 11605 7848 13511 7850
rect 11605 7792 11610 7848
rect 11666 7792 13450 7848
rect 13506 7792 13511 7848
rect 11605 7790 13511 7792
rect 11605 7787 11671 7790
rect 13445 7787 13511 7790
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 7925 7442 7991 7445
rect 12893 7442 12959 7445
rect 7925 7440 12959 7442
rect 7925 7384 7930 7440
rect 7986 7384 12898 7440
rect 12954 7384 12959 7440
rect 7925 7382 12959 7384
rect 7925 7379 7991 7382
rect 12893 7379 12959 7382
rect 0 7306 480 7336
rect 2405 7306 2471 7309
rect 0 7304 2471 7306
rect 0 7248 2410 7304
rect 2466 7248 2471 7304
rect 0 7246 2471 7248
rect 0 7216 480 7246
rect 2405 7243 2471 7246
rect 12525 7306 12591 7309
rect 12525 7304 12634 7306
rect 12525 7248 12530 7304
rect 12586 7248 12634 7304
rect 12525 7243 12634 7248
rect 12574 7170 12634 7243
rect 12709 7170 12775 7173
rect 12574 7168 12775 7170
rect 12574 7112 12714 7168
rect 12770 7112 12775 7168
rect 12574 7110 12775 7112
rect 12709 7107 12775 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 12065 7034 12131 7037
rect 12249 7034 12315 7037
rect 12065 7032 12315 7034
rect 12065 6976 12070 7032
rect 12126 6976 12254 7032
rect 12310 6976 12315 7032
rect 12065 6974 12315 6976
rect 12065 6971 12131 6974
rect 12249 6971 12315 6974
rect 0 6898 480 6928
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6808 480 6838
rect 4061 6835 4127 6838
rect 9213 6898 9279 6901
rect 17493 6898 17559 6901
rect 9213 6896 17559 6898
rect 9213 6840 9218 6896
rect 9274 6840 17498 6896
rect 17554 6840 17559 6896
rect 9213 6838 17559 6840
rect 9213 6835 9279 6838
rect 17493 6835 17559 6838
rect 10501 6762 10567 6765
rect 798 6760 10567 6762
rect 798 6704 10506 6760
rect 10562 6704 10567 6760
rect 798 6702 10567 6704
rect 0 6354 480 6384
rect 798 6354 858 6702
rect 10501 6699 10567 6702
rect 11053 6762 11119 6765
rect 14089 6762 14155 6765
rect 11053 6760 14155 6762
rect 11053 6704 11058 6760
rect 11114 6704 14094 6760
rect 14150 6704 14155 6760
rect 11053 6702 14155 6704
rect 11053 6699 11119 6702
rect 14089 6699 14155 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6294 858 6354
rect 10593 6354 10659 6357
rect 13169 6354 13235 6357
rect 10593 6352 13235 6354
rect 10593 6296 10598 6352
rect 10654 6296 13174 6352
rect 13230 6296 13235 6352
rect 10593 6294 13235 6296
rect 0 6264 480 6294
rect 10593 6291 10659 6294
rect 13169 6291 13235 6294
rect 6913 6218 6979 6221
rect 14089 6218 14155 6221
rect 6913 6216 14155 6218
rect 6913 6160 6918 6216
rect 6974 6160 14094 6216
rect 14150 6160 14155 6216
rect 6913 6158 14155 6160
rect 6913 6155 6979 6158
rect 14089 6155 14155 6158
rect 10041 6082 10107 6085
rect 11973 6082 12039 6085
rect 10041 6080 12039 6082
rect 10041 6024 10046 6080
rect 10102 6024 11978 6080
rect 12034 6024 12039 6080
rect 10041 6022 12039 6024
rect 10041 6019 10107 6022
rect 11973 6019 12039 6022
rect 7808 6016 8128 6017
rect 0 5946 480 5976
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 4521 5946 4587 5949
rect 0 5944 4587 5946
rect 0 5888 4526 5944
rect 4582 5888 4587 5944
rect 0 5886 4587 5888
rect 0 5856 480 5886
rect 4521 5883 4587 5886
rect 3141 5810 3207 5813
rect 17953 5810 18019 5813
rect 3141 5808 18019 5810
rect 3141 5752 3146 5808
rect 3202 5752 17958 5808
rect 18014 5752 18019 5808
rect 3141 5750 18019 5752
rect 3141 5747 3207 5750
rect 17953 5747 18019 5750
rect 18689 5810 18755 5813
rect 22320 5810 22800 5840
rect 18689 5808 22800 5810
rect 18689 5752 18694 5808
rect 18750 5752 22800 5808
rect 18689 5750 22800 5752
rect 18689 5747 18755 5750
rect 22320 5720 22800 5750
rect 9857 5674 9923 5677
rect 10409 5674 10475 5677
rect 18873 5674 18939 5677
rect 9857 5672 18939 5674
rect 9857 5616 9862 5672
rect 9918 5616 10414 5672
rect 10470 5616 18878 5672
rect 18934 5616 18939 5672
rect 9857 5614 18939 5616
rect 9857 5611 9923 5614
rect 10409 5611 10475 5614
rect 18873 5611 18939 5614
rect 4376 5472 4696 5473
rect 0 5402 480 5432
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 3969 5402 4035 5405
rect 0 5400 4035 5402
rect 0 5344 3974 5400
rect 4030 5344 4035 5400
rect 0 5342 4035 5344
rect 0 5312 480 5342
rect 3969 5339 4035 5342
rect 10133 5266 10199 5269
rect 14825 5266 14891 5269
rect 10133 5264 14891 5266
rect 10133 5208 10138 5264
rect 10194 5208 14830 5264
rect 14886 5208 14891 5264
rect 10133 5206 14891 5208
rect 10133 5203 10199 5206
rect 14825 5203 14891 5206
rect 0 4994 480 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 0 4904 480 4934
rect 4061 4931 4127 4934
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 7925 4722 7991 4725
rect 4156 4720 7991 4722
rect 4156 4664 7930 4720
rect 7986 4664 7991 4720
rect 4156 4662 7991 4664
rect 0 4450 480 4480
rect 4156 4450 4216 4662
rect 7925 4659 7991 4662
rect 6085 4586 6151 4589
rect 7925 4586 7991 4589
rect 6085 4584 7991 4586
rect 6085 4528 6090 4584
rect 6146 4528 7930 4584
rect 7986 4528 7991 4584
rect 6085 4526 7991 4528
rect 6085 4523 6151 4526
rect 7925 4523 7991 4526
rect 0 4390 4216 4450
rect 0 4360 480 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 10593 4178 10659 4181
rect 14457 4178 14523 4181
rect 10593 4176 14523 4178
rect 10593 4120 10598 4176
rect 10654 4120 14462 4176
rect 14518 4120 14523 4176
rect 10593 4118 14523 4120
rect 10593 4115 10659 4118
rect 14457 4115 14523 4118
rect 0 4042 480 4072
rect 2773 4042 2839 4045
rect 0 4040 2839 4042
rect 0 3984 2778 4040
rect 2834 3984 2839 4040
rect 0 3982 2839 3984
rect 0 3952 480 3982
rect 2773 3979 2839 3982
rect 6729 4042 6795 4045
rect 14038 4042 14044 4044
rect 6729 4040 14044 4042
rect 6729 3984 6734 4040
rect 6790 3984 14044 4040
rect 6729 3982 14044 3984
rect 6729 3979 6795 3982
rect 14038 3980 14044 3982
rect 14108 3980 14114 4044
rect 3141 3906 3207 3909
rect 7097 3906 7163 3909
rect 3141 3904 7163 3906
rect 3141 3848 3146 3904
rect 3202 3848 7102 3904
rect 7158 3848 7163 3904
rect 3141 3846 7163 3848
rect 3141 3843 3207 3846
rect 7097 3843 7163 3846
rect 8661 3906 8727 3909
rect 11094 3906 11100 3908
rect 8661 3904 11100 3906
rect 8661 3848 8666 3904
rect 8722 3848 11100 3904
rect 8661 3846 11100 3848
rect 8661 3843 8727 3846
rect 11094 3844 11100 3846
rect 11164 3844 11170 3908
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 6177 3634 6243 3637
rect 15469 3634 15535 3637
rect 6177 3632 15535 3634
rect 6177 3576 6182 3632
rect 6238 3576 15474 3632
rect 15530 3576 15535 3632
rect 6177 3574 15535 3576
rect 6177 3571 6243 3574
rect 15469 3571 15535 3574
rect 0 3498 480 3528
rect 4889 3498 4955 3501
rect 5165 3498 5231 3501
rect 0 3496 5231 3498
rect 0 3440 4894 3496
rect 4950 3440 5170 3496
rect 5226 3440 5231 3496
rect 0 3438 5231 3440
rect 0 3408 480 3438
rect 4889 3435 4955 3438
rect 5165 3435 5231 3438
rect 9765 3498 9831 3501
rect 10869 3498 10935 3501
rect 11421 3498 11487 3501
rect 9765 3496 11487 3498
rect 9765 3440 9770 3496
rect 9826 3440 10874 3496
rect 10930 3440 11426 3496
rect 11482 3440 11487 3496
rect 9765 3438 11487 3440
rect 9765 3435 9831 3438
rect 10869 3435 10935 3438
rect 11421 3435 11487 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 3090 480 3120
rect 2957 3090 3023 3093
rect 0 3088 3023 3090
rect 0 3032 2962 3088
rect 3018 3032 3023 3088
rect 0 3030 3023 3032
rect 0 3000 480 3030
rect 2957 3027 3023 3030
rect 7281 3090 7347 3093
rect 9213 3090 9279 3093
rect 7281 3088 9279 3090
rect 7281 3032 7286 3088
rect 7342 3032 9218 3088
rect 9274 3032 9279 3088
rect 7281 3030 9279 3032
rect 7281 3027 7347 3030
rect 9213 3027 9279 3030
rect 5809 2954 5875 2957
rect 10317 2954 10383 2957
rect 14733 2954 14799 2957
rect 5809 2952 14799 2954
rect 5809 2896 5814 2952
rect 5870 2896 10322 2952
rect 10378 2896 14738 2952
rect 14794 2896 14799 2952
rect 5809 2894 14799 2896
rect 5809 2891 5875 2894
rect 10317 2891 10383 2894
rect 14733 2891 14799 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 480 2486
rect 4061 2483 4127 2486
rect 5441 2546 5507 2549
rect 8109 2546 8175 2549
rect 5441 2544 8175 2546
rect 5441 2488 5446 2544
rect 5502 2488 8114 2544
rect 8170 2488 8175 2544
rect 5441 2486 8175 2488
rect 5441 2483 5507 2486
rect 8109 2483 8175 2486
rect 4376 2208 4696 2209
rect 0 2138 480 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 3049 2138 3115 2141
rect 0 2136 3115 2138
rect 0 2080 3054 2136
rect 3110 2080 3115 2136
rect 0 2078 3115 2080
rect 0 2048 480 2078
rect 3049 2075 3115 2078
rect 0 1594 480 1624
rect 3325 1594 3391 1597
rect 0 1592 3391 1594
rect 0 1536 3330 1592
rect 3386 1536 3391 1592
rect 0 1534 3391 1536
rect 0 1504 480 1534
rect 3325 1531 3391 1534
rect 0 1186 480 1216
rect 2773 1186 2839 1189
rect 0 1184 2839 1186
rect 0 1128 2778 1184
rect 2834 1128 2839 1184
rect 0 1126 2839 1128
rect 0 1096 480 1126
rect 2773 1123 2839 1126
rect 0 642 480 672
rect 5533 642 5599 645
rect 0 640 5599 642
rect 0 584 5538 640
rect 5594 584 5599 640
rect 0 582 5599 584
rect 0 552 480 582
rect 5533 579 5599 582
rect 0 234 480 264
rect 4153 234 4219 237
rect 0 232 4219 234
rect 0 176 4158 232
rect 4214 176 4219 232
rect 0 174 4219 176
rect 0 144 480 174
rect 4153 171 4219 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 5212 16960 5276 16964
rect 5212 16904 5262 16960
rect 5262 16904 5276 16960
rect 5212 16900 5276 16904
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 12572 13152 12636 13156
rect 12572 13096 12586 13152
rect 12586 13096 12636 13152
rect 12572 13092 12636 13096
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 5212 11732 5276 11796
rect 12572 11732 12636 11796
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 14044 9556 14108 9620
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 11100 8936 11164 8940
rect 11100 8880 11150 8936
rect 11150 8880 11164 8936
rect 11100 8876 11164 8880
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 14044 3980 14108 4044
rect 11100 3844 11164 3908
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 5211 16964 5277 16965
rect 5211 16900 5212 16964
rect 5276 16900 5277 16964
rect 5211 16899 5277 16900
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 5214 11797 5274 16899
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 5211 11796 5277 11797
rect 5211 11732 5212 11796
rect 5276 11732 5277 11796
rect 5211 11731 5277 11732
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 12571 13156 12637 13157
rect 12571 13092 12572 13156
rect 12636 13092 12637 13156
rect 12571 13091 12637 13092
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 12574 11797 12634 13091
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 12571 11796 12637 11797
rect 12571 11732 12572 11796
rect 12636 11732 12637 11796
rect 12571 11731 12637 11732
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11099 8940 11165 8941
rect 11099 8876 11100 8940
rect 11164 8876 11165 8940
rect 11099 8875 11165 8876
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 11102 3909 11162 8875
rect 11240 8736 11560 9760
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14043 9620 14109 9621
rect 14043 9556 14044 9620
rect 14108 9556 14109 9620
rect 14043 9555 14109 9556
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11099 3908 11165 3909
rect 11099 3844 11100 3908
rect 11164 3844 11165 3908
rect 11099 3843 11165 3844
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 3296 11560 4320
rect 14046 4045 14106 9555
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14043 4044 14109 4045
rect 14043 3980 14044 4044
rect 14108 3980 14109 4044
rect 14043 3979 14109 3980
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2300 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1606256979
transform 1 0 2208 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 3680 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21
timestamp 1606256979
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606256979
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 4876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_22 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3128 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1606256979
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1606256979
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45
timestamp 1606256979
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5336 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606256979
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1606256979
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55
timestamp 1606256979
transform 1 0 6164 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1606256979
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8188 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606256979
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1606256979
transform 1 0 7544 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606256979
transform 1 0 8648 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1606256979
transform 1 0 7452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_79
timestamp 1606256979
transform 1 0 8372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1606256979
transform 1 0 7820 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9844 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1606256979
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606256979
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_93
timestamp 1606256979
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1606256979
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1606256979
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10764 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10856 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1606256979
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1606256979
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1606256979
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _090_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 11776 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606256979
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606256979
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606256979
transform 1 0 13984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13432 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1606256979
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1606256979
transform 1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_144
timestamp 1606256979
transform 1 0 14352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1606256979
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1606256979
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1606256979
transform 1 0 15088 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1606256979
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1606256979
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606256979
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606256979
transform 1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1606256979
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606256979
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606256979
transform 1 0 15272 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp 1606256979
transform 1 0 16008 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1606256979
transform 1 0 16008 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606256979
transform 1 0 16100 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_177
timestamp 1606256979
transform 1 0 17388 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_167
timestamp 1606256979
transform 1 0 16468 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_172
timestamp 1606256979
transform 1 0 16928 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606256979
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606256979
transform 1 0 17020 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1606256979
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1606256979
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606256979
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606256979
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606256979
transform 1 0 18860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606256979
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 1606256979
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_197
timestamp 1606256979
transform 1 0 19228 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606256979
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606256979
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_209
timestamp 1606256979
transform 1 0 20332 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_217
timestamp 1606256979
transform 1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1748 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4140 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1606256979
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1606256979
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1606256979
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1606256979
transform 1 0 5796 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1606256979
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1606256979
transform 1 0 6624 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6992 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8648 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_80
timestamp 1606256979
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 9752 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1606256979
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1606256979
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11408 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_110
timestamp 1606256979
transform 1 0 11224 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13064 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14076 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1606256979
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_139
timestamp 1606256979
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606256979
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_147
timestamp 1606256979
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_160
timestamp 1606256979
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606256979
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606256979
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606256979
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606256979
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606256979
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606256979
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1748 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3404 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_23
timestamp 1606256979
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_41
timestamp 1606256979
transform 1 0 4876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606256979
transform 1 0 5152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5612 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1606256979
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_58
timestamp 1606256979
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_62
timestamp 1606256979
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1606256979
transform 1 0 7084 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1606256979
transform 1 0 8096 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1606256979
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606256979
transform 1 0 10396 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_85
timestamp 1606256979
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_98
timestamp 1606256979
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10948 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1606256979
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116
timestamp 1606256979
transform 1 0 11776 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1606256979
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606256979
transform 1 0 15088 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_150
timestamp 1606256979
transform 1 0 14904 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1606256979
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_168
timestamp 1606256979
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1606256979
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606256979
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606256979
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606256979
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1840 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1606256979
transform 1 0 1748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_17
timestamp 1606256979
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4140 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1606256979
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1606256979
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6256 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_49
timestamp 1606256979
transform 1 0 5612 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1606256979
transform 1 0 6164 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8372 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp 1606256979
transform 1 0 7084 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1606256979
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1606256979
transform 1 0 10672 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 1606256979
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1606256979
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11224 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_4_107
timestamp 1606256979
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1606256979
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_137
timestamp 1606256979
transform 1 0 13708 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1606256979
transform 1 0 14076 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1606256979
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1606256979
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606256979
transform 1 0 17848 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 17020 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_171
timestamp 1606256979
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_179
timestamp 1606256979
transform 1 0 17572 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_186
timestamp 1606256979
transform 1 0 18216 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_198
timestamp 1606256979
transform 1 0 19320 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1606256979
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2024 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1606256979
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4600 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3680 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1606256979
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_34
timestamp 1606256979
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_54
timestamp 1606256979
transform 1 0 6072 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1606256979
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8464 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1606256979
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_89
timestamp 1606256979
transform 1 0 9292 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_104
timestamp 1606256979
transform 1 0 10672 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1606256979
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606256979
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1606256979
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606256979
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13340 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606256979
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1606256979
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1606256979
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15364 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_153
timestamp 1606256979
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1606256979
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1606256979
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606256979
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606256979
transform 1 0 19780 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_196
timestamp 1606256979
transform 1 0 19136 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_202
timestamp 1606256979
transform 1 0 19688 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1606256979
transform 1 0 20148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606256979
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1564 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2576 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_14
timestamp 1606256979
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4784 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3220 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_25
timestamp 1606256979
transform 1 0 3404 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1606256979
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1606256979
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_32
timestamp 1606256979
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5244 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606256979
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1606256979
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1606256979
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606256979
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7912 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7360 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_7_71
timestamp 1606256979
transform 1 0 7636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1606256979
transform 1 0 10488 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1606256979
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_93
timestamp 1606256979
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1606256979
transform 1 0 10396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_90
timestamp 1606256979
transform 1 0 9384 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1606256979
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 11500 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1606256979
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1606256979
transform 1 0 11316 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1606256979
transform 1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1606256979
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606256979
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606256979
transform 1 0 13432 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 14168 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_6_129
timestamp 1606256979
transform 1 0 12972 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1606256979
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1606256979
transform 1 0 13708 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp 1606256979
transform 1 0 14076 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 15824 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1606256979
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1606256979
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1606256979
transform 1 0 16928 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1606256979
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_181
timestamp 1606256979
transform 1 0 17756 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1606256979
transform 1 0 16652 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606256979
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606256979
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18860 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1606256979
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1606256979
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606256979
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1606256979
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1656 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606256979
transform 1 0 3312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4048 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_22
timestamp 1606256979
transform 1 0 3128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5888 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1606256979
transform 1 0 5520 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8556 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1606256979
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1606256979
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1606256979
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11684 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1606256979
transform 1 0 11132 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_131
timestamp 1606256979
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_142
timestamp 1606256979
transform 1 0 14168 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606256979
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1606256979
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606256979
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1606256979
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_175
timestamp 1606256979
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_187
timestamp 1606256979
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_199
timestamp 1606256979
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1606256979
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1606256979
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1606256979
transform 1 0 2944 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1606256979
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606256979
transform 1 0 4140 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 4600 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1606256979
transform 1 0 3772 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1606256979
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1606256979
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606256979
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7820 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1606256979
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_82
timestamp 1606256979
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606256979
transform 1 0 8832 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9568 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10580 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_87
timestamp 1606256979
transform 1 0 9108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_91
timestamp 1606256979
transform 1 0 9476 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1606256979
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_106
timestamp 1606256979
transform 1 0 10856 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_110
timestamp 1606256979
transform 1 0 11224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1606256979
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13432 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1606256979
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_143
timestamp 1606256979
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1606256979
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_166
timestamp 1606256979
transform 1 0 16376 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1606256979
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606256979
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606256979
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1606256979
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1606256979
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1606256979
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1606256979
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1606256979
transform 1 0 4232 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606256979
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1606256979
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5428 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_43
timestamp 1606256979
transform 1 0 5060 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7452 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8464 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1606256979
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp 1606256979
transform 1 0 8280 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1606256979
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606256979
transform 1 0 11316 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 11776 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1606256979
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_114
timestamp 1606256979
transform 1 0 11592 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13432 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1606256979
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1606256979
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606256979
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1606256979
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1606256979
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1606256979
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1606256979
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1606256979
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1606256979
transform 1 0 4048 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606256979
transform 1 0 3036 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1606256979
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1606256979
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5060 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606256979
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1606256979
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7084 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8740 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1606256979
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10672 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1606256979
transform 1 0 10212 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1606256979
transform 1 0 10580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606256979
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14444 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_143
timestamp 1606256979
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1606256979
transform 1 0 15272 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1606256979
transform 1 0 16376 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1606256979
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1606256979
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606256979
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606256979
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606256979
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606256979
transform 1 0 1564 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2024 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_8
timestamp 1606256979
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1606256979
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1606256979
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5152 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1606256979
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7820 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1606256979
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1606256979
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606256979
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1606256979
transform 1 0 10672 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1606256979
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1606256979
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1606256979
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1606256979
transform 1 0 11684 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_113
timestamp 1606256979
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp 1606256979
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12696 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1606256979
transform 1 0 13708 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_135
timestamp 1606256979
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1606256979
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1606256979
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606256979
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606256979
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606256979
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606256979
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606256979
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1932 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1606256979
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_18
timestamp 1606256979
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606256979
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1606256979
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_40
timestamp 1606256979
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1606256979
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1606256979
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp 1606256979
transform 1 0 5888 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1606256979
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1606256979
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1606256979
transform 1 0 4968 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1606256979
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_56
timestamp 1606256979
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606256979
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6348 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8096 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8188 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 7820 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606256979
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_73
timestamp 1606256979
transform 1 0 7820 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1606256979
transform 1 0 9568 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1606256979
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_85
timestamp 1606256979
transform 1 0 8924 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_91
timestamp 1606256979
transform 1 0 9476 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1606256979
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1606256979
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606256979
transform 1 0 11592 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11408 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1606256979
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_117
timestamp 1606256979
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1606256979
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_109
timestamp 1606256979
transform 1 0 11132 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14444 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1606256979
transform 1 0 13064 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1606256979
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1606256979
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp 1606256979
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1606256979
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1606256979
transform 1 0 15272 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1606256979
transform 1 0 16376 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606256979
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1606256979
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1606256979
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1606256979
transform 1 0 17480 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1606256979
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606256979
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1606256979
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606256979
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606256979
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1606256979
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1606256979
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2024 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1606256979
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606256979
transform 1 0 3956 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4416 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_26
timestamp 1606256979
transform 1 0 3496 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_30
timestamp 1606256979
transform 1 0 3864 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1606256979
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1606256979
transform 1 0 5888 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1606256979
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606256979
transform 1 0 7084 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7544 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_68
timestamp 1606256979
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10580 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1606256979
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1606256979
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1606256979
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1606256979
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1606256979
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1606256979
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606256979
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_152
timestamp 1606256979
transform 1 0 15088 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_164
timestamp 1606256979
transform 1 0 16192 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_176
timestamp 1606256979
transform 1 0 17296 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1606256979
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1606256979
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1606256979
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1606256979
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1606256979
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606256979
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 4784 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3036 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1606256979
transform 1 0 4324 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1606256979
transform 1 0 4692 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1606256979
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_71
timestamp 1606256979
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606256979
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11132 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11960 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12788 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14076 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1606256979
transform 1 0 13616 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_140
timestamp 1606256979
transform 1 0 13984 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_150
timestamp 1606256979
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1606256979
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1606256979
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1606256979
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1606256979
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1606256979
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2300 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1564 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1606256979
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606256979
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 1606256979
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1606256979
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606256979
transform 1 0 5980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1606256979
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1606256979
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1606256979
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1606256979
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7360 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 8372 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1606256979
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_99
timestamp 1606256979
transform 1 0 10212 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10856 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 1606256979
transform 1 0 10764 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1606256979
transform 1 0 11684 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606256979
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1606256979
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1606256979
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_150
timestamp 1606256979
transform 1 0 14904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1606256979
transform 1 0 16008 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16652 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_168
timestamp 1606256979
transform 1 0 16560 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1606256979
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1606256979
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1606256979
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1606256979
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606256979
transform 1 0 2760 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1748 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1606256979
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_41
timestamp 1606256979
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606256979
transform 1 0 5060 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5888 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1606256979
transform 1 0 5428 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_51
timestamp 1606256979
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1606256979
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1606256979
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1606256979
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606256979
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10212 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1606256979
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_96
timestamp 1606256979
transform 1 0 9936 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11868 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1606256979
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606256979
transform 1 0 13064 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1606256979
transform 1 0 12696 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1606256979
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1606256979
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1606256979
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1606256979
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1606256979
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1606256979
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1606256979
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606256979
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606256979
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1606256979
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606256979
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1606256979
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1606256979
transform 1 0 2116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1606256979
transform 1 0 2760 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_20
timestamp 1606256979
transform 1 0 2944 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606256979
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1606256979
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1606256979
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606256979
transform 1 0 3772 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606256979
transform 1 0 3128 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1606256979
transform 1 0 4508 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1606256979
transform 1 0 4140 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4600 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 5704 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_54
timestamp 1606256979
transform 1 0 6072 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1606256979
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1606256979
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7820 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1606256979
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1606256979
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1606256979
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1606256979
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_89
timestamp 1606256979
transform 1 0 9292 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1606256979
transform 1 0 9660 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1606256979
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1606256979
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 9844 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10580 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 10672 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606256979
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11592 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606256979
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1606256979
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_123
timestamp 1606256979
transform 1 0 12420 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 12880 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1606256979
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1606256979
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_127
timestamp 1606256979
transform 1 0 12788 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1606256979
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606256979
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1606256979
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1606256979
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606256979
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1606256979
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606256979
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1606256979
transform 1 0 15548 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1606256979
transform 1 0 16284 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_166
timestamp 1606256979
transform 1 0 16376 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1606256979
transform 1 0 17480 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1606256979
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_174
timestamp 1606256979
transform 1 0 17112 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_186
timestamp 1606256979
transform 1 0 18216 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1606256979
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1606256979
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_198
timestamp 1606256979
transform 1 0 19320 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1606256979
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 2484 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1606256979
transform 1 0 1472 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_13
timestamp 1606256979
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1606256979
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1606256979
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1606256979
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1606256979
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1606256979
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1606256979
transform 1 0 7820 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1606256979
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1606256979
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606256979
transform 1 0 10304 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1606256979
transform 1 0 9292 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 8832 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_87
timestamp 1606256979
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_98
timestamp 1606256979
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_103
timestamp 1606256979
transform 1 0 10580 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10948 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 11960 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_116
timestamp 1606256979
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1606256979
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_139
timestamp 1606256979
transform 1 0 13892 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14628 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_163
timestamp 1606256979
transform 1 0 16100 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1606256979
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606256979
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1606256979
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1606256979
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606256979
transform 1 0 1472 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 2024 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_8
timestamp 1606256979
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1606256979
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1606256979
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1606256979
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 5060 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6072 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1606256979
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 8188 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1606256979
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_63
timestamp 1606256979
transform 1 0 6900 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1606256979
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1606256979
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 10672 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_86
timestamp 1606256979
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1606256979
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11132 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1606256979
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1606256979
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12788 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_22_143
timestamp 1606256979
transform 1 0 14260 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1606256979
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606256979
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1606256979
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1606256979
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_187
timestamp 1606256979
transform 1 0 18308 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1606256979
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1606256979
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606256979
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606256979
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1472 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1606256979
transform 1 0 2208 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1606256979
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606256979
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1606256979
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1606256979
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1606256979
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_48
timestamp 1606256979
transform 1 0 5520 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606256979
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 8464 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1606256979
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_83
timestamp 1606256979
transform 1 0 8740 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10304 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1606256979
transform 1 0 9108 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_96
timestamp 1606256979
transform 1 0 9936 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1606256979
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1606256979
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12788 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606256979
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1606256979
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 14996 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1606256979
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_160
timestamp 1606256979
transform 1 0 15824 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1606256979
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1606256979
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606256979
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1606256979
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1606256979
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606256979
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1606256979
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1606256979
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606256979
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1606256979
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606256979
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5060 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6716 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1606256979
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1606256979
transform 1 0 6348 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 7912 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_70
timestamp 1606256979
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606256979
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606256979
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12604 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1606256979
transform 1 0 11592 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_109
timestamp 1606256979
transform 1 0 11132 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_113
timestamp 1606256979
transform 1 0 11500 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1606256979
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606256979
transform 1 0 14260 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1606256979
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1606256979
transform 1 0 14536 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1606256979
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606256979
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606256979
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606256979
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606256979
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1606256979
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606256979
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 2944 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1606256979
transform 1 0 1932 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1606256979
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1606256979
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3956 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1606256979
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_40
timestamp 1606256979
transform 1 0 4784 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606256979
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606256979
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1606256979
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606256979
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_71
timestamp 1606256979
transform 1 0 7636 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_83
timestamp 1606256979
transform 1 0 8740 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9016 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1606256979
transform 1 0 10028 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1606256979
transform 1 0 9844 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1606256979
transform 1 0 12512 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1606256979
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1606256979
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606256979
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_123
timestamp 1606256979
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13524 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1606256979
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_141
timestamp 1606256979
transform 1 0 14076 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_153
timestamp 1606256979
transform 1 0 15180 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_165
timestamp 1606256979
transform 1 0 16284 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_177
timestamp 1606256979
transform 1 0 17388 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606256979
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1606256979
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1606256979
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606256979
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606256979
transform 1 0 1656 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606256979
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_17
timestamp 1606256979
transform 1 0 2668 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1606256979
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_10
timestamp 1606256979
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606256979
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4600 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3220 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1606256979
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1606256979
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1606256979
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606256979
transform 1 0 5888 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6256 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_54
timestamp 1606256979
transform 1 0 6072 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1606256979
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_56
timestamp 1606256979
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8096 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_72
timestamp 1606256979
transform 1 0 7728 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_78
timestamp 1606256979
transform 1 0 8280 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606256979
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10304 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1606256979
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606256979
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1606256979
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1606256979
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1606256979
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1606256979
transform 1 0 10948 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1606256979
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1606256979
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_121
timestamp 1606256979
transform 1 0 12236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_116
timestamp 1606256979
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606256979
transform 1 0 11960 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606256979
transform 1 0 11960 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12604 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606256979
transform 1 0 13984 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1606256979
transform 1 0 13432 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14260 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1606256979
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1606256979
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1606256979
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_144
timestamp 1606256979
transform 1 0 14352 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1606256979
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1606256979
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1606256979
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606256979
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1606256979
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1606256979
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606256979
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606256979
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1606256979
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606256979
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1606256979
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606256979
transform 1 0 2944 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 1472 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606256979
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1606256979
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606256979
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_24
timestamp 1606256979
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1606256979
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606256979
transform 1 0 5704 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1606256979
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp 1606256979
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1606256979
transform 1 0 6072 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7452 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1606256979
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606256979
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1606256979
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1606256979
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606256979
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_102
timestamp 1606256979
transform 1 0 10488 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10856 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12512 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1606256979
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606256979
transform 1 0 14260 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_140
timestamp 1606256979
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_147
timestamp 1606256979
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1606256979
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1606256979
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1606256979
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1606256979
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1606256979
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606256979
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606256979
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606256979
transform 1 0 1472 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2024 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2760 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1606256979
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_16
timestamp 1606256979
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3496 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_24
timestamp 1606256979
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606256979
transform 1 0 6164 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_42
timestamp 1606256979
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1606256979
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606256979
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1606256979
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_71
timestamp 1606256979
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1606256979
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_97
timestamp 1606256979
transform 1 0 10028 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606256979
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10856 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_105
timestamp 1606256979
transform 1 0 10764 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1606256979
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606256979
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606256979
transform 1 0 14444 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606256979
transform 1 0 13432 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1606256979
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1606256979
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1606256979
transform 1 0 14812 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_161
timestamp 1606256979
transform 1 0 15916 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1606256979
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606256979
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606256979
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606256979
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1606256979
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606256979
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606256979
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1606256979
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1606256979
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606256979
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_41
timestamp 1606256979
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606256979
transform 1 0 6808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5152 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_60
timestamp 1606256979
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7268 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_65
timestamp 1606256979
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_83
timestamp 1606256979
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606256979
transform 1 0 8924 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1606256979
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606256979
transform 1 0 11316 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11868 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp 1606256979
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1606256979
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13524 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 14260 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1606256979
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1606256979
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1606256979
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_160
timestamp 1606256979
transform 1 0 15824 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_172
timestamp 1606256979
transform 1 0 16928 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1606256979
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18400 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_194
timestamp 1606256979
transform 1 0 18952 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1606256979
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606256979
transform 1 0 1564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 2944 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2116 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1606256979
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_17
timestamp 1606256979
transform 1 0 2668 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606256979
transform 1 0 4600 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1606256979
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1606256979
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606256979
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1606256979
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7360 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1606256979
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606256979
transform 1 0 9016 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9476 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_84
timestamp 1606256979
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1606256979
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606256979
transform 1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1606256979
transform 1 0 10948 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1606256979
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1606256979
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606256979
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_145
timestamp 1606256979
transform 1 0 14444 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1606256979
transform 1 0 16008 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 14720 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_160
timestamp 1606256979
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1606256979
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606256979
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606256979
transform 1 0 17112 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606256979
transform 1 0 16560 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1606256979
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1606256979
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1606256979
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606256979
transform 1 0 19320 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606256979
transform 1 0 18584 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1606256979
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_194
timestamp 1606256979
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_202
timestamp 1606256979
transform 1 0 19688 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_214
timestamp 1606256979
transform 1 0 20792 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606256979
transform 1 0 1656 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 2208 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1606256979
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_18
timestamp 1606256979
transform 1 0 2760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3036 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606256979
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_41
timestamp 1606256979
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5152 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1606256979
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7820 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 7084 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1606256979
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1606256979
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606256979
transform 1 0 9752 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1606256979
transform 1 0 10212 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 8832 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_90
timestamp 1606256979
transform 1 0 9384 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1606256979
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606256979
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1606256979
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11224 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_108
timestamp 1606256979
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_116
timestamp 1606256979
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606256979
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1606256979
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1606256979
transform 1 0 13156 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_129
timestamp 1606256979
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_135
timestamp 1606256979
transform 1 0 13524 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1606256979
transform 1 0 14076 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1606256979
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1606256979
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1606256979
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_146
timestamp 1606256979
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_152
timestamp 1606256979
transform 1 0 15088 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1606256979
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_166
timestamp 1606256979
transform 1 0 16376 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606256979
transform 1 0 17112 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_178
timestamp 1606256979
transform 1 0 17480 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606256979
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606256979
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1606256979
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2962 0 3018 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 22466 0 22522 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 ccff_head
port 9 nsew default input
rlabel metal3 s 22320 17144 22800 17264 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 17866 0 17922 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 20166 0 20222 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 21086 0 21142 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 14094 0 14150 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 15014 0 15070 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 15566 0 15622 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 3790 22320 3846 22800 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 8390 22320 8446 22800 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 8850 22320 8906 22800 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 9310 22320 9366 22800 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 9770 22320 9826 22800 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 10230 22320 10286 22800 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 10690 22320 10746 22800 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 12438 22320 12494 22800 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 4250 22320 4306 22800 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 4710 22320 4766 22800 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 5170 22320 5226 22800 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 5630 22320 5686 22800 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 6090 22320 6146 22800 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 6550 22320 6606 22800 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 7010 22320 7066 22800 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 7470 22320 7526 22800 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 7930 22320 7986 22800 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 12898 22320 12954 22800 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 17958 22320 18014 22800 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 18418 22320 18474 22800 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 18878 22320 18934 22800 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 19338 22320 19394 22800 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 19798 22320 19854 22800 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 20258 22320 20314 22800 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 20718 22320 20774 22800 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 21178 22320 21234 22800 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 21638 22320 21694 22800 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 13358 22320 13414 22800 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 13818 22320 13874 22800 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 14278 22320 14334 22800 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 14738 22320 14794 22800 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 15198 22320 15254 22800 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 15658 22320 15714 22800 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 16118 22320 16174 22800 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 16578 22320 16634 22800 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 17038 22320 17094 22800 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 131 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 132 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_36_
port 133 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 134 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_38_
port 135 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 136 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_40_
port 137 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 138 nsew default input
rlabel metal2 s 22098 22320 22154 22800 6 prog_clk_0_N_in
port 139 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 140 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_43_
port 141 nsew default input
rlabel metal2 s 1030 22320 1086 22800 6 top_left_grid_pin_44_
port 142 nsew default input
rlabel metal2 s 1490 22320 1546 22800 6 top_left_grid_pin_45_
port 143 nsew default input
rlabel metal2 s 1950 22320 2006 22800 6 top_left_grid_pin_46_
port 144 nsew default input
rlabel metal2 s 2410 22320 2466 22800 6 top_left_grid_pin_47_
port 145 nsew default input
rlabel metal2 s 2870 22320 2926 22800 6 top_left_grid_pin_48_
port 146 nsew default input
rlabel metal2 s 3330 22320 3386 22800 6 top_left_grid_pin_49_
port 147 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 149 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
