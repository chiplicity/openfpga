magic
tech EFS8A
magscale 1 2
timestamp 1602269422
<< locali >>
rect 6595 19873 6630 19907
rect 8493 19873 8654 19907
rect 8493 19771 8527 19873
rect 1903 18785 2030 18819
rect 1443 18173 1478 18207
rect 2547 17697 2582 17731
rect 11483 17289 11621 17323
rect 10051 16745 10057 16779
rect 17043 16745 17049 16779
rect 10051 16677 10085 16745
rect 17043 16677 17077 16745
rect 22511 16609 22546 16643
rect 4807 15895 4841 15963
rect 14289 15895 14323 16201
rect 4807 15861 4813 15895
rect 7015 15657 7021 15691
rect 19435 15657 19441 15691
rect 7015 15589 7049 15657
rect 19435 15589 19469 15657
rect 8619 15521 8654 15555
rect 5583 14909 5618 14943
rect 16899 13345 16934 13379
rect 19809 12631 19843 12801
rect 17411 12393 17417 12427
rect 17411 12325 17445 12393
rect 9413 11747 9447 11849
rect 23949 10455 23983 10557
rect 6101 9911 6135 10081
rect 10609 9367 10643 9605
rect 13093 9503 13127 9673
rect 16491 9367 16525 9435
rect 16491 9333 16497 9367
rect 13363 9129 13369 9163
rect 13363 9061 13397 9129
rect 25087 8993 25122 9027
rect 11483 7225 11621 7259
rect 19291 6885 19336 6919
rect 15611 6817 15646 6851
rect 10517 6239 10551 6341
rect 19073 6103 19107 6341
rect 19441 6171 19475 6341
rect 21373 6205 21465 6239
rect 15439 4777 15577 4811
rect 1443 4641 1478 4675
rect 15243 4641 15370 4675
rect 21051 3689 21097 3723
rect 15243 3553 15370 3587
rect 18705 3553 18866 3587
rect 20855 3553 20982 3587
rect 18705 3383 18739 3553
<< viali >>
rect 21256 24225 21290 24259
rect 21327 24021 21361 24055
rect 8769 23817 8803 23851
rect 12633 23817 12667 23851
rect 13737 23817 13771 23851
rect 19349 23817 19383 23851
rect 21557 23817 21591 23851
rect 22569 23817 22603 23851
rect 21281 23749 21315 23783
rect 1869 23681 1903 23715
rect 1476 23613 1510 23647
rect 8585 23613 8619 23647
rect 9137 23613 9171 23647
rect 12449 23613 12483 23647
rect 13001 23613 13035 23647
rect 13553 23613 13587 23647
rect 14105 23613 14139 23647
rect 19165 23613 19199 23647
rect 19717 23613 19751 23647
rect 20637 23613 20671 23647
rect 22068 23613 22102 23647
rect 22155 23545 22189 23579
rect 1547 23477 1581 23511
rect 20821 23477 20855 23511
rect 1593 23273 1627 23307
rect 1409 23137 1443 23171
rect 12909 22729 12943 22763
rect 13369 22729 13403 22763
rect 1685 22593 1719 22627
rect 12725 22525 12759 22559
rect 18128 22525 18162 22559
rect 18199 22389 18233 22423
rect 18613 22389 18647 22423
rect 6904 20349 6938 20383
rect 6975 20213 7009 20247
rect 7389 20213 7423 20247
rect 12403 20009 12437 20043
rect 6561 19873 6595 19907
rect 12332 19873 12366 19907
rect 12725 19873 12759 19907
rect 8493 19737 8527 19771
rect 6699 19669 6733 19703
rect 8723 19669 8757 19703
rect 1593 19465 1627 19499
rect 3893 19465 3927 19499
rect 5871 19465 5905 19499
rect 7849 19465 7883 19499
rect 9597 19465 9631 19499
rect 25145 19465 25179 19499
rect 1409 19261 1443 19295
rect 3484 19261 3518 19295
rect 5800 19261 5834 19295
rect 7941 19261 7975 19295
rect 9112 19261 9146 19295
rect 11380 19261 11414 19295
rect 11805 19261 11839 19295
rect 12541 19261 12575 19295
rect 24660 19261 24694 19295
rect 3571 19193 3605 19227
rect 8677 19193 8711 19227
rect 2053 19125 2087 19159
rect 6285 19125 6319 19159
rect 6653 19125 6687 19159
rect 6929 19125 6963 19159
rect 8125 19125 8159 19159
rect 9183 19125 9217 19159
rect 11483 19125 11517 19159
rect 12265 19125 12299 19159
rect 12725 19125 12759 19159
rect 24731 19125 24765 19159
rect 1593 18921 1627 18955
rect 7205 18921 7239 18955
rect 6377 18853 6411 18887
rect 7849 18853 7883 18887
rect 7941 18853 7975 18887
rect 9873 18853 9907 18887
rect 12265 18853 12299 18887
rect 12357 18853 12391 18887
rect 1869 18785 1903 18819
rect 5064 18785 5098 18819
rect 13804 18785 13838 18819
rect 18772 18785 18806 18819
rect 2099 18717 2133 18751
rect 6285 18717 6319 18751
rect 8493 18717 8527 18751
rect 9781 18717 9815 18751
rect 10425 18717 10459 18751
rect 17693 18717 17727 18751
rect 6837 18649 6871 18683
rect 12817 18649 12851 18683
rect 5135 18581 5169 18615
rect 13875 18581 13909 18615
rect 18843 18581 18877 18615
rect 1961 18377 1995 18411
rect 5181 18377 5215 18411
rect 6561 18377 6595 18411
rect 12725 18377 12759 18411
rect 13921 18377 13955 18411
rect 19349 18377 19383 18411
rect 24777 18377 24811 18411
rect 5871 18309 5905 18343
rect 10241 18309 10275 18343
rect 10563 18309 10597 18343
rect 18889 18309 18923 18343
rect 7113 18241 7147 18275
rect 8953 18241 8987 18275
rect 9229 18241 9263 18275
rect 10885 18241 10919 18275
rect 13185 18241 13219 18275
rect 19901 18241 19935 18275
rect 20177 18241 20211 18275
rect 1409 18173 1443 18207
rect 5800 18173 5834 18207
rect 10460 18173 10494 18207
rect 14540 18173 14574 18207
rect 14933 18173 14967 18207
rect 16992 18173 17026 18207
rect 17417 18173 17451 18207
rect 24593 18173 24627 18207
rect 25145 18173 25179 18207
rect 7205 18105 7239 18139
rect 7757 18105 7791 18139
rect 8769 18105 8803 18139
rect 9045 18105 9079 18139
rect 12265 18105 12299 18139
rect 12909 18105 12943 18139
rect 13001 18105 13035 18139
rect 17095 18105 17129 18139
rect 18337 18105 18371 18139
rect 18438 18105 18472 18139
rect 19717 18105 19751 18139
rect 19993 18105 20027 18139
rect 1547 18037 1581 18071
rect 4721 18037 4755 18071
rect 6285 18037 6319 18071
rect 8125 18037 8159 18071
rect 9965 18037 9999 18071
rect 11897 18037 11931 18071
rect 14611 18037 14645 18071
rect 17877 18037 17911 18071
rect 1593 17833 1627 17867
rect 6285 17833 6319 17867
rect 8217 17833 8251 17867
rect 8953 17833 8987 17867
rect 11621 17833 11655 17867
rect 12265 17833 12299 17867
rect 17049 17833 17083 17867
rect 18337 17833 18371 17867
rect 19901 17833 19935 17867
rect 20177 17833 20211 17867
rect 21557 17833 21591 17867
rect 24501 17833 24535 17867
rect 7297 17765 7331 17799
rect 7389 17765 7423 17799
rect 9873 17765 9907 17799
rect 12817 17765 12851 17799
rect 17325 17765 17359 17799
rect 17417 17765 17451 17799
rect 18889 17765 18923 17799
rect 18981 17765 19015 17799
rect 1409 17697 1443 17731
rect 2513 17697 2547 17731
rect 5457 17697 5491 17731
rect 15393 17697 15427 17731
rect 22604 17697 22638 17731
rect 22707 17697 22741 17731
rect 24317 17697 24351 17731
rect 7757 17629 7791 17663
rect 9781 17629 9815 17663
rect 12725 17629 12759 17663
rect 13185 17629 13219 17663
rect 14197 17629 14231 17663
rect 17969 17629 18003 17663
rect 19165 17629 19199 17663
rect 10333 17561 10367 17595
rect 2651 17493 2685 17527
rect 3525 17493 3559 17527
rect 5089 17493 5123 17527
rect 7113 17493 7147 17527
rect 15761 17493 15795 17527
rect 18613 17493 18647 17527
rect 3341 17289 3375 17323
rect 4629 17289 4663 17323
rect 4997 17289 5031 17323
rect 6101 17289 6135 17323
rect 6561 17289 6595 17323
rect 9137 17289 9171 17323
rect 10609 17289 10643 17323
rect 11621 17289 11655 17323
rect 15393 17289 15427 17323
rect 17325 17289 17359 17323
rect 17785 17289 17819 17323
rect 22569 17289 22603 17323
rect 24317 17289 24351 17323
rect 7757 17221 7791 17255
rect 20545 17221 20579 17255
rect 2881 17153 2915 17187
rect 3617 17153 3651 17187
rect 5181 17153 5215 17187
rect 7205 17153 7239 17187
rect 8125 17153 8159 17187
rect 11897 17153 11931 17187
rect 12541 17153 12575 17187
rect 12817 17153 12851 17187
rect 18245 17153 18279 17187
rect 18521 17153 18555 17187
rect 19993 17153 20027 17187
rect 21557 17153 21591 17187
rect 1961 17085 1995 17119
rect 2488 17085 2522 17119
rect 11253 17085 11287 17119
rect 11380 17085 11414 17119
rect 13921 17085 13955 17119
rect 14105 17085 14139 17119
rect 15669 17085 15703 17119
rect 16589 17085 16623 17119
rect 3709 17017 3743 17051
rect 4261 17017 4295 17051
rect 5273 17017 5307 17051
rect 5825 17017 5859 17051
rect 7297 17017 7331 17051
rect 9689 17017 9723 17051
rect 9781 17017 9815 17051
rect 10333 17017 10367 17051
rect 12633 17017 12667 17051
rect 14013 17017 14047 17051
rect 15577 17017 15611 17051
rect 18337 17017 18371 17051
rect 20085 17017 20119 17051
rect 21373 17017 21407 17051
rect 21649 17017 21683 17051
rect 22201 17017 22235 17051
rect 1409 16949 1443 16983
rect 2559 16949 2593 16983
rect 8769 16949 8803 16983
rect 9505 16949 9539 16983
rect 12265 16949 12299 16983
rect 13553 16949 13587 16983
rect 19165 16949 19199 16983
rect 19809 16949 19843 16983
rect 2513 16745 2547 16779
rect 7205 16745 7239 16779
rect 10057 16745 10091 16779
rect 10609 16745 10643 16779
rect 12817 16745 12851 16779
rect 17049 16745 17083 16779
rect 17601 16745 17635 16779
rect 4813 16677 4847 16711
rect 6377 16677 6411 16711
rect 7849 16677 7883 16711
rect 7941 16677 7975 16711
rect 11850 16677 11884 16711
rect 13461 16677 13495 16711
rect 19441 16677 19475 16711
rect 19993 16677 20027 16711
rect 21097 16677 21131 16711
rect 1869 16609 1903 16643
rect 12449 16609 12483 16643
rect 15301 16609 15335 16643
rect 15485 16609 15519 16643
rect 22477 16609 22511 16643
rect 4721 16541 4755 16575
rect 4997 16541 5031 16575
rect 6009 16541 6043 16575
rect 6285 16541 6319 16575
rect 6561 16541 6595 16575
rect 8125 16541 8159 16575
rect 9689 16541 9723 16575
rect 11529 16541 11563 16575
rect 13369 16541 13403 16575
rect 13645 16541 13679 16575
rect 15853 16541 15887 16575
rect 16129 16541 16163 16575
rect 16681 16541 16715 16575
rect 19349 16541 19383 16575
rect 21005 16541 21039 16575
rect 22615 16541 22649 16575
rect 18245 16473 18279 16507
rect 21557 16473 21591 16507
rect 1777 16405 1811 16439
rect 3617 16405 3651 16439
rect 4445 16405 4479 16439
rect 7665 16405 7699 16439
rect 8769 16405 8803 16439
rect 10885 16405 10919 16439
rect 18889 16405 18923 16439
rect 5365 16201 5399 16235
rect 6193 16201 6227 16235
rect 7941 16201 7975 16235
rect 9505 16201 9539 16235
rect 11529 16201 11563 16235
rect 13277 16201 13311 16235
rect 14289 16201 14323 16235
rect 14933 16201 14967 16235
rect 18337 16201 18371 16235
rect 19717 16201 19751 16235
rect 19993 16201 20027 16235
rect 21741 16201 21775 16235
rect 3617 16133 3651 16167
rect 10977 16133 11011 16167
rect 12909 16133 12943 16167
rect 14013 16133 14047 16167
rect 1593 16065 1627 16099
rect 2881 16065 2915 16099
rect 3985 16065 4019 16099
rect 7573 16065 7607 16099
rect 10425 16065 10459 16099
rect 13461 16065 13495 16099
rect 3132 15997 3166 16031
rect 4445 15997 4479 16031
rect 8585 15997 8619 16031
rect 1685 15929 1719 15963
rect 2237 15929 2271 15963
rect 5825 15929 5859 15963
rect 6929 15929 6963 15963
rect 7021 15929 7055 15963
rect 8906 15929 8940 15963
rect 9781 15929 9815 15963
rect 10517 15929 10551 15963
rect 13553 15929 13587 15963
rect 15163 16133 15197 16167
rect 16773 16065 16807 16099
rect 17417 16065 17451 16099
rect 18797 16065 18831 16099
rect 20821 16065 20855 16099
rect 22201 16065 22235 16099
rect 15060 15997 15094 16031
rect 15485 15997 15519 16031
rect 16037 15997 16071 16031
rect 16497 15997 16531 16031
rect 20545 15997 20579 16031
rect 19118 15929 19152 15963
rect 20913 15929 20947 15963
rect 21465 15929 21499 15963
rect 2513 15861 2547 15895
rect 3203 15861 3237 15895
rect 4353 15861 4387 15895
rect 4813 15861 4847 15895
rect 6653 15861 6687 15895
rect 8401 15861 8435 15895
rect 10149 15861 10183 15895
rect 11989 15861 12023 15895
rect 14289 15861 14323 15895
rect 14381 15861 14415 15895
rect 15853 15861 15887 15895
rect 17049 15861 17083 15895
rect 18613 15861 18647 15895
rect 22477 15861 22511 15895
rect 2697 15657 2731 15691
rect 3893 15657 3927 15691
rect 4997 15657 5031 15691
rect 7021 15657 7055 15691
rect 7849 15657 7883 15691
rect 8723 15657 8757 15691
rect 10609 15657 10643 15691
rect 12357 15657 12391 15691
rect 16037 15657 16071 15691
rect 17325 15657 17359 15691
rect 19441 15657 19475 15691
rect 19993 15657 20027 15691
rect 20729 15657 20763 15691
rect 24777 15657 24811 15691
rect 1777 15589 1811 15623
rect 1869 15589 1903 15623
rect 2421 15589 2455 15623
rect 4398 15589 4432 15623
rect 10051 15589 10085 15623
rect 11758 15589 11792 15623
rect 13737 15589 13771 15623
rect 13829 15589 13863 15623
rect 16726 15589 16760 15623
rect 21189 15589 21223 15623
rect 21741 15589 21775 15623
rect 22753 15589 22787 15623
rect 7573 15521 7607 15555
rect 8585 15521 8619 15555
rect 15368 15521 15402 15555
rect 24593 15521 24627 15555
rect 4077 15453 4111 15487
rect 6653 15453 6687 15487
rect 9689 15453 9723 15487
rect 11437 15453 11471 15487
rect 12633 15453 12667 15487
rect 14381 15453 14415 15487
rect 16405 15453 16439 15487
rect 19073 15453 19107 15487
rect 20361 15453 20395 15487
rect 21097 15453 21131 15487
rect 22661 15453 22695 15487
rect 22937 15453 22971 15487
rect 13001 15385 13035 15419
rect 3065 15317 3099 15351
rect 5549 15317 5583 15351
rect 6193 15317 6227 15351
rect 6561 15317 6595 15351
rect 9045 15317 9079 15351
rect 9413 15317 9447 15351
rect 10977 15317 11011 15351
rect 11253 15317 11287 15351
rect 13369 15317 13403 15351
rect 15439 15317 15473 15351
rect 18061 15317 18095 15351
rect 18981 15317 19015 15351
rect 2697 15113 2731 15147
rect 2973 15113 3007 15147
rect 5687 15113 5721 15147
rect 7757 15113 7791 15147
rect 8585 15113 8619 15147
rect 9781 15113 9815 15147
rect 11621 15113 11655 15147
rect 12173 15113 12207 15147
rect 13369 15113 13403 15147
rect 15393 15113 15427 15147
rect 17417 15113 17451 15147
rect 18981 15113 19015 15147
rect 20913 15113 20947 15147
rect 22845 15113 22879 15147
rect 5365 15045 5399 15079
rect 24777 15045 24811 15079
rect 3985 14977 4019 15011
rect 4997 14977 5031 15011
rect 6837 14977 6871 15011
rect 8861 14977 8895 15011
rect 14289 14977 14323 15011
rect 14565 14977 14599 15011
rect 17141 14977 17175 15011
rect 18061 14977 18095 15011
rect 23121 14977 23155 15011
rect 1777 14909 1811 14943
rect 3341 14909 3375 14943
rect 4629 14909 4663 14943
rect 5549 14909 5583 14943
rect 10057 14909 10091 14943
rect 10517 14909 10551 14943
rect 10885 14909 10919 14943
rect 11161 14909 11195 14943
rect 12449 14909 12483 14943
rect 16405 14909 16439 14943
rect 16865 14909 16899 14943
rect 19993 14909 20027 14943
rect 21741 14909 21775 14943
rect 22201 14909 22235 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 2098 14841 2132 14875
rect 3801 14841 3835 14875
rect 6193 14841 6227 14875
rect 6561 14841 6595 14875
rect 7158 14841 7192 14875
rect 8217 14841 8251 14875
rect 9182 14841 9216 14875
rect 12770 14841 12804 14875
rect 14381 14841 14415 14875
rect 18382 14841 18416 14875
rect 19257 14841 19291 14875
rect 19809 14841 19843 14875
rect 20314 14841 20348 14875
rect 1685 14773 1719 14807
rect 10701 14773 10735 14807
rect 13737 14773 13771 14807
rect 14105 14773 14139 14807
rect 15853 14773 15887 14807
rect 16221 14773 16255 14807
rect 17785 14773 17819 14807
rect 21189 14773 21223 14807
rect 21649 14773 21683 14807
rect 21833 14773 21867 14807
rect 24409 14773 24443 14807
rect 2605 14569 2639 14603
rect 4169 14569 4203 14603
rect 6745 14569 6779 14603
rect 9137 14569 9171 14603
rect 9505 14569 9539 14603
rect 12909 14569 12943 14603
rect 14289 14569 14323 14603
rect 14749 14569 14783 14603
rect 16773 14569 16807 14603
rect 17417 14569 17451 14603
rect 20729 14569 20763 14603
rect 22661 14569 22695 14603
rect 23765 14569 23799 14603
rect 1777 14501 1811 14535
rect 7573 14501 7607 14535
rect 7941 14501 7975 14535
rect 8769 14501 8803 14535
rect 12265 14501 12299 14535
rect 13414 14501 13448 14535
rect 15945 14501 15979 14535
rect 19717 14501 19751 14535
rect 19993 14501 20027 14535
rect 2973 14433 3007 14467
rect 4261 14433 4295 14467
rect 4721 14433 4755 14467
rect 5089 14433 5123 14467
rect 5457 14433 5491 14467
rect 6561 14433 6595 14467
rect 7021 14433 7055 14467
rect 8033 14433 8067 14467
rect 8585 14433 8619 14467
rect 9848 14433 9882 14467
rect 10701 14433 10735 14467
rect 10793 14433 10827 14467
rect 11529 14433 11563 14467
rect 11621 14433 11655 14467
rect 11989 14433 12023 14467
rect 17325 14433 17359 14467
rect 17785 14433 17819 14467
rect 18981 14433 19015 14467
rect 19441 14433 19475 14467
rect 20913 14433 20947 14467
rect 21373 14433 21407 14467
rect 22477 14433 22511 14467
rect 23581 14433 23615 14467
rect 1685 14365 1719 14399
rect 3525 14365 3559 14399
rect 6377 14365 6411 14399
rect 13093 14365 13127 14399
rect 15853 14365 15887 14399
rect 21465 14365 21499 14399
rect 2237 14297 2271 14331
rect 14013 14297 14047 14331
rect 16405 14297 16439 14331
rect 3893 14229 3927 14263
rect 9919 14229 9953 14263
rect 10333 14229 10367 14263
rect 12541 14229 12575 14263
rect 21925 14229 21959 14263
rect 2881 14025 2915 14059
rect 9597 14025 9631 14059
rect 15577 14025 15611 14059
rect 16773 14025 16807 14059
rect 17325 14025 17359 14059
rect 17785 14025 17819 14059
rect 18429 14025 18463 14059
rect 21373 14025 21407 14059
rect 22661 14025 22695 14059
rect 24133 14025 24167 14059
rect 3157 13957 3191 13991
rect 4169 13957 4203 13991
rect 11437 13957 11471 13991
rect 24501 13957 24535 13991
rect 1501 13889 1535 13923
rect 2145 13889 2179 13923
rect 6561 13889 6595 13923
rect 11805 13889 11839 13923
rect 16405 13889 16439 13923
rect 23811 13889 23845 13923
rect 2973 13821 3007 13855
rect 4261 13821 4295 13855
rect 4721 13821 4755 13855
rect 5089 13821 5123 13855
rect 5457 13821 5491 13855
rect 7113 13821 7147 13855
rect 7389 13821 7423 13855
rect 8677 13821 8711 13855
rect 8861 13821 8895 13855
rect 9873 13821 9907 13855
rect 10057 13821 10091 13855
rect 10517 13821 10551 13855
rect 11069 13821 11103 13855
rect 11253 13821 11287 13855
rect 12449 13821 12483 13855
rect 12909 13821 12943 13855
rect 13277 13821 13311 13855
rect 13645 13821 13679 13855
rect 13921 13821 13955 13855
rect 14197 13821 14231 13855
rect 15209 13821 15243 13855
rect 18889 13821 18923 13855
rect 19165 13821 19199 13855
rect 19441 13821 19475 13855
rect 23708 13821 23742 13855
rect 1593 13753 1627 13787
rect 2421 13753 2455 13787
rect 3801 13753 3835 13787
rect 6101 13753 6135 13787
rect 14841 13753 14875 13787
rect 15761 13753 15795 13787
rect 15853 13753 15887 13787
rect 19717 13753 19751 13787
rect 21741 13753 21775 13787
rect 21833 13753 21867 13787
rect 22385 13753 22419 13787
rect 4353 13685 4387 13719
rect 6929 13685 6963 13719
rect 8033 13685 8067 13719
rect 8493 13685 8527 13719
rect 12265 13685 12299 13719
rect 20545 13685 20579 13719
rect 21005 13685 21039 13719
rect 2421 13481 2455 13515
rect 2697 13481 2731 13515
rect 4169 13481 4203 13515
rect 7849 13481 7883 13515
rect 9045 13481 9079 13515
rect 10793 13481 10827 13515
rect 12081 13481 12115 13515
rect 12633 13481 12667 13515
rect 13093 13481 13127 13515
rect 14381 13481 14415 13515
rect 19441 13481 19475 13515
rect 1822 13413 1856 13447
rect 6561 13413 6595 13447
rect 7113 13413 7147 13447
rect 8769 13413 8803 13447
rect 13782 13413 13816 13447
rect 15301 13413 15335 13447
rect 18153 13413 18187 13447
rect 21465 13413 21499 13447
rect 3525 13345 3559 13379
rect 4353 13345 4387 13379
rect 4537 13345 4571 13379
rect 5089 13345 5123 13379
rect 5457 13345 5491 13379
rect 8309 13345 8343 13379
rect 8493 13345 8527 13379
rect 10425 13345 10459 13379
rect 11161 13345 11195 13379
rect 11621 13345 11655 13379
rect 11713 13345 11747 13379
rect 12265 13345 12299 13379
rect 15393 13345 15427 13379
rect 16865 13345 16899 13379
rect 19533 13345 19567 13379
rect 24660 13345 24694 13379
rect 1501 13277 1535 13311
rect 3065 13277 3099 13311
rect 6469 13277 6503 13311
rect 9873 13277 9907 13311
rect 13461 13277 13495 13311
rect 18061 13277 18095 13311
rect 21373 13277 21407 13311
rect 5917 13209 5951 13243
rect 17785 13209 17819 13243
rect 18613 13209 18647 13243
rect 21925 13209 21959 13243
rect 3801 13141 3835 13175
rect 6285 13141 6319 13175
rect 7481 13141 7515 13175
rect 9413 13141 9447 13175
rect 17003 13141 17037 13175
rect 19073 13141 19107 13175
rect 19717 13141 19751 13175
rect 22293 13141 22327 13175
rect 24731 13141 24765 13175
rect 1685 12937 1719 12971
rect 3525 12937 3559 12971
rect 5825 12937 5859 12971
rect 9413 12937 9447 12971
rect 11529 12937 11563 12971
rect 14197 12937 14231 12971
rect 15393 12937 15427 12971
rect 16865 12937 16899 12971
rect 17509 12937 17543 12971
rect 18981 12937 19015 12971
rect 21005 12937 21039 12971
rect 21373 12937 21407 12971
rect 24501 12937 24535 12971
rect 24777 12937 24811 12971
rect 7849 12869 7883 12903
rect 8493 12869 8527 12903
rect 11161 12869 11195 12903
rect 12265 12869 12299 12903
rect 21833 12869 21867 12903
rect 2789 12801 2823 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 8861 12801 8895 12835
rect 15577 12801 15611 12835
rect 16497 12801 16531 12835
rect 19809 12801 19843 12835
rect 22109 12801 22143 12835
rect 22477 12801 22511 12835
rect 23029 12801 23063 12835
rect 2053 12733 2087 12767
rect 3893 12733 3927 12767
rect 4169 12733 4203 12767
rect 4629 12733 4663 12767
rect 4997 12733 5031 12767
rect 8401 12733 8435 12767
rect 8677 12733 8711 12767
rect 10701 12733 10735 12767
rect 12449 12733 12483 12767
rect 13093 12733 13127 12767
rect 13277 12733 13311 12767
rect 13645 12733 13679 12767
rect 18061 12733 18095 12767
rect 3157 12665 3191 12699
rect 7021 12665 7055 12699
rect 9873 12665 9907 12699
rect 10057 12665 10091 12699
rect 11897 12665 11931 12699
rect 13921 12665 13955 12699
rect 14565 12665 14599 12699
rect 15025 12665 15059 12699
rect 15669 12665 15703 12699
rect 16221 12665 16255 12699
rect 18382 12665 18416 12699
rect 19625 12665 19659 12699
rect 20085 12733 20119 12767
rect 24593 12733 24627 12767
rect 20406 12665 20440 12699
rect 22201 12665 22235 12699
rect 25237 12665 25271 12699
rect 3709 12597 3743 12631
rect 5365 12597 5399 12631
rect 6377 12597 6411 12631
rect 8217 12597 8251 12631
rect 17785 12597 17819 12631
rect 19809 12597 19843 12631
rect 19901 12597 19935 12631
rect 3709 12393 3743 12427
rect 4261 12393 4295 12427
rect 12449 12393 12483 12427
rect 12909 12393 12943 12427
rect 16221 12393 16255 12427
rect 17417 12393 17451 12427
rect 18613 12393 18647 12427
rect 18889 12393 18923 12427
rect 22293 12393 22327 12427
rect 1685 12325 1719 12359
rect 2053 12325 2087 12359
rect 2513 12325 2547 12359
rect 7894 12325 7928 12359
rect 9873 12325 9907 12359
rect 11345 12325 11379 12359
rect 11437 12325 11471 12359
rect 15622 12325 15656 12359
rect 21373 12325 21407 12359
rect 21925 12325 21959 12359
rect 22937 12325 22971 12359
rect 24501 12325 24535 12359
rect 4077 12257 4111 12291
rect 5549 12257 5583 12291
rect 5733 12257 5767 12291
rect 6285 12257 6319 12291
rect 6653 12257 6687 12291
rect 7481 12257 7515 12291
rect 10977 12257 11011 12291
rect 13737 12257 13771 12291
rect 14197 12257 14231 12291
rect 18981 12257 19015 12291
rect 19349 12257 19383 12291
rect 2421 12189 2455 12223
rect 4721 12189 4755 12223
rect 6745 12189 6779 12223
rect 7573 12189 7607 12223
rect 9137 12189 9171 12223
rect 9781 12189 9815 12223
rect 10149 12189 10183 12223
rect 11989 12189 12023 12223
rect 14381 12189 14415 12223
rect 15301 12189 15335 12223
rect 17049 12189 17083 12223
rect 21281 12189 21315 12223
rect 22845 12189 22879 12223
rect 23121 12189 23155 12223
rect 24409 12189 24443 12223
rect 24685 12189 24719 12223
rect 2973 12121 3007 12155
rect 4997 12121 5031 12155
rect 13369 12121 13403 12155
rect 7021 12053 7055 12087
rect 8493 12053 8527 12087
rect 8861 12053 8895 12087
rect 17969 12053 18003 12087
rect 18245 12053 18279 12087
rect 20085 12053 20119 12087
rect 2145 11849 2179 11883
rect 3709 11849 3743 11883
rect 7665 11849 7699 11883
rect 9413 11849 9447 11883
rect 11989 11849 12023 11883
rect 14749 11849 14783 11883
rect 16497 11849 16531 11883
rect 20913 11849 20947 11883
rect 21281 11849 21315 11883
rect 23397 11849 23431 11883
rect 24041 11849 24075 11883
rect 24317 11849 24351 11883
rect 24777 11849 24811 11883
rect 3985 11781 4019 11815
rect 6653 11781 6687 11815
rect 21833 11781 21867 11815
rect 2973 11713 3007 11747
rect 5733 11713 5767 11747
rect 7297 11713 7331 11747
rect 9413 11713 9447 11747
rect 9505 11713 9539 11747
rect 9873 11713 9907 11747
rect 14473 11713 14507 11747
rect 16819 11713 16853 11747
rect 18153 11713 18187 11747
rect 18429 11713 18463 11747
rect 19441 11713 19475 11747
rect 19993 11713 20027 11747
rect 22109 11713 22143 11747
rect 22477 11713 22511 11747
rect 1409 11645 1443 11679
rect 4261 11645 4295 11679
rect 8033 11645 8067 11679
rect 8401 11645 8435 11679
rect 8769 11645 8803 11679
rect 8953 11645 8987 11679
rect 9229 11645 9263 11679
rect 10057 11645 10091 11679
rect 13277 11645 13311 11679
rect 13645 11645 13679 11679
rect 13829 11645 13863 11679
rect 14105 11645 14139 11679
rect 14933 11645 14967 11679
rect 16716 11645 16750 11679
rect 17141 11645 17175 11679
rect 19809 11645 19843 11679
rect 23029 11645 23063 11679
rect 24593 11645 24627 11679
rect 25145 11645 25179 11679
rect 2697 11577 2731 11611
rect 2789 11577 2823 11611
rect 4169 11577 4203 11611
rect 10378 11577 10412 11611
rect 11345 11577 11379 11611
rect 11713 11577 11747 11611
rect 15254 11577 15288 11611
rect 16129 11577 16163 11611
rect 17509 11577 17543 11611
rect 18245 11577 18279 11611
rect 20314 11577 20348 11611
rect 22201 11577 22235 11611
rect 1593 11509 1627 11543
rect 2513 11509 2547 11543
rect 5365 11509 5399 11543
rect 6285 11509 6319 11543
rect 10977 11509 11011 11543
rect 12817 11509 12851 11543
rect 15853 11509 15887 11543
rect 19073 11509 19107 11543
rect 4169 11305 4203 11339
rect 5917 11305 5951 11339
rect 6193 11305 6227 11339
rect 9045 11305 9079 11339
rect 10609 11305 10643 11339
rect 10885 11305 10919 11339
rect 12817 11305 12851 11339
rect 14933 11305 14967 11339
rect 16957 11305 16991 11339
rect 17141 11305 17175 11339
rect 18153 11305 18187 11339
rect 20453 11305 20487 11339
rect 21097 11305 21131 11339
rect 21419 11305 21453 11339
rect 23995 11305 24029 11339
rect 2558 11237 2592 11271
rect 6377 11237 6411 11271
rect 8677 11237 8711 11271
rect 10030 11237 10064 11271
rect 11253 11237 11287 11271
rect 11621 11237 11655 11271
rect 15669 11237 15703 11271
rect 16221 11237 16255 11271
rect 19809 11237 19843 11271
rect 22477 11237 22511 11271
rect 4353 11169 4387 11203
rect 4813 11169 4847 11203
rect 4997 11169 5031 11203
rect 5457 11169 5491 11203
rect 7021 11169 7055 11203
rect 8033 11169 8067 11203
rect 13461 11169 13495 11203
rect 17049 11169 17083 11203
rect 17601 11169 17635 11203
rect 19073 11169 19107 11203
rect 19533 11169 19567 11203
rect 21316 11169 21350 11203
rect 23892 11169 23926 11203
rect 2237 11101 2271 11135
rect 3893 11101 3927 11135
rect 9689 11101 9723 11135
rect 11529 11101 11563 11135
rect 11805 11101 11839 11135
rect 13001 11101 13035 11135
rect 14657 11101 14691 11135
rect 15577 11101 15611 11135
rect 22385 11101 22419 11135
rect 22661 11101 22695 11135
rect 3157 11033 3191 11067
rect 1685 10965 1719 10999
rect 1961 10965 1995 10999
rect 3433 10965 3467 10999
rect 7481 10965 7515 10999
rect 7757 10965 7791 10999
rect 9321 10965 9355 10999
rect 12541 10965 12575 10999
rect 20085 10965 20119 10999
rect 22109 10965 22143 10999
rect 2421 10761 2455 10795
rect 2789 10761 2823 10795
rect 4445 10761 4479 10795
rect 9965 10761 9999 10795
rect 10333 10761 10367 10795
rect 13461 10761 13495 10795
rect 17095 10761 17129 10795
rect 22017 10761 22051 10795
rect 22707 10761 22741 10795
rect 23811 10761 23845 10795
rect 4077 10693 4111 10727
rect 22385 10693 22419 10727
rect 1501 10625 1535 10659
rect 3065 10625 3099 10659
rect 5917 10625 5951 10659
rect 7389 10625 7423 10659
rect 10609 10625 10643 10659
rect 10977 10625 11011 10659
rect 12817 10625 12851 10659
rect 14933 10625 14967 10659
rect 18521 10625 18555 10659
rect 20177 10625 20211 10659
rect 24501 10625 24535 10659
rect 5181 10557 5215 10591
rect 5273 10557 5307 10591
rect 5457 10557 5491 10591
rect 6837 10557 6871 10591
rect 7021 10557 7055 10591
rect 8217 10557 8251 10591
rect 8677 10557 8711 10591
rect 9229 10557 9263 10591
rect 9413 10557 9447 10591
rect 13829 10557 13863 10591
rect 14013 10557 14047 10591
rect 14197 10557 14231 10591
rect 14565 10557 14599 10591
rect 15301 10557 15335 10591
rect 15577 10557 15611 10591
rect 15945 10557 15979 10591
rect 16129 10557 16163 10591
rect 16992 10557 17026 10591
rect 17877 10557 17911 10591
rect 18245 10557 18279 10591
rect 22604 10557 22638 10591
rect 23121 10557 23155 10591
rect 23740 10557 23774 10591
rect 23949 10557 23983 10591
rect 24720 10557 24754 10591
rect 25145 10557 25179 10591
rect 1593 10489 1627 10523
rect 2145 10489 2179 10523
rect 3157 10489 3191 10523
rect 3709 10489 3743 10523
rect 9689 10489 9723 10523
rect 10701 10489 10735 10523
rect 12541 10489 12575 10523
rect 12633 10489 12667 10523
rect 17417 10489 17451 10523
rect 18061 10489 18095 10523
rect 19257 10489 19291 10523
rect 19533 10489 19567 10523
rect 19625 10489 19659 10523
rect 21097 10489 21131 10523
rect 21189 10489 21223 10523
rect 21741 10489 21775 10523
rect 24823 10489 24857 10523
rect 4997 10421 5031 10455
rect 6193 10421 6227 10455
rect 6561 10421 6595 10455
rect 7665 10421 7699 10455
rect 8033 10421 8067 10455
rect 11621 10421 11655 10455
rect 12265 10421 12299 10455
rect 16497 10421 16531 10455
rect 16773 10421 16807 10455
rect 18981 10421 19015 10455
rect 20453 10421 20487 10455
rect 20913 10421 20947 10455
rect 23949 10421 23983 10455
rect 24225 10421 24259 10455
rect 2605 10217 2639 10251
rect 3065 10217 3099 10251
rect 3893 10217 3927 10251
rect 4353 10217 4387 10251
rect 7757 10217 7791 10251
rect 9413 10217 9447 10251
rect 9873 10217 9907 10251
rect 11621 10217 11655 10251
rect 11989 10217 12023 10251
rect 15117 10217 15151 10251
rect 16957 10217 16991 10251
rect 19625 10217 19659 10251
rect 21833 10217 21867 10251
rect 24317 10217 24351 10251
rect 2047 10149 2081 10183
rect 7113 10149 7147 10183
rect 10793 10149 10827 10183
rect 17141 10149 17175 10183
rect 17233 10149 17267 10183
rect 19067 10149 19101 10183
rect 19901 10149 19935 10183
rect 21234 10149 21268 10183
rect 22845 10149 22879 10183
rect 4077 10081 4111 10115
rect 4813 10081 4847 10115
rect 5089 10081 5123 10115
rect 5457 10081 5491 10115
rect 6101 10081 6135 10115
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 7389 10081 7423 10115
rect 8125 10081 8159 10115
rect 12173 10081 12207 10115
rect 12725 10081 12759 10115
rect 13737 10081 13771 10115
rect 13921 10081 13955 10115
rect 15669 10081 15703 10115
rect 15853 10081 15887 10115
rect 18153 10081 18187 10115
rect 24225 10081 24259 10115
rect 24777 10081 24811 10115
rect 1685 10013 1719 10047
rect 5917 9945 5951 9979
rect 8033 10013 8067 10047
rect 9045 10013 9079 10047
rect 10701 10013 10735 10047
rect 10977 10013 11011 10047
rect 12909 10013 12943 10047
rect 14197 10013 14231 10047
rect 16129 10013 16163 10047
rect 18705 10013 18739 10047
rect 20913 10013 20947 10047
rect 22753 10013 22787 10047
rect 23029 10013 23063 10047
rect 6469 9945 6503 9979
rect 14565 9945 14599 9979
rect 17693 9945 17727 9979
rect 20269 9945 20303 9979
rect 3433 9877 3467 9911
rect 6101 9877 6135 9911
rect 6193 9877 6227 9911
rect 10241 9877 10275 9911
rect 16405 9877 16439 9911
rect 22293 9877 22327 9911
rect 1685 9673 1719 9707
rect 2421 9673 2455 9707
rect 2973 9673 3007 9707
rect 4077 9673 4111 9707
rect 6193 9673 6227 9707
rect 8953 9673 8987 9707
rect 10793 9673 10827 9707
rect 11483 9673 11517 9707
rect 13093 9673 13127 9707
rect 13277 9673 13311 9707
rect 13645 9673 13679 9707
rect 15117 9673 15151 9707
rect 16037 9673 16071 9707
rect 19165 9673 19199 9707
rect 19441 9673 19475 9707
rect 22661 9673 22695 9707
rect 25053 9673 25087 9707
rect 25789 9673 25823 9707
rect 10609 9605 10643 9639
rect 11253 9605 11287 9639
rect 5273 9537 5307 9571
rect 6653 9537 6687 9571
rect 2053 9469 2087 9503
rect 3525 9469 3559 9503
rect 4261 9469 4295 9503
rect 5181 9469 5215 9503
rect 5457 9469 5491 9503
rect 7481 9469 7515 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 8585 9469 8619 9503
rect 5089 9401 5123 9435
rect 5917 9401 5951 9435
rect 7113 9401 7147 9435
rect 9873 9401 9907 9435
rect 9965 9401 9999 9435
rect 10517 9401 10551 9435
rect 21373 9605 21407 9639
rect 13829 9537 13863 9571
rect 18429 9537 18463 9571
rect 21925 9537 21959 9571
rect 23029 9537 23063 9571
rect 23397 9537 23431 9571
rect 11396 9469 11430 9503
rect 11897 9469 11931 9503
rect 12776 9469 12810 9503
rect 13093 9469 13127 9503
rect 16129 9469 16163 9503
rect 17325 9469 17359 9503
rect 19625 9469 19659 9503
rect 23673 9469 23707 9503
rect 24225 9469 24259 9503
rect 24685 9469 24719 9503
rect 25304 9469 25338 9503
rect 13921 9401 13955 9435
rect 14473 9401 14507 9435
rect 18153 9401 18187 9435
rect 18245 9401 18279 9435
rect 19946 9401 19980 9435
rect 20913 9401 20947 9435
rect 21649 9401 21683 9435
rect 21741 9401 21775 9435
rect 4721 9333 4755 9367
rect 7297 9333 7331 9367
rect 9597 9333 9631 9367
rect 10609 9333 10643 9367
rect 12173 9333 12207 9367
rect 12863 9333 12897 9367
rect 15485 9333 15519 9367
rect 16497 9333 16531 9367
rect 17049 9333 17083 9367
rect 17877 9333 17911 9367
rect 20545 9333 20579 9367
rect 23765 9333 23799 9367
rect 25375 9333 25409 9367
rect 1409 9129 1443 9163
rect 1961 9129 1995 9163
rect 2329 9129 2363 9163
rect 3525 9129 3559 9163
rect 6377 9129 6411 9163
rect 6745 9129 6779 9163
rect 7205 9129 7239 9163
rect 12541 9129 12575 9163
rect 13369 9129 13403 9163
rect 14197 9129 14231 9163
rect 17325 9129 17359 9163
rect 18797 9129 18831 9163
rect 19165 9129 19199 9163
rect 23673 9129 23707 9163
rect 5825 9061 5859 9095
rect 9873 9061 9907 9095
rect 16450 9061 16484 9095
rect 18198 9061 18232 9095
rect 21097 9061 21131 9095
rect 21925 9061 21959 9095
rect 22661 9061 22695 9095
rect 23213 9061 23247 9095
rect 2421 8993 2455 9027
rect 2697 8993 2731 9027
rect 4144 8993 4178 9027
rect 4537 8993 4571 9027
rect 5549 8993 5583 9027
rect 7573 8993 7607 9027
rect 7849 8993 7883 9027
rect 8125 8993 8159 9027
rect 8677 8993 8711 9027
rect 11713 8993 11747 9027
rect 11989 8993 12023 9027
rect 13921 8993 13955 9027
rect 14565 8993 14599 9027
rect 16129 8993 16163 9027
rect 17877 8993 17911 9027
rect 19860 8993 19894 9027
rect 25053 8993 25087 9027
rect 3157 8925 3191 8959
rect 3801 8925 3835 8959
rect 8769 8925 8803 8959
rect 9781 8925 9815 8959
rect 12173 8925 12207 8959
rect 13001 8925 13035 8959
rect 19947 8925 19981 8959
rect 21005 8925 21039 8959
rect 21281 8925 21315 8959
rect 22569 8925 22603 8959
rect 24041 8925 24075 8959
rect 2513 8857 2547 8891
rect 10333 8857 10367 8891
rect 19717 8857 19751 8891
rect 4215 8789 4249 8823
rect 4997 8789 5031 8823
rect 17049 8789 17083 8823
rect 17693 8789 17727 8823
rect 20637 8789 20671 8823
rect 25191 8789 25225 8823
rect 2513 8585 2547 8619
rect 2789 8585 2823 8619
rect 5825 8585 5859 8619
rect 6653 8585 6687 8619
rect 9413 8585 9447 8619
rect 10793 8585 10827 8619
rect 17785 8585 17819 8619
rect 21097 8585 21131 8619
rect 22661 8585 22695 8619
rect 22937 8585 22971 8619
rect 25145 8585 25179 8619
rect 3157 8517 3191 8551
rect 11253 8517 11287 8551
rect 16037 8517 16071 8551
rect 17509 8517 17543 8551
rect 20729 8517 20763 8551
rect 2145 8449 2179 8483
rect 3617 8449 3651 8483
rect 7849 8449 7883 8483
rect 9597 8449 9631 8483
rect 11345 8449 11379 8483
rect 12909 8449 12943 8483
rect 14105 8449 14139 8483
rect 15025 8449 15059 8483
rect 15761 8449 15795 8483
rect 19165 8449 19199 8483
rect 19717 8449 19751 8483
rect 20361 8449 20395 8483
rect 21281 8449 21315 8483
rect 21649 8449 21683 8483
rect 1685 8381 1719 8415
rect 2973 8381 3007 8415
rect 4353 8381 4387 8415
rect 4813 8381 4847 8415
rect 5089 8381 5123 8415
rect 5457 8381 5491 8415
rect 7389 8381 7423 8415
rect 16497 8381 16531 8415
rect 16681 8381 16715 8415
rect 18337 8381 18371 8415
rect 18613 8381 18647 8415
rect 18797 8381 18831 8415
rect 3985 8313 4019 8347
rect 8170 8313 8204 8347
rect 9918 8313 9952 8347
rect 12173 8313 12207 8347
rect 12725 8313 12759 8347
rect 13230 8313 13264 8347
rect 14749 8313 14783 8347
rect 14841 8313 14875 8347
rect 19533 8313 19567 8347
rect 19809 8313 19843 8347
rect 21373 8313 21407 8347
rect 4169 8245 4203 8279
rect 7665 8245 7699 8279
rect 8769 8245 8803 8279
rect 9137 8245 9171 8279
rect 10517 8245 10551 8279
rect 11805 8245 11839 8279
rect 13829 8245 13863 8279
rect 14473 8245 14507 8279
rect 16313 8245 16347 8279
rect 22201 8245 22235 8279
rect 1547 8041 1581 8075
rect 2237 8041 2271 8075
rect 3525 8041 3559 8075
rect 4353 8041 4387 8075
rect 7481 8041 7515 8075
rect 7849 8041 7883 8075
rect 9413 8041 9447 8075
rect 12817 8041 12851 8075
rect 14841 8041 14875 8075
rect 16957 8041 16991 8075
rect 18245 8041 18279 8075
rect 18521 8041 18555 8075
rect 20637 8041 20671 8075
rect 2605 7973 2639 8007
rect 8217 7973 8251 8007
rect 9873 7973 9907 8007
rect 11437 7973 11471 8007
rect 17325 7973 17359 8007
rect 18889 7973 18923 8007
rect 21097 7973 21131 8007
rect 21649 7973 21683 8007
rect 1476 7905 1510 7939
rect 4629 7905 4663 7939
rect 5365 7905 5399 7939
rect 5641 7905 5675 7939
rect 6009 7905 6043 7939
rect 6964 7905 6998 7939
rect 13001 7905 13035 7939
rect 13277 7905 13311 7939
rect 15853 7905 15887 7939
rect 16129 7905 16163 7939
rect 22544 7905 22578 7939
rect 2513 7837 2547 7871
rect 3157 7837 3191 7871
rect 6101 7837 6135 7871
rect 6377 7837 6411 7871
rect 8125 7837 8159 7871
rect 8769 7837 8803 7871
rect 9781 7837 9815 7871
rect 10057 7837 10091 7871
rect 11345 7837 11379 7871
rect 11621 7837 11655 7871
rect 13737 7837 13771 7871
rect 16313 7837 16347 7871
rect 17233 7837 17267 7871
rect 17693 7837 17727 7871
rect 18797 7837 18831 7871
rect 21005 7837 21039 7871
rect 1869 7769 1903 7803
rect 3893 7769 3927 7803
rect 13093 7769 13127 7803
rect 19349 7769 19383 7803
rect 22615 7769 22649 7803
rect 7067 7701 7101 7735
rect 14565 7701 14599 7735
rect 16589 7701 16623 7735
rect 19901 7701 19935 7735
rect 21925 7701 21959 7735
rect 1593 7497 1627 7531
rect 2145 7497 2179 7531
rect 6193 7497 6227 7531
rect 6653 7497 6687 7531
rect 8033 7497 8067 7531
rect 8953 7497 8987 7531
rect 11253 7497 11287 7531
rect 12265 7497 12299 7531
rect 12817 7497 12851 7531
rect 14013 7497 14047 7531
rect 16221 7497 16255 7531
rect 17417 7497 17451 7531
rect 21603 7497 21637 7531
rect 23029 7497 23063 7531
rect 23811 7497 23845 7531
rect 8401 7429 8435 7463
rect 10057 7429 10091 7463
rect 15669 7429 15703 7463
rect 21005 7429 21039 7463
rect 3249 7361 3283 7395
rect 4997 7361 5031 7395
rect 7205 7361 7239 7395
rect 13001 7361 13035 7395
rect 13461 7361 13495 7395
rect 14565 7361 14599 7395
rect 18153 7361 18187 7395
rect 22615 7361 22649 7395
rect 1409 7293 1443 7327
rect 4721 7293 4755 7327
rect 11412 7293 11446 7327
rect 14289 7293 14323 7327
rect 16405 7293 16439 7327
rect 16865 7293 16899 7327
rect 21500 7293 21534 7327
rect 21925 7293 21959 7327
rect 22528 7293 22562 7327
rect 23305 7293 23339 7327
rect 23740 7293 23774 7327
rect 24133 7293 24167 7327
rect 3065 7225 3099 7259
rect 3570 7225 3604 7259
rect 5359 7225 5393 7259
rect 6929 7225 6963 7259
rect 7021 7225 7055 7259
rect 9505 7225 9539 7259
rect 9597 7225 9631 7259
rect 11621 7225 11655 7259
rect 13093 7225 13127 7259
rect 14657 7225 14691 7259
rect 15209 7225 15243 7259
rect 17141 7225 17175 7259
rect 18245 7225 18279 7259
rect 18797 7225 18831 7259
rect 19993 7225 20027 7259
rect 20085 7225 20119 7259
rect 20637 7225 20671 7259
rect 2421 7157 2455 7191
rect 4169 7157 4203 7191
rect 5917 7157 5951 7191
rect 9321 7157 9355 7191
rect 10425 7157 10459 7191
rect 10793 7157 10827 7191
rect 11897 7157 11931 7191
rect 17785 7157 17819 7191
rect 19073 7157 19107 7191
rect 19717 7157 19751 7191
rect 21281 7157 21315 7191
rect 1869 6953 1903 6987
rect 3525 6953 3559 6987
rect 3801 6953 3835 6987
rect 5181 6953 5215 6987
rect 5549 6953 5583 6987
rect 7665 6953 7699 6987
rect 9505 6953 9539 6987
rect 11161 6953 11195 6987
rect 13001 6953 13035 6987
rect 13369 6953 13403 6987
rect 15715 6953 15749 6987
rect 18153 6953 18187 6987
rect 18521 6953 18555 6987
rect 19901 6953 19935 6987
rect 2421 6885 2455 6919
rect 4261 6885 4295 6919
rect 6009 6885 6043 6919
rect 6561 6885 6595 6919
rect 8769 6885 8803 6919
rect 13829 6885 13863 6919
rect 14381 6885 14415 6919
rect 16129 6885 16163 6919
rect 16405 6885 16439 6919
rect 16910 6885 16944 6919
rect 19257 6885 19291 6919
rect 21097 6885 21131 6919
rect 21649 6885 21683 6919
rect 1444 6817 1478 6851
rect 1547 6817 1581 6851
rect 2237 6817 2271 6851
rect 3065 6817 3099 6851
rect 8677 6817 8711 6851
rect 9689 6817 9723 6851
rect 10333 6817 10367 6851
rect 11253 6817 11287 6851
rect 11713 6817 11747 6851
rect 15577 6817 15611 6851
rect 16589 6817 16623 6851
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 5917 6749 5951 6783
rect 11989 6749 12023 6783
rect 13737 6749 13771 6783
rect 18981 6749 19015 6783
rect 21005 6749 21039 6783
rect 6837 6613 6871 6647
rect 7389 6613 7423 6647
rect 17509 6613 17543 6647
rect 18797 6613 18831 6647
rect 1547 6409 1581 6443
rect 1961 6409 1995 6443
rect 2329 6409 2363 6443
rect 2973 6409 3007 6443
rect 3571 6409 3605 6443
rect 4261 6409 4295 6443
rect 4721 6409 4755 6443
rect 7113 6409 7147 6443
rect 8401 6409 8435 6443
rect 10333 6409 10367 6443
rect 11805 6409 11839 6443
rect 12173 6409 12207 6443
rect 13369 6409 13403 6443
rect 14013 6409 14047 6443
rect 17141 6409 17175 6443
rect 7389 6341 7423 6375
rect 10517 6341 10551 6375
rect 10609 6341 10643 6375
rect 16405 6341 16439 6375
rect 19073 6341 19107 6375
rect 2421 6273 2455 6307
rect 5917 6273 5951 6307
rect 6193 6273 6227 6307
rect 6653 6273 6687 6307
rect 12449 6273 12483 6307
rect 14289 6273 14323 6307
rect 14657 6273 14691 6307
rect 15853 6273 15887 6307
rect 18797 6273 18831 6307
rect 1476 6205 1510 6239
rect 3500 6205 3534 6239
rect 5089 6205 5123 6239
rect 5273 6205 5307 6239
rect 7297 6205 7331 6239
rect 7573 6205 7607 6239
rect 9229 6205 9263 6239
rect 9781 6205 9815 6239
rect 10517 6205 10551 6239
rect 10793 6205 10827 6239
rect 11253 6205 11287 6239
rect 18153 6205 18187 6239
rect 18613 6205 18647 6239
rect 9965 6137 9999 6171
rect 11529 6137 11563 6171
rect 12771 6137 12805 6171
rect 14381 6137 14415 6171
rect 15209 6137 15243 6171
rect 15945 6137 15979 6171
rect 17785 6137 17819 6171
rect 19441 6341 19475 6375
rect 19533 6341 19567 6375
rect 20637 6341 20671 6375
rect 22477 6341 22511 6375
rect 20913 6273 20947 6307
rect 19717 6205 19751 6239
rect 21465 6205 21499 6239
rect 21925 6205 21959 6239
rect 19441 6137 19475 6171
rect 20038 6137 20072 6171
rect 3985 6069 4019 6103
rect 7757 6069 7791 6103
rect 9045 6069 9079 6103
rect 13645 6069 13679 6103
rect 15577 6069 15611 6103
rect 16773 6069 16807 6103
rect 19073 6069 19107 6103
rect 19165 6069 19199 6103
rect 21557 6069 21591 6103
rect 2559 5865 2593 5899
rect 4353 5865 4387 5899
rect 5365 5865 5399 5899
rect 9321 5865 9355 5899
rect 10103 5865 10137 5899
rect 10885 5865 10919 5899
rect 12449 5865 12483 5899
rect 18153 5865 18187 5899
rect 19901 5865 19935 5899
rect 11523 5797 11557 5831
rect 13230 5797 13264 5831
rect 15485 5797 15519 5831
rect 17325 5797 17359 5831
rect 17877 5797 17911 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 1476 5729 1510 5763
rect 2488 5729 2522 5763
rect 5549 5729 5583 5763
rect 7849 5729 7883 5763
rect 10032 5729 10066 5763
rect 11161 5729 11195 5763
rect 12909 5729 12943 5763
rect 18797 5729 18831 5763
rect 19257 5729 19291 5763
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 17233 5661 17267 5695
rect 19533 5661 19567 5695
rect 21005 5661 21039 5695
rect 1547 5593 1581 5627
rect 12081 5593 12115 5627
rect 14105 5593 14139 5627
rect 7297 5525 7331 5559
rect 8125 5525 8159 5559
rect 13829 5525 13863 5559
rect 14473 5525 14507 5559
rect 16313 5525 16347 5559
rect 20729 5525 20763 5559
rect 1547 5321 1581 5355
rect 2237 5321 2271 5355
rect 2697 5321 2731 5355
rect 4997 5321 5031 5355
rect 9137 5321 9171 5355
rect 11897 5321 11931 5355
rect 12725 5321 12759 5355
rect 13047 5321 13081 5355
rect 15669 5321 15703 5355
rect 19073 5321 19107 5355
rect 19533 5321 19567 5355
rect 20637 5321 20671 5355
rect 21005 5321 21039 5355
rect 7205 5253 7239 5287
rect 7573 5253 7607 5287
rect 8125 5253 8159 5287
rect 13737 5253 13771 5287
rect 22477 5253 22511 5287
rect 7941 5185 7975 5219
rect 8769 5185 8803 5219
rect 10057 5185 10091 5219
rect 14013 5185 14047 5219
rect 14933 5185 14967 5219
rect 15393 5185 15427 5219
rect 19717 5185 19751 5219
rect 21833 5185 21867 5219
rect 1476 5117 1510 5151
rect 1869 5117 1903 5151
rect 8033 5117 8067 5151
rect 8309 5117 8343 5151
rect 12976 5117 13010 5151
rect 13369 5117 13403 5151
rect 14657 5117 14691 5151
rect 16221 5117 16255 5151
rect 10885 5049 10919 5083
rect 10977 5049 11011 5083
rect 11529 5049 11563 5083
rect 14105 5049 14139 5083
rect 16542 5049 16576 5083
rect 17877 5049 17911 5083
rect 18153 5049 18187 5083
rect 18245 5049 18279 5083
rect 18797 5049 18831 5083
rect 20038 5049 20072 5083
rect 21557 5049 21591 5083
rect 21649 5049 21683 5083
rect 10701 4981 10735 5015
rect 16037 4981 16071 5015
rect 17141 4981 17175 5015
rect 17417 4981 17451 5015
rect 21373 4981 21407 5015
rect 1547 4777 1581 4811
rect 10149 4777 10183 4811
rect 10885 4777 10919 4811
rect 11161 4777 11195 4811
rect 12265 4777 12299 4811
rect 14197 4777 14231 4811
rect 15577 4777 15611 4811
rect 15853 4777 15887 4811
rect 17785 4777 17819 4811
rect 19257 4777 19291 4811
rect 20177 4777 20211 4811
rect 11707 4709 11741 4743
rect 13277 4709 13311 4743
rect 16589 4709 16623 4743
rect 18331 4709 18365 4743
rect 1409 4641 1443 4675
rect 8309 4641 8343 4675
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 15209 4641 15243 4675
rect 17969 4641 18003 4675
rect 19752 4641 19786 4675
rect 19855 4641 19889 4675
rect 21465 4641 21499 4675
rect 11345 4573 11379 4607
rect 13185 4573 13219 4607
rect 13461 4573 13495 4607
rect 16497 4573 16531 4607
rect 17141 4573 17175 4607
rect 9781 4505 9815 4539
rect 7941 4437 7975 4471
rect 16313 4437 16347 4471
rect 17417 4437 17451 4471
rect 18889 4437 18923 4471
rect 21097 4437 21131 4471
rect 1593 4233 1627 4267
rect 7573 4233 7607 4267
rect 10701 4233 10735 4267
rect 11897 4233 11931 4267
rect 12817 4233 12851 4267
rect 13093 4233 13127 4267
rect 15393 4233 15427 4267
rect 16773 4233 16807 4267
rect 17417 4233 17451 4267
rect 17877 4233 17911 4267
rect 19073 4233 19107 4267
rect 9781 4165 9815 4199
rect 14381 4165 14415 4199
rect 20177 4165 20211 4199
rect 8493 4097 8527 4131
rect 10057 4097 10091 4131
rect 13461 4097 13495 4131
rect 13737 4097 13771 4131
rect 16313 4097 16347 4131
rect 19533 4097 19567 4131
rect 20821 4097 20855 4131
rect 7757 4029 7791 4063
rect 7849 4029 7883 4063
rect 8033 4029 8067 4063
rect 8769 4029 8803 4063
rect 9321 4029 9355 4063
rect 10793 4029 10827 4063
rect 11253 4029 11287 4063
rect 15761 4029 15795 4063
rect 16221 4029 16255 4063
rect 18096 4029 18130 4063
rect 11529 3961 11563 3995
rect 12173 3961 12207 3995
rect 13553 3961 13587 3995
rect 18521 3961 18555 3995
rect 19257 3961 19291 3995
rect 19349 3961 19383 3995
rect 20913 3961 20947 3995
rect 21465 3961 21499 3995
rect 7297 3893 7331 3927
rect 18199 3893 18233 3927
rect 20637 3893 20671 3927
rect 10885 3689 10919 3723
rect 13645 3689 13679 3723
rect 15761 3689 15795 3723
rect 18935 3689 18969 3723
rect 19257 3689 19291 3723
rect 21097 3689 21131 3723
rect 3111 3621 3145 3655
rect 8769 3621 8803 3655
rect 13461 3621 13495 3655
rect 15439 3621 15473 3655
rect 16405 3621 16439 3655
rect 17325 3621 17359 3655
rect 3008 3553 3042 3587
rect 8033 3553 8067 3587
rect 8309 3553 8343 3587
rect 12700 3553 12734 3587
rect 15209 3553 15243 3587
rect 20821 3553 20855 3587
rect 17233 3485 17267 3519
rect 17509 3485 17543 3519
rect 7757 3417 7791 3451
rect 8125 3417 8159 3451
rect 12771 3349 12805 3383
rect 18705 3349 18739 3383
rect 8033 3145 8067 3179
rect 10149 3145 10183 3179
rect 13093 3145 13127 3179
rect 13783 3145 13817 3179
rect 15393 3145 15427 3179
rect 17233 3145 17267 3179
rect 20407 3145 20441 3179
rect 21005 3145 21039 3179
rect 23903 3145 23937 3179
rect 7297 3077 7331 3111
rect 8217 3077 8251 3111
rect 9137 3077 9171 3111
rect 8861 3009 8895 3043
rect 17509 3009 17543 3043
rect 18061 3009 18095 3043
rect 8125 2941 8159 2975
rect 8401 2941 8435 2975
rect 9756 2941 9790 2975
rect 12265 2941 12299 2975
rect 12449 2941 12483 2975
rect 13680 2941 13714 2975
rect 20177 2941 20211 2975
rect 20336 2941 20370 2975
rect 23832 2941 23866 2975
rect 3065 2805 3099 2839
rect 7573 2805 7607 2839
rect 9827 2805 9861 2839
rect 12633 2805 12667 2839
rect 14197 2805 14231 2839
rect 18797 2805 18831 2839
rect 24317 2805 24351 2839
rect 8125 2601 8159 2635
rect 10011 2601 10045 2635
rect 19763 2601 19797 2635
rect 21511 2601 21545 2635
rect 22799 2601 22833 2635
rect 9045 2533 9079 2567
rect 24179 2533 24213 2567
rect 7849 2465 7883 2499
rect 8401 2465 8435 2499
rect 9940 2465 9974 2499
rect 13553 2465 13587 2499
rect 19692 2465 19726 2499
rect 21440 2465 21474 2499
rect 22728 2465 22762 2499
rect 23121 2465 23155 2499
rect 24092 2465 24126 2499
rect 8585 2329 8619 2363
rect 13737 2329 13771 2363
rect 10425 2261 10459 2295
rect 14197 2261 14231 2295
rect 20085 2261 20119 2295
rect 21925 2261 21959 2295
rect 24593 2261 24627 2295
<< metal1 >>
rect 19242 27480 19248 27532
rect 19300 27520 19306 27532
rect 19886 27520 19892 27532
rect 19300 27492 19892 27520
rect 19300 27480 19306 27492
rect 19886 27480 19892 27492
rect 19944 27480 19950 27532
rect 24854 27480 24860 27532
rect 24912 27520 24918 27532
rect 25774 27520 25780 27532
rect 24912 27492 25780 27520
rect 24912 27480 24918 27492
rect 25774 27480 25780 27492
rect 25832 27480 25838 27532
rect 26234 27480 26240 27532
rect 26292 27520 26298 27532
rect 27246 27520 27252 27532
rect 26292 27492 27252 27520
rect 26292 27480 26298 27492
rect 27246 27480 27252 27492
rect 27304 27480 27310 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 19058 24596 19064 24608
rect 15528 24568 19064 24596
rect 15528 24556 15534 24568
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 21244 24259 21302 24265
rect 21244 24225 21256 24259
rect 21290 24256 21302 24259
rect 21358 24256 21364 24268
rect 21290 24228 21364 24256
rect 21290 24225 21302 24228
rect 21244 24219 21302 24225
rect 21358 24216 21364 24228
rect 21416 24216 21422 24268
rect 21315 24055 21373 24061
rect 21315 24021 21327 24055
rect 21361 24052 21373 24055
rect 21542 24052 21548 24064
rect 21361 24024 21548 24052
rect 21361 24021 21373 24024
rect 21315 24015 21373 24021
rect 21542 24012 21548 24024
rect 21600 24012 21606 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 8757 23851 8815 23857
rect 8757 23817 8769 23851
rect 8803 23848 8815 23851
rect 11054 23848 11060 23860
rect 8803 23820 11060 23848
rect 8803 23817 8815 23820
rect 8757 23811 8815 23817
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 12618 23848 12624 23860
rect 12579 23820 12624 23848
rect 12618 23808 12624 23820
rect 12676 23808 12682 23860
rect 13722 23848 13728 23860
rect 13683 23820 13728 23848
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 21082 23848 21088 23860
rect 19383 23820 21088 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 21358 23808 21364 23860
rect 21416 23848 21422 23860
rect 21545 23851 21603 23857
rect 21545 23848 21557 23851
rect 21416 23820 21557 23848
rect 21416 23808 21422 23820
rect 21545 23817 21557 23820
rect 21591 23817 21603 23851
rect 22554 23848 22560 23860
rect 22515 23820 22560 23848
rect 21545 23811 21603 23817
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 21269 23783 21327 23789
rect 21269 23749 21281 23783
rect 21315 23780 21327 23783
rect 22002 23780 22008 23792
rect 21315 23752 22008 23780
rect 21315 23749 21327 23752
rect 21269 23743 21327 23749
rect 1118 23672 1124 23724
rect 1176 23712 1182 23724
rect 1857 23715 1915 23721
rect 1857 23712 1869 23715
rect 1176 23684 1869 23712
rect 1176 23672 1182 23684
rect 1479 23653 1507 23684
rect 1857 23681 1869 23684
rect 1903 23681 1915 23715
rect 1857 23675 1915 23681
rect 1464 23647 1522 23653
rect 1464 23613 1476 23647
rect 1510 23613 1522 23647
rect 1464 23607 1522 23613
rect 6086 23604 6092 23656
rect 6144 23644 6150 23656
rect 8573 23647 8631 23653
rect 8573 23644 8585 23647
rect 6144 23616 8585 23644
rect 6144 23604 6150 23616
rect 8573 23613 8585 23616
rect 8619 23644 8631 23647
rect 9125 23647 9183 23653
rect 9125 23644 9137 23647
rect 8619 23616 9137 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 9125 23613 9137 23616
rect 9171 23613 9183 23647
rect 9125 23607 9183 23613
rect 11514 23604 11520 23656
rect 11572 23644 11578 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 11572 23616 12449 23644
rect 11572 23604 11578 23616
rect 12437 23613 12449 23616
rect 12483 23644 12495 23647
rect 12989 23647 13047 23653
rect 12989 23644 13001 23647
rect 12483 23616 13001 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12989 23613 13001 23616
rect 13035 23613 13047 23647
rect 13538 23644 13544 23656
rect 13451 23616 13544 23644
rect 12989 23607 13047 23613
rect 13538 23604 13544 23616
rect 13596 23644 13602 23656
rect 14093 23647 14151 23653
rect 14093 23644 14105 23647
rect 13596 23616 14105 23644
rect 13596 23604 13602 23616
rect 14093 23613 14105 23616
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 19058 23604 19064 23656
rect 19116 23644 19122 23656
rect 19153 23647 19211 23653
rect 19153 23644 19165 23647
rect 19116 23616 19165 23644
rect 19116 23604 19122 23616
rect 19153 23613 19165 23616
rect 19199 23644 19211 23647
rect 19705 23647 19763 23653
rect 19705 23644 19717 23647
rect 19199 23616 19717 23644
rect 19199 23613 19211 23616
rect 19153 23607 19211 23613
rect 19705 23613 19717 23616
rect 19751 23613 19763 23647
rect 19705 23607 19763 23613
rect 20625 23647 20683 23653
rect 20625 23613 20637 23647
rect 20671 23644 20683 23647
rect 21284 23644 21312 23743
rect 22002 23740 22008 23752
rect 22060 23740 22066 23792
rect 20671 23616 21312 23644
rect 22056 23647 22114 23653
rect 20671 23613 20683 23616
rect 20625 23607 20683 23613
rect 22056 23613 22068 23647
rect 22102 23644 22114 23647
rect 22554 23644 22560 23656
rect 22102 23616 22560 23644
rect 22102 23613 22114 23616
rect 22056 23607 22114 23613
rect 22554 23604 22560 23616
rect 22612 23604 22618 23656
rect 21266 23536 21272 23588
rect 21324 23576 21330 23588
rect 22143 23579 22201 23585
rect 22143 23576 22155 23579
rect 21324 23548 22155 23576
rect 21324 23536 21330 23548
rect 22143 23545 22155 23548
rect 22189 23545 22201 23579
rect 22143 23539 22201 23545
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1762 23508 1768 23520
rect 1581 23480 1768 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1762 23468 1768 23480
rect 1820 23468 1826 23520
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23508 20867 23511
rect 22830 23508 22836 23520
rect 20855 23480 22836 23508
rect 20855 23477 20867 23480
rect 20809 23471 20867 23477
rect 22830 23468 22836 23480
rect 22888 23468 22894 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 106 23264 112 23316
rect 164 23304 170 23316
rect 1581 23307 1639 23313
rect 1581 23304 1593 23307
rect 164 23276 1593 23304
rect 164 23264 170 23276
rect 1581 23273 1593 23276
rect 1627 23273 1639 23307
rect 1581 23267 1639 23273
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 1670 23168 1676 23180
rect 1443 23140 1676 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 1670 23128 1676 23140
rect 1728 23128 1734 23180
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 12894 22760 12900 22772
rect 12855 22732 12900 22760
rect 12894 22720 12900 22732
rect 12952 22720 12958 22772
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 15746 22760 15752 22772
rect 13403 22732 15752 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 1670 22624 1676 22636
rect 1631 22596 1676 22624
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22556 12771 22559
rect 13372 22556 13400 22723
rect 15746 22720 15752 22732
rect 15804 22760 15810 22772
rect 16942 22760 16948 22772
rect 15804 22732 16948 22760
rect 15804 22720 15810 22732
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 12759 22528 13400 22556
rect 18116 22559 18174 22565
rect 12759 22525 12771 22528
rect 12713 22519 12771 22525
rect 18116 22525 18128 22559
rect 18162 22556 18174 22559
rect 18162 22528 18644 22556
rect 18162 22525 18174 22528
rect 18116 22519 18174 22525
rect 18616 22432 18644 22528
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18187 22423 18245 22429
rect 18187 22420 18199 22423
rect 18104 22392 18199 22420
rect 18104 22380 18110 22392
rect 18187 22389 18199 22392
rect 18233 22389 18245 22423
rect 18598 22420 18604 22432
rect 18559 22392 18604 22420
rect 18187 22383 18245 22389
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 6892 20383 6950 20389
rect 6892 20349 6904 20383
rect 6938 20380 6950 20383
rect 6938 20352 7420 20380
rect 6938 20349 6950 20352
rect 6892 20343 6950 20349
rect 6963 20247 7021 20253
rect 6963 20213 6975 20247
rect 7009 20244 7021 20247
rect 7098 20244 7104 20256
rect 7009 20216 7104 20244
rect 7009 20213 7021 20216
rect 6963 20207 7021 20213
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 7392 20253 7420 20352
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 8662 20244 8668 20256
rect 7423 20216 8668 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 8662 20204 8668 20216
rect 8720 20204 8726 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 12391 20043 12449 20049
rect 12391 20009 12403 20043
rect 12437 20040 12449 20043
rect 13538 20040 13544 20052
rect 12437 20012 13544 20040
rect 12437 20009 12449 20012
rect 12391 20003 12449 20009
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 5166 19864 5172 19916
rect 5224 19904 5230 19916
rect 6549 19907 6607 19913
rect 6549 19904 6561 19907
rect 5224 19876 6561 19904
rect 5224 19864 5230 19876
rect 6549 19873 6561 19876
rect 6595 19904 6607 19907
rect 6638 19904 6644 19916
rect 6595 19876 6644 19904
rect 6595 19873 6607 19876
rect 6549 19867 6607 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 12320 19907 12378 19913
rect 12320 19873 12332 19907
rect 12366 19904 12378 19907
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 12366 19876 12725 19904
rect 12366 19873 12378 19876
rect 12320 19867 12378 19873
rect 12713 19873 12725 19876
rect 12759 19904 12771 19907
rect 13170 19904 13176 19916
rect 12759 19876 13176 19904
rect 12759 19873 12771 19876
rect 12713 19867 12771 19873
rect 13170 19864 13176 19876
rect 13228 19864 13234 19916
rect 8478 19768 8484 19780
rect 8439 19740 8484 19768
rect 8478 19728 8484 19740
rect 8536 19728 8542 19780
rect 6687 19703 6745 19709
rect 6687 19669 6699 19703
rect 6733 19700 6745 19703
rect 7190 19700 7196 19712
rect 6733 19672 7196 19700
rect 6733 19669 6745 19672
rect 6687 19663 6745 19669
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 7834 19660 7840 19712
rect 7892 19700 7898 19712
rect 8711 19703 8769 19709
rect 8711 19700 8723 19703
rect 7892 19672 8723 19700
rect 7892 19660 7898 19672
rect 8711 19669 8723 19672
rect 8757 19669 8769 19703
rect 8711 19663 8769 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1578 19496 1584 19508
rect 1539 19468 1584 19496
rect 1578 19456 1584 19468
rect 1636 19456 1642 19508
rect 3878 19496 3884 19508
rect 3839 19468 3884 19496
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 5859 19499 5917 19505
rect 5859 19465 5871 19499
rect 5905 19496 5917 19499
rect 6086 19496 6092 19508
rect 5905 19468 6092 19496
rect 5905 19465 5917 19468
rect 5859 19459 5917 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 7834 19496 7840 19508
rect 7795 19468 7840 19496
rect 7834 19456 7840 19468
rect 7892 19456 7898 19508
rect 9582 19496 9588 19508
rect 9543 19468 9588 19496
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 25130 19496 25136 19508
rect 25091 19468 25136 19496
rect 25130 19456 25136 19468
rect 25188 19456 25194 19508
rect 7650 19360 7656 19372
rect 4126 19332 7656 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 3472 19295 3530 19301
rect 1443 19264 2084 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 2056 19165 2084 19264
rect 3472 19261 3484 19295
rect 3518 19292 3530 19295
rect 3878 19292 3884 19304
rect 3518 19264 3884 19292
rect 3518 19261 3530 19264
rect 3472 19255 3530 19261
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 3559 19227 3617 19233
rect 3559 19193 3571 19227
rect 3605 19224 3617 19227
rect 4126 19224 4154 19332
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8628 19332 11411 19360
rect 8628 19320 8634 19332
rect 5788 19295 5846 19301
rect 5788 19261 5800 19295
rect 5834 19292 5846 19295
rect 5834 19264 6316 19292
rect 5834 19261 5846 19264
rect 5788 19255 5846 19261
rect 3605 19196 4154 19224
rect 3605 19193 3617 19196
rect 3559 19187 3617 19193
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2498 19156 2504 19168
rect 2087 19128 2504 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2498 19116 2504 19128
rect 2556 19116 2562 19168
rect 6288 19165 6316 19264
rect 7834 19252 7840 19304
rect 7892 19292 7898 19304
rect 7929 19295 7987 19301
rect 7929 19292 7941 19295
rect 7892 19264 7941 19292
rect 7892 19252 7898 19264
rect 7929 19261 7941 19264
rect 7975 19261 7987 19295
rect 7929 19255 7987 19261
rect 9100 19295 9158 19301
rect 9100 19261 9112 19295
rect 9146 19292 9158 19295
rect 9582 19292 9588 19304
rect 9146 19264 9588 19292
rect 9146 19261 9158 19264
rect 9100 19255 9158 19261
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 11383 19301 11411 19332
rect 11368 19295 11426 19301
rect 11368 19261 11380 19295
rect 11414 19292 11426 19295
rect 11790 19292 11796 19304
rect 11414 19264 11796 19292
rect 11414 19261 11426 19264
rect 11368 19255 11426 19261
rect 11790 19252 11796 19264
rect 11848 19252 11854 19304
rect 12529 19295 12587 19301
rect 12529 19292 12541 19295
rect 12360 19264 12541 19292
rect 8478 19184 8484 19236
rect 8536 19224 8542 19236
rect 8665 19227 8723 19233
rect 8665 19224 8677 19227
rect 8536 19196 8677 19224
rect 8536 19184 8542 19196
rect 8665 19193 8677 19196
rect 8711 19224 8723 19227
rect 9858 19224 9864 19236
rect 8711 19196 9864 19224
rect 8711 19193 8723 19196
rect 8665 19187 8723 19193
rect 9858 19184 9864 19196
rect 9916 19184 9922 19236
rect 12360 19168 12388 19264
rect 12529 19261 12541 19264
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 24648 19295 24706 19301
rect 24648 19261 24660 19295
rect 24694 19292 24706 19295
rect 25130 19292 25136 19304
rect 24694 19264 25136 19292
rect 24694 19261 24706 19264
rect 24648 19255 24706 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 6273 19159 6331 19165
rect 6273 19125 6285 19159
rect 6319 19156 6331 19159
rect 6454 19156 6460 19168
rect 6319 19128 6460 19156
rect 6319 19125 6331 19128
rect 6273 19119 6331 19125
rect 6454 19116 6460 19128
rect 6512 19116 6518 19168
rect 6638 19156 6644 19168
rect 6599 19128 6644 19156
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 6914 19156 6920 19168
rect 6875 19128 6920 19156
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 8113 19159 8171 19165
rect 8113 19156 8125 19159
rect 7064 19128 8125 19156
rect 7064 19116 7070 19128
rect 8113 19125 8125 19128
rect 8159 19125 8171 19159
rect 8113 19119 8171 19125
rect 8938 19116 8944 19168
rect 8996 19156 9002 19168
rect 9171 19159 9229 19165
rect 9171 19156 9183 19159
rect 8996 19128 9183 19156
rect 8996 19116 9002 19128
rect 9171 19125 9183 19128
rect 9217 19125 9229 19159
rect 9171 19119 9229 19125
rect 11471 19159 11529 19165
rect 11471 19125 11483 19159
rect 11517 19156 11529 19159
rect 11698 19156 11704 19168
rect 11517 19128 11704 19156
rect 11517 19125 11529 19128
rect 11471 19119 11529 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12342 19156 12348 19168
rect 12299 19128 12348 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 12342 19116 12348 19128
rect 12400 19116 12406 19168
rect 12710 19156 12716 19168
rect 12671 19128 12716 19156
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 16758 19116 16764 19168
rect 16816 19156 16822 19168
rect 24719 19159 24777 19165
rect 24719 19156 24731 19159
rect 16816 19128 24731 19156
rect 16816 19116 16822 19128
rect 24719 19125 24731 19128
rect 24765 19125 24777 19159
rect 24719 19119 24777 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1486 18912 1492 18964
rect 1544 18952 1550 18964
rect 1581 18955 1639 18961
rect 1581 18952 1593 18955
rect 1544 18924 1593 18952
rect 1544 18912 1550 18924
rect 1581 18921 1593 18924
rect 1627 18921 1639 18955
rect 7006 18952 7012 18964
rect 1581 18915 1639 18921
rect 4126 18924 7012 18952
rect 106 18844 112 18896
rect 164 18884 170 18896
rect 4126 18884 4154 18924
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7190 18952 7196 18964
rect 7151 18924 7196 18952
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 6362 18884 6368 18896
rect 164 18856 4154 18884
rect 6323 18856 6368 18884
rect 164 18844 170 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 7650 18844 7656 18896
rect 7708 18884 7714 18896
rect 7834 18884 7840 18896
rect 7708 18856 7840 18884
rect 7708 18844 7714 18856
rect 7834 18844 7840 18856
rect 7892 18844 7898 18896
rect 7926 18844 7932 18896
rect 7984 18884 7990 18896
rect 9861 18887 9919 18893
rect 7984 18856 8029 18884
rect 7984 18844 7990 18856
rect 9861 18853 9873 18887
rect 9907 18884 9919 18887
rect 10134 18884 10140 18896
rect 9907 18856 10140 18884
rect 9907 18853 9919 18856
rect 9861 18847 9919 18853
rect 10134 18844 10140 18856
rect 10192 18844 10198 18896
rect 11698 18844 11704 18896
rect 11756 18884 11762 18896
rect 12250 18884 12256 18896
rect 11756 18856 12256 18884
rect 11756 18844 11762 18856
rect 12250 18844 12256 18856
rect 12308 18844 12314 18896
rect 12345 18887 12403 18893
rect 12345 18853 12357 18887
rect 12391 18884 12403 18887
rect 12434 18884 12440 18896
rect 12391 18856 12440 18884
rect 12391 18853 12403 18856
rect 12345 18847 12403 18853
rect 12434 18844 12440 18856
rect 12492 18844 12498 18896
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 1946 18816 1952 18828
rect 1903 18788 1952 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 1946 18776 1952 18788
rect 2004 18776 2010 18828
rect 5052 18819 5110 18825
rect 5052 18785 5064 18819
rect 5098 18816 5110 18819
rect 5166 18816 5172 18828
rect 5098 18788 5172 18816
rect 5098 18785 5110 18788
rect 5052 18779 5110 18785
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 13792 18819 13850 18825
rect 13792 18785 13804 18819
rect 13838 18816 13850 18819
rect 13906 18816 13912 18828
rect 13838 18788 13912 18816
rect 13838 18785 13850 18788
rect 13792 18779 13850 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 18760 18819 18818 18825
rect 18760 18785 18772 18819
rect 18806 18816 18818 18819
rect 19334 18816 19340 18828
rect 18806 18788 19340 18816
rect 18806 18785 18818 18788
rect 18760 18779 18818 18785
rect 19334 18776 19340 18788
rect 19392 18816 19398 18828
rect 24210 18816 24216 18828
rect 19392 18788 24216 18816
rect 19392 18776 19398 18788
rect 24210 18776 24216 18788
rect 24268 18776 24274 18828
rect 2087 18751 2145 18757
rect 2087 18717 2099 18751
rect 2133 18748 2145 18751
rect 6270 18748 6276 18760
rect 2133 18720 6276 18748
rect 2133 18717 2145 18720
rect 2087 18711 2145 18717
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 8478 18748 8484 18760
rect 8439 18720 8484 18748
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 9766 18748 9772 18760
rect 9727 18720 9772 18748
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 9858 18708 9864 18760
rect 9916 18748 9922 18760
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 9916 18720 10425 18748
rect 9916 18708 9922 18720
rect 10413 18717 10425 18720
rect 10459 18748 10471 18751
rect 10962 18748 10968 18760
rect 10459 18720 10968 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 10962 18708 10968 18720
rect 11020 18708 11026 18760
rect 17678 18748 17684 18760
rect 17639 18720 17684 18748
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 6825 18683 6883 18689
rect 6825 18649 6837 18683
rect 6871 18680 6883 18683
rect 8496 18680 8524 18708
rect 12802 18680 12808 18692
rect 6871 18652 8524 18680
rect 12763 18652 12808 18680
rect 6871 18649 6883 18652
rect 6825 18643 6883 18649
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 5123 18615 5181 18621
rect 5123 18612 5135 18615
rect 4856 18584 5135 18612
rect 4856 18572 4862 18584
rect 5123 18581 5135 18584
rect 5169 18581 5181 18615
rect 5123 18575 5181 18581
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 8294 18612 8300 18624
rect 7800 18584 8300 18612
rect 7800 18572 7806 18584
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 13863 18615 13921 18621
rect 13863 18612 13875 18615
rect 12584 18584 13875 18612
rect 12584 18572 12590 18584
rect 13863 18581 13875 18584
rect 13909 18581 13921 18615
rect 13863 18575 13921 18581
rect 18831 18615 18889 18621
rect 18831 18581 18843 18615
rect 18877 18612 18889 18615
rect 19886 18612 19892 18624
rect 18877 18584 19892 18612
rect 18877 18581 18889 18584
rect 18831 18575 18889 18581
rect 19886 18572 19892 18584
rect 19944 18572 19950 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 5166 18408 5172 18420
rect 5127 18380 5172 18408
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 6362 18368 6368 18420
rect 6420 18408 6426 18420
rect 6546 18408 6552 18420
rect 6420 18380 6552 18408
rect 6420 18368 6426 18380
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 12710 18408 12716 18420
rect 12671 18380 12716 18408
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13906 18408 13912 18420
rect 13819 18380 13912 18408
rect 13906 18368 13912 18380
rect 13964 18408 13970 18420
rect 19334 18408 19340 18420
rect 13964 18380 19340 18408
rect 13964 18368 13970 18380
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 24762 18408 24768 18420
rect 24723 18380 24768 18408
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 5859 18343 5917 18349
rect 5859 18309 5871 18343
rect 5905 18340 5917 18343
rect 7558 18340 7564 18352
rect 5905 18312 7564 18340
rect 5905 18309 5917 18312
rect 5859 18303 5917 18309
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 7742 18300 7748 18352
rect 7800 18340 7806 18352
rect 9766 18340 9772 18352
rect 7800 18312 9772 18340
rect 7800 18300 7806 18312
rect 7101 18275 7159 18281
rect 7101 18241 7113 18275
rect 7147 18272 7159 18275
rect 7190 18272 7196 18284
rect 7147 18244 7196 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 8938 18272 8944 18284
rect 8899 18244 8944 18272
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9232 18281 9260 18312
rect 9766 18300 9772 18312
rect 9824 18340 9830 18352
rect 10229 18343 10287 18349
rect 10229 18340 10241 18343
rect 9824 18312 10241 18340
rect 9824 18300 9830 18312
rect 10229 18309 10241 18312
rect 10275 18309 10287 18343
rect 10229 18303 10287 18309
rect 10551 18343 10609 18349
rect 10551 18309 10563 18343
rect 10597 18340 10609 18343
rect 17034 18340 17040 18352
rect 10597 18312 17040 18340
rect 10597 18309 10609 18312
rect 10551 18303 10609 18309
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 18877 18343 18935 18349
rect 18877 18309 18889 18343
rect 18923 18340 18935 18343
rect 18923 18312 20208 18340
rect 18923 18309 18935 18312
rect 18877 18303 18935 18309
rect 20180 18284 20208 18312
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10873 18275 10931 18281
rect 10873 18272 10885 18275
rect 9640 18244 10885 18272
rect 9640 18232 9646 18244
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 1486 18204 1492 18216
rect 1443 18176 1492 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1486 18164 1492 18176
rect 1544 18164 1550 18216
rect 10463 18213 10491 18244
rect 10873 18241 10885 18244
rect 10919 18241 10931 18275
rect 13170 18272 13176 18284
rect 13131 18244 13176 18272
rect 10873 18235 10931 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 17494 18232 17500 18284
rect 17552 18272 17558 18284
rect 19886 18272 19892 18284
rect 17552 18244 19334 18272
rect 19847 18244 19892 18272
rect 17552 18232 17558 18244
rect 5788 18207 5846 18213
rect 5788 18204 5800 18207
rect 4126 18176 5800 18204
rect 3326 18096 3332 18148
rect 3384 18136 3390 18148
rect 4126 18136 4154 18176
rect 5788 18173 5800 18176
rect 5834 18204 5846 18207
rect 10448 18207 10506 18213
rect 5834 18176 6316 18204
rect 5834 18173 5846 18176
rect 5788 18167 5846 18173
rect 3384 18108 4154 18136
rect 3384 18096 3390 18108
rect 1535 18071 1593 18077
rect 1535 18037 1547 18071
rect 1581 18068 1593 18071
rect 1670 18068 1676 18080
rect 1581 18040 1676 18068
rect 1581 18037 1593 18040
rect 1535 18031 1593 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 4706 18068 4712 18080
rect 4667 18040 4712 18068
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 6288 18077 6316 18176
rect 10448 18173 10460 18207
rect 10494 18173 10506 18207
rect 10448 18167 10506 18173
rect 14528 18207 14586 18213
rect 14528 18173 14540 18207
rect 14574 18204 14586 18207
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14574 18176 14933 18204
rect 14574 18173 14586 18176
rect 14528 18167 14586 18173
rect 14921 18173 14933 18176
rect 14967 18204 14979 18207
rect 16298 18204 16304 18216
rect 14967 18176 16304 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 16298 18164 16304 18176
rect 16356 18164 16362 18216
rect 16574 18164 16580 18216
rect 16632 18204 16638 18216
rect 16980 18207 17038 18213
rect 16980 18204 16992 18207
rect 16632 18176 16992 18204
rect 16632 18164 16638 18176
rect 16980 18173 16992 18176
rect 17026 18204 17038 18207
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 17026 18176 17417 18204
rect 17026 18173 17038 18176
rect 16980 18167 17038 18173
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 7193 18139 7251 18145
rect 7193 18105 7205 18139
rect 7239 18136 7251 18139
rect 7374 18136 7380 18148
rect 7239 18108 7380 18136
rect 7239 18105 7251 18108
rect 7193 18099 7251 18105
rect 7374 18096 7380 18108
rect 7432 18096 7438 18148
rect 7745 18139 7803 18145
rect 7745 18105 7757 18139
rect 7791 18136 7803 18139
rect 8478 18136 8484 18148
rect 7791 18108 8484 18136
rect 7791 18105 7803 18108
rect 7745 18099 7803 18105
rect 8478 18096 8484 18108
rect 8536 18096 8542 18148
rect 8757 18139 8815 18145
rect 8757 18105 8769 18139
rect 8803 18136 8815 18139
rect 9033 18139 9091 18145
rect 9033 18136 9045 18139
rect 8803 18108 9045 18136
rect 8803 18105 8815 18108
rect 8757 18099 8815 18105
rect 9033 18105 9045 18108
rect 9079 18136 9091 18139
rect 9766 18136 9772 18148
rect 9079 18108 9772 18136
rect 9079 18105 9091 18108
rect 9033 18099 9091 18105
rect 6273 18071 6331 18077
rect 6273 18037 6285 18071
rect 6319 18068 6331 18071
rect 6362 18068 6368 18080
rect 6319 18040 6368 18068
rect 6319 18037 6331 18040
rect 6273 18031 6331 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7984 18040 8125 18068
rect 7984 18028 7990 18040
rect 8113 18037 8125 18040
rect 8159 18068 8171 18071
rect 8772 18068 8800 18099
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 11606 18096 11612 18148
rect 11664 18136 11670 18148
rect 12253 18139 12311 18145
rect 12253 18136 12265 18139
rect 11664 18108 12265 18136
rect 11664 18096 11670 18108
rect 12253 18105 12265 18108
rect 12299 18136 12311 18139
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 12299 18108 12909 18136
rect 12299 18105 12311 18108
rect 12253 18099 12311 18105
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 12989 18139 13047 18145
rect 12989 18105 13001 18139
rect 13035 18105 13047 18139
rect 12989 18099 13047 18105
rect 17083 18139 17141 18145
rect 17083 18105 17095 18139
rect 17129 18136 17141 18139
rect 18322 18136 18328 18148
rect 17129 18108 18328 18136
rect 17129 18105 17141 18108
rect 17083 18099 17141 18105
rect 8159 18040 8800 18068
rect 9953 18071 10011 18077
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 9953 18037 9965 18071
rect 9999 18068 10011 18071
rect 10134 18068 10140 18080
rect 9999 18040 10140 18068
rect 9999 18037 10011 18040
rect 9953 18031 10011 18037
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 11885 18071 11943 18077
rect 11885 18037 11897 18071
rect 11931 18068 11943 18071
rect 12434 18068 12440 18080
rect 11931 18040 12440 18068
rect 11931 18037 11943 18040
rect 11885 18031 11943 18037
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13004 18068 13032 18099
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 18426 18139 18484 18145
rect 18426 18105 18438 18139
rect 18472 18105 18484 18139
rect 19306 18136 19334 18244
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 20162 18272 20168 18284
rect 20075 18244 20168 18272
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24268 18176 24593 18204
rect 24268 18164 24274 18176
rect 24581 18173 24593 18176
rect 24627 18204 24639 18207
rect 25133 18207 25191 18213
rect 25133 18204 25145 18207
rect 24627 18176 25145 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 25133 18173 25145 18176
rect 25179 18173 25191 18207
rect 25133 18167 25191 18173
rect 19705 18139 19763 18145
rect 19705 18136 19717 18139
rect 19306 18108 19717 18136
rect 18426 18099 18484 18105
rect 19705 18105 19717 18108
rect 19751 18136 19763 18139
rect 19981 18139 20039 18145
rect 19981 18136 19993 18139
rect 19751 18108 19993 18136
rect 19751 18105 19763 18108
rect 19705 18099 19763 18105
rect 19981 18105 19993 18108
rect 20027 18136 20039 18139
rect 21358 18136 21364 18148
rect 20027 18108 21364 18136
rect 20027 18105 20039 18108
rect 19981 18099 20039 18105
rect 12768 18040 13032 18068
rect 12768 18028 12774 18040
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 14599 18071 14657 18077
rect 14599 18068 14611 18071
rect 14332 18040 14611 18068
rect 14332 18028 14338 18040
rect 14599 18037 14611 18040
rect 14645 18037 14657 18071
rect 14599 18031 14657 18037
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18230 18068 18236 18080
rect 17911 18040 18236 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 18230 18028 18236 18040
rect 18288 18068 18294 18080
rect 18432 18068 18460 18099
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 18288 18040 18460 18068
rect 18288 18028 18294 18040
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 6270 17864 6276 17876
rect 6231 17836 6276 17864
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 8205 17867 8263 17873
rect 8205 17864 8217 17867
rect 7892 17836 8217 17864
rect 7892 17824 7898 17836
rect 8205 17833 8217 17836
rect 8251 17833 8263 17867
rect 8938 17864 8944 17876
rect 8899 17836 8944 17864
rect 8205 17827 8263 17833
rect 8938 17824 8944 17836
rect 8996 17824 9002 17876
rect 11606 17864 11612 17876
rect 11567 17836 11612 17864
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 12250 17864 12256 17876
rect 12211 17836 12256 17864
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 17034 17864 17040 17876
rect 16995 17836 17040 17864
rect 17034 17824 17040 17836
rect 17092 17824 17098 17876
rect 18322 17864 18328 17876
rect 18283 17836 18328 17864
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 19889 17867 19947 17873
rect 19889 17833 19901 17867
rect 19935 17864 19947 17867
rect 19978 17864 19984 17876
rect 19935 17836 19984 17864
rect 19935 17833 19947 17836
rect 19889 17827 19947 17833
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 20162 17864 20168 17876
rect 20123 17836 20168 17864
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 21542 17864 21548 17876
rect 21503 17836 21548 17864
rect 21542 17824 21548 17836
rect 21600 17824 21606 17876
rect 24489 17867 24547 17873
rect 24489 17833 24501 17867
rect 24535 17864 24547 17867
rect 25498 17864 25504 17876
rect 24535 17836 25504 17864
rect 24535 17833 24547 17836
rect 24489 17827 24547 17833
rect 25498 17824 25504 17836
rect 25556 17824 25562 17876
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 7285 17799 7343 17805
rect 7285 17796 7297 17799
rect 6972 17768 7297 17796
rect 6972 17756 6978 17768
rect 7285 17765 7297 17768
rect 7331 17765 7343 17799
rect 7285 17759 7343 17765
rect 7374 17756 7380 17808
rect 7432 17796 7438 17808
rect 7650 17796 7656 17808
rect 7432 17768 7656 17796
rect 7432 17756 7438 17768
rect 7650 17756 7656 17768
rect 7708 17756 7714 17808
rect 9858 17796 9864 17808
rect 9819 17768 9864 17796
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 12342 17756 12348 17808
rect 12400 17796 12406 17808
rect 12805 17799 12863 17805
rect 12805 17796 12817 17799
rect 12400 17768 12817 17796
rect 12400 17756 12406 17768
rect 12805 17765 12817 17768
rect 12851 17796 12863 17799
rect 13538 17796 13544 17808
rect 12851 17768 13544 17796
rect 12851 17765 12863 17768
rect 12805 17759 12863 17765
rect 13538 17756 13544 17768
rect 13596 17756 13602 17808
rect 17052 17796 17080 17824
rect 17313 17799 17371 17805
rect 17313 17796 17325 17799
rect 17052 17768 17325 17796
rect 17313 17765 17325 17768
rect 17359 17765 17371 17799
rect 17313 17759 17371 17765
rect 17405 17799 17463 17805
rect 17405 17765 17417 17799
rect 17451 17796 17463 17799
rect 17494 17796 17500 17808
rect 17451 17768 17500 17796
rect 17451 17765 17463 17768
rect 17405 17759 17463 17765
rect 17494 17756 17500 17768
rect 17552 17756 17558 17808
rect 18414 17756 18420 17808
rect 18472 17796 18478 17808
rect 18877 17799 18935 17805
rect 18877 17796 18889 17799
rect 18472 17768 18889 17796
rect 18472 17756 18478 17768
rect 18877 17765 18889 17768
rect 18923 17765 18935 17799
rect 18877 17759 18935 17765
rect 18969 17799 19027 17805
rect 18969 17765 18981 17799
rect 19015 17796 19027 17799
rect 19150 17796 19156 17808
rect 19015 17768 19156 17796
rect 19015 17765 19027 17768
rect 18969 17759 19027 17765
rect 19150 17756 19156 17768
rect 19208 17756 19214 17808
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 2501 17731 2559 17737
rect 2501 17697 2513 17731
rect 2547 17728 2559 17731
rect 2590 17728 2596 17740
rect 2547 17700 2596 17728
rect 2547 17697 2559 17700
rect 2501 17691 2559 17697
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 5442 17728 5448 17740
rect 5403 17700 5448 17728
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 15378 17728 15384 17740
rect 15339 17700 15384 17728
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22592 17731 22650 17737
rect 22592 17728 22604 17731
rect 22520 17700 22604 17728
rect 22520 17688 22526 17700
rect 22592 17697 22604 17700
rect 22638 17697 22650 17731
rect 22592 17691 22650 17697
rect 22695 17731 22753 17737
rect 22695 17697 22707 17731
rect 22741 17728 22753 17731
rect 24210 17728 24216 17740
rect 22741 17700 24216 17728
rect 22741 17697 22753 17700
rect 22695 17691 22753 17697
rect 24210 17688 24216 17700
rect 24268 17728 24274 17740
rect 24305 17731 24363 17737
rect 24305 17728 24317 17731
rect 24268 17700 24317 17728
rect 24268 17688 24274 17700
rect 24305 17697 24317 17700
rect 24351 17697 24363 17731
rect 24305 17691 24363 17697
rect 7742 17660 7748 17672
rect 7703 17632 7748 17660
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 8536 17632 9781 17660
rect 8536 17620 8542 17632
rect 9769 17629 9781 17632
rect 9815 17660 9827 17663
rect 10594 17660 10600 17672
rect 9815 17632 10600 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 12802 17660 12808 17672
rect 12759 17632 12808 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 12802 17620 12808 17632
rect 12860 17620 12866 17672
rect 13170 17660 13176 17672
rect 13131 17632 13176 17660
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13412 17632 14197 17660
rect 13412 17620 13418 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 18506 17660 18512 17672
rect 18003 17632 18512 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 19153 17663 19211 17669
rect 19153 17629 19165 17663
rect 19199 17629 19211 17663
rect 19153 17623 19211 17629
rect 1762 17552 1768 17604
rect 1820 17592 1826 17604
rect 8202 17592 8208 17604
rect 1820 17564 8208 17592
rect 1820 17552 1826 17564
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 10321 17595 10379 17601
rect 10321 17561 10333 17595
rect 10367 17592 10379 17595
rect 10962 17592 10968 17604
rect 10367 17564 10968 17592
rect 10367 17561 10379 17564
rect 10321 17555 10379 17561
rect 10962 17552 10968 17564
rect 11020 17552 11026 17604
rect 18524 17592 18552 17620
rect 19168 17592 19196 17623
rect 18524 17564 19196 17592
rect 2639 17527 2697 17533
rect 2639 17493 2651 17527
rect 2685 17524 2697 17527
rect 3513 17527 3571 17533
rect 3513 17524 3525 17527
rect 2685 17496 3525 17524
rect 2685 17493 2697 17496
rect 2639 17487 2697 17493
rect 3513 17493 3525 17496
rect 3559 17524 3571 17527
rect 3602 17524 3608 17536
rect 3559 17496 3608 17524
rect 3559 17493 3571 17496
rect 3513 17487 3571 17493
rect 3602 17484 3608 17496
rect 3660 17484 3666 17536
rect 5074 17524 5080 17536
rect 5035 17496 5080 17524
rect 5074 17484 5080 17496
rect 5132 17484 5138 17536
rect 7101 17527 7159 17533
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7650 17524 7656 17536
rect 7147 17496 7656 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 15749 17527 15807 17533
rect 15749 17493 15761 17527
rect 15795 17524 15807 17527
rect 15930 17524 15936 17536
rect 15795 17496 15936 17524
rect 15795 17493 15807 17496
rect 15749 17487 15807 17493
rect 15930 17484 15936 17496
rect 15988 17484 15994 17536
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 18472 17496 18613 17524
rect 18472 17484 18478 17496
rect 18601 17493 18613 17496
rect 18647 17493 18659 17527
rect 18601 17487 18659 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 3326 17320 3332 17332
rect 3287 17292 3332 17320
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 4617 17323 4675 17329
rect 4617 17289 4629 17323
rect 4663 17320 4675 17323
rect 4706 17320 4712 17332
rect 4663 17292 4712 17320
rect 4663 17289 4675 17292
rect 4617 17283 4675 17289
rect 4706 17280 4712 17292
rect 4764 17280 4770 17332
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 5074 17320 5080 17332
rect 5031 17292 5080 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 6089 17323 6147 17329
rect 6089 17320 6101 17323
rect 5500 17292 6101 17320
rect 5500 17280 5506 17292
rect 6089 17289 6101 17292
rect 6135 17320 6147 17323
rect 6362 17320 6368 17332
rect 6135 17292 6368 17320
rect 6135 17289 6147 17292
rect 6089 17283 6147 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 6546 17320 6552 17332
rect 6507 17292 6552 17320
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9490 17320 9496 17332
rect 9171 17292 9496 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 9490 17280 9496 17292
rect 9548 17320 9554 17332
rect 9858 17320 9864 17332
rect 9548 17292 9864 17320
rect 9548 17280 9554 17292
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10594 17320 10600 17332
rect 10555 17292 10600 17320
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11572 17292 11621 17320
rect 11572 17280 11578 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 11609 17283 11667 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 17313 17323 17371 17329
rect 17313 17289 17325 17323
rect 17359 17320 17371 17323
rect 17494 17320 17500 17332
rect 17359 17292 17500 17320
rect 17359 17289 17371 17292
rect 17313 17283 17371 17289
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 17736 17292 17785 17320
rect 17736 17280 17742 17292
rect 17773 17289 17785 17292
rect 17819 17289 17831 17323
rect 17773 17283 17831 17289
rect 106 17144 112 17196
rect 164 17184 170 17196
rect 2590 17184 2596 17196
rect 164 17156 2596 17184
rect 164 17144 170 17156
rect 2590 17144 2596 17156
rect 2648 17184 2654 17196
rect 2869 17187 2927 17193
rect 2869 17184 2881 17187
rect 2648 17156 2881 17184
rect 2648 17144 2654 17156
rect 2869 17153 2881 17156
rect 2915 17153 2927 17187
rect 3602 17184 3608 17196
rect 3563 17156 3608 17184
rect 2869 17147 2927 17153
rect 3602 17144 3608 17156
rect 3660 17144 3666 17196
rect 4724 17184 4752 17280
rect 7098 17212 7104 17264
rect 7156 17252 7162 17264
rect 7742 17252 7748 17264
rect 7156 17224 7236 17252
rect 7703 17224 7748 17252
rect 7156 17212 7162 17224
rect 7208 17193 7236 17224
rect 7742 17212 7748 17224
rect 7800 17212 7806 17264
rect 5169 17187 5227 17193
rect 5169 17184 5181 17187
rect 4724 17156 5181 17184
rect 5169 17153 5181 17156
rect 5215 17153 5227 17187
rect 5169 17147 5227 17153
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17184 7251 17187
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7239 17156 8125 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 8113 17147 8171 17153
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12526 17184 12532 17196
rect 11931 17156 12532 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 17788 17184 17816 17283
rect 22462 17280 22468 17332
rect 22520 17320 22526 17332
rect 22557 17323 22615 17329
rect 22557 17320 22569 17323
rect 22520 17292 22569 17320
rect 22520 17280 22526 17292
rect 22557 17289 22569 17292
rect 22603 17289 22615 17323
rect 22557 17283 22615 17289
rect 24210 17280 24216 17332
rect 24268 17320 24274 17332
rect 24305 17323 24363 17329
rect 24305 17320 24317 17323
rect 24268 17292 24317 17320
rect 24268 17280 24274 17292
rect 24305 17289 24317 17292
rect 24351 17289 24363 17323
rect 24305 17283 24363 17289
rect 20530 17252 20536 17264
rect 20443 17224 20536 17252
rect 20530 17212 20536 17224
rect 20588 17252 20594 17264
rect 21726 17252 21732 17264
rect 20588 17224 21732 17252
rect 20588 17212 20594 17224
rect 21726 17212 21732 17224
rect 21784 17252 21790 17264
rect 22480 17252 22508 17280
rect 21784 17224 22508 17252
rect 21784 17212 21790 17224
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 17788 17156 18245 17184
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18506 17184 18512 17196
rect 18467 17156 18512 17184
rect 18233 17147 18291 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20162 17184 20168 17196
rect 20027 17156 20168 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 21542 17184 21548 17196
rect 21503 17156 21548 17184
rect 21542 17144 21548 17156
rect 21600 17144 21606 17196
rect 1394 17076 1400 17128
rect 1452 17116 1458 17128
rect 1949 17119 2007 17125
rect 1949 17116 1961 17119
rect 1452 17088 1961 17116
rect 1452 17076 1458 17088
rect 1949 17085 1961 17088
rect 1995 17116 2007 17119
rect 2476 17119 2534 17125
rect 2476 17116 2488 17119
rect 1995 17088 2488 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2476 17085 2488 17088
rect 2522 17116 2534 17119
rect 3326 17116 3332 17128
rect 2522 17088 3332 17116
rect 2522 17085 2534 17088
rect 2476 17079 2534 17085
rect 3326 17076 3332 17088
rect 3384 17076 3390 17128
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 11368 17119 11426 17125
rect 11368 17116 11380 17119
rect 11287 17088 11380 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 11368 17085 11380 17088
rect 11414 17116 11426 17119
rect 12342 17116 12348 17128
rect 11414 17088 12348 17116
rect 11414 17085 11426 17088
rect 11368 17079 11426 17085
rect 12342 17076 12348 17088
rect 12400 17076 12406 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13228 17088 13921 17116
rect 13228 17076 13234 17088
rect 13909 17085 13921 17088
rect 13955 17116 13967 17119
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13955 17088 14105 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 15654 17116 15660 17128
rect 15615 17088 15660 17116
rect 14093 17079 14151 17085
rect 15654 17076 15660 17088
rect 15712 17116 15718 17128
rect 16577 17119 16635 17125
rect 16577 17116 16589 17119
rect 15712 17088 16589 17116
rect 15712 17076 15718 17088
rect 16577 17085 16589 17088
rect 16623 17085 16635 17119
rect 16577 17079 16635 17085
rect 3697 17051 3755 17057
rect 3697 17017 3709 17051
rect 3743 17048 3755 17051
rect 3970 17048 3976 17060
rect 3743 17020 3976 17048
rect 3743 17017 3755 17020
rect 3697 17011 3755 17017
rect 3970 17008 3976 17020
rect 4028 17008 4034 17060
rect 4249 17051 4307 17057
rect 4249 17017 4261 17051
rect 4295 17048 4307 17051
rect 4982 17048 4988 17060
rect 4295 17020 4988 17048
rect 4295 17017 4307 17020
rect 4249 17011 4307 17017
rect 4982 17008 4988 17020
rect 5040 17008 5046 17060
rect 5261 17051 5319 17057
rect 5261 17017 5273 17051
rect 5307 17017 5319 17051
rect 5261 17011 5319 17017
rect 5813 17051 5871 17057
rect 5813 17017 5825 17051
rect 5859 17048 5871 17051
rect 6454 17048 6460 17060
rect 5859 17020 6460 17048
rect 5859 17017 5871 17020
rect 5813 17011 5871 17017
rect 1397 16983 1455 16989
rect 1397 16949 1409 16983
rect 1443 16980 1455 16983
rect 1486 16980 1492 16992
rect 1443 16952 1492 16980
rect 1443 16949 1455 16952
rect 1397 16943 1455 16949
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 2547 16983 2605 16989
rect 2547 16949 2559 16983
rect 2593 16980 2605 16983
rect 2682 16980 2688 16992
rect 2593 16952 2688 16980
rect 2593 16949 2605 16952
rect 2547 16943 2605 16949
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 5074 16940 5080 16992
rect 5132 16980 5138 16992
rect 5276 16980 5304 17011
rect 6454 17008 6460 17020
rect 6512 17008 6518 17060
rect 6546 17008 6552 17060
rect 6604 17048 6610 17060
rect 7285 17051 7343 17057
rect 7285 17048 7297 17051
rect 6604 17020 7297 17048
rect 6604 17008 6610 17020
rect 7285 17017 7297 17020
rect 7331 17048 7343 17051
rect 7926 17048 7932 17060
rect 7331 17020 7932 17048
rect 7331 17017 7343 17020
rect 7285 17011 7343 17017
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 9677 17051 9735 17057
rect 9677 17048 9689 17051
rect 8864 17020 9689 17048
rect 8864 16992 8892 17020
rect 9677 17017 9689 17020
rect 9723 17017 9735 17051
rect 9677 17011 9735 17017
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 10321 17051 10379 17057
rect 9824 17020 9869 17048
rect 9824 17008 9830 17020
rect 10321 17017 10333 17051
rect 10367 17048 10379 17051
rect 10870 17048 10876 17060
rect 10367 17020 10876 17048
rect 10367 17017 10379 17020
rect 10321 17011 10379 17017
rect 10870 17008 10876 17020
rect 10928 17008 10934 17060
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17017 12679 17051
rect 14001 17051 14059 17057
rect 14001 17048 14013 17051
rect 12621 17011 12679 17017
rect 13280 17020 14013 17048
rect 5132 16952 5304 16980
rect 8757 16983 8815 16989
rect 5132 16940 5138 16952
rect 8757 16949 8769 16983
rect 8803 16980 8815 16983
rect 8846 16980 8852 16992
rect 8803 16952 8852 16980
rect 8803 16949 8815 16952
rect 8757 16943 8815 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9784 16980 9812 17008
rect 9539 16952 9812 16980
rect 12253 16983 12311 16989
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 12253 16949 12265 16983
rect 12299 16980 12311 16983
rect 12636 16980 12664 17011
rect 13280 16980 13308 17020
rect 14001 17017 14013 17020
rect 14047 17017 14059 17051
rect 15562 17048 15568 17060
rect 15523 17020 15568 17048
rect 14001 17011 14059 17017
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 18322 17048 18328 17060
rect 18283 17020 18328 17048
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 20070 17008 20076 17060
rect 20128 17048 20134 17060
rect 21358 17048 21364 17060
rect 20128 17020 20173 17048
rect 21271 17020 21364 17048
rect 20128 17008 20134 17020
rect 21358 17008 21364 17020
rect 21416 17048 21422 17060
rect 21637 17051 21695 17057
rect 21637 17048 21649 17051
rect 21416 17020 21649 17048
rect 21416 17008 21422 17020
rect 21637 17017 21649 17020
rect 21683 17017 21695 17051
rect 22186 17048 22192 17060
rect 22147 17020 22192 17048
rect 21637 17011 21695 17017
rect 22186 17008 22192 17020
rect 22244 17008 22250 17060
rect 13538 16980 13544 16992
rect 12299 16952 13308 16980
rect 13499 16952 13544 16980
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 19150 16980 19156 16992
rect 19111 16952 19156 16980
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 19797 16983 19855 16989
rect 19797 16949 19809 16983
rect 19843 16980 19855 16983
rect 20088 16980 20116 17008
rect 19843 16952 20116 16980
rect 19843 16949 19855 16952
rect 19797 16943 19855 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 2501 16779 2559 16785
rect 2501 16776 2513 16779
rect 1728 16748 2513 16776
rect 1728 16736 1734 16748
rect 2501 16745 2513 16748
rect 2547 16745 2559 16779
rect 2501 16739 2559 16745
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7193 16779 7251 16785
rect 7193 16776 7205 16779
rect 6972 16748 7205 16776
rect 6972 16736 6978 16748
rect 7193 16745 7205 16748
rect 7239 16745 7251 16779
rect 10042 16776 10048 16788
rect 10003 16748 10048 16776
rect 7193 16739 7251 16745
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 10597 16779 10655 16785
rect 10597 16776 10609 16779
rect 10192 16748 10609 16776
rect 10192 16736 10198 16748
rect 10597 16745 10609 16748
rect 10643 16745 10655 16779
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 10597 16739 10655 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 17034 16776 17040 16788
rect 16995 16748 17040 16776
rect 17034 16736 17040 16748
rect 17092 16736 17098 16788
rect 17494 16736 17500 16788
rect 17552 16776 17558 16788
rect 17589 16779 17647 16785
rect 17589 16776 17601 16779
rect 17552 16748 17601 16776
rect 17552 16736 17558 16748
rect 17589 16745 17601 16748
rect 17635 16745 17647 16779
rect 17589 16739 17647 16745
rect 19150 16736 19156 16788
rect 19208 16776 19214 16788
rect 19208 16748 21128 16776
rect 19208 16736 19214 16748
rect 21100 16720 21128 16748
rect 4798 16708 4804 16720
rect 4759 16680 4804 16708
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 6362 16708 6368 16720
rect 6323 16680 6368 16708
rect 6362 16668 6368 16680
rect 6420 16668 6426 16720
rect 7558 16668 7564 16720
rect 7616 16708 7622 16720
rect 7837 16711 7895 16717
rect 7837 16708 7849 16711
rect 7616 16680 7849 16708
rect 7616 16668 7622 16680
rect 7837 16677 7849 16680
rect 7883 16677 7895 16711
rect 7837 16671 7895 16677
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 7984 16680 8029 16708
rect 7984 16668 7990 16680
rect 11606 16668 11612 16720
rect 11664 16708 11670 16720
rect 11838 16711 11896 16717
rect 11838 16708 11850 16711
rect 11664 16680 11850 16708
rect 11664 16668 11670 16680
rect 11838 16677 11850 16680
rect 11884 16677 11896 16711
rect 13446 16708 13452 16720
rect 13407 16680 13452 16708
rect 11838 16671 11896 16677
rect 13446 16668 13452 16680
rect 13504 16708 13510 16720
rect 15562 16708 15568 16720
rect 13504 16680 15568 16708
rect 13504 16668 13510 16680
rect 15562 16668 15568 16680
rect 15620 16668 15626 16720
rect 19426 16708 19432 16720
rect 19387 16680 19432 16708
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 19981 16711 20039 16717
rect 19981 16677 19993 16711
rect 20027 16708 20039 16711
rect 20530 16708 20536 16720
rect 20027 16680 20536 16708
rect 20027 16677 20039 16680
rect 19981 16671 20039 16677
rect 20530 16668 20536 16680
rect 20588 16668 20594 16720
rect 21082 16708 21088 16720
rect 20995 16680 21088 16708
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 12434 16640 12440 16652
rect 12347 16612 12440 16640
rect 12434 16600 12440 16612
rect 12492 16640 12498 16652
rect 13170 16640 13176 16652
rect 12492 16612 13176 16640
rect 12492 16600 12498 16612
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 22002 16600 22008 16652
rect 22060 16640 22066 16652
rect 22462 16640 22468 16652
rect 22060 16612 22468 16640
rect 22060 16600 22066 16612
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 4706 16572 4712 16584
rect 4667 16544 4712 16572
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 4982 16572 4988 16584
rect 4943 16544 4988 16572
rect 4982 16532 4988 16544
rect 5040 16572 5046 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5040 16544 6009 16572
rect 5040 16532 5046 16544
rect 5997 16541 6009 16544
rect 6043 16572 6055 16575
rect 6273 16575 6331 16581
rect 6273 16572 6285 16575
rect 6043 16544 6285 16572
rect 6043 16541 6055 16544
rect 5997 16535 6055 16541
rect 6273 16541 6285 16544
rect 6319 16541 6331 16575
rect 6273 16535 6331 16541
rect 6454 16532 6460 16584
rect 6512 16572 6518 16584
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6512 16544 6561 16572
rect 6512 16532 6518 16544
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 8110 16572 8116 16584
rect 8071 16544 8116 16572
rect 6549 16535 6607 16541
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 9677 16575 9735 16581
rect 9677 16572 9689 16575
rect 9456 16544 9689 16572
rect 9456 16532 9462 16544
rect 9677 16541 9689 16544
rect 9723 16541 9735 16575
rect 9677 16535 9735 16541
rect 11517 16575 11575 16581
rect 11517 16541 11529 16575
rect 11563 16572 11575 16575
rect 12066 16572 12072 16584
rect 11563 16544 12072 16572
rect 11563 16541 11575 16544
rect 11517 16535 11575 16541
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 13354 16572 13360 16584
rect 13315 16544 13360 16572
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 13633 16575 13691 16581
rect 13633 16541 13645 16575
rect 13679 16572 13691 16575
rect 13998 16572 14004 16584
rect 13679 16544 14004 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 13648 16504 13676 16535
rect 13998 16532 14004 16544
rect 14056 16532 14062 16584
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15887 16544 16129 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 16117 16541 16129 16544
rect 16163 16572 16175 16575
rect 16482 16572 16488 16584
rect 16163 16544 16488 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 16666 16572 16672 16584
rect 16627 16544 16672 16572
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 19337 16575 19395 16581
rect 19337 16572 19349 16575
rect 18564 16544 19349 16572
rect 18564 16532 18570 16544
rect 19337 16541 19349 16544
rect 19383 16541 19395 16575
rect 19337 16535 19395 16541
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 20772 16544 21005 16572
rect 20772 16532 20778 16544
rect 20993 16541 21005 16544
rect 21039 16572 21051 16575
rect 22603 16575 22661 16581
rect 22603 16572 22615 16575
rect 21039 16544 22615 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 22603 16541 22615 16544
rect 22649 16541 22661 16575
rect 22603 16535 22661 16541
rect 12400 16476 13676 16504
rect 18233 16507 18291 16513
rect 12400 16464 12406 16476
rect 18233 16473 18245 16507
rect 18279 16504 18291 16507
rect 18322 16504 18328 16516
rect 18279 16476 18328 16504
rect 18279 16473 18291 16476
rect 18233 16467 18291 16473
rect 18322 16464 18328 16476
rect 18380 16504 18386 16516
rect 18966 16504 18972 16516
rect 18380 16476 18972 16504
rect 18380 16464 18386 16476
rect 18966 16464 18972 16476
rect 19024 16464 19030 16516
rect 20162 16464 20168 16516
rect 20220 16504 20226 16516
rect 21545 16507 21603 16513
rect 21545 16504 21557 16507
rect 20220 16476 21557 16504
rect 20220 16464 20226 16476
rect 21545 16473 21557 16476
rect 21591 16473 21603 16507
rect 21545 16467 21603 16473
rect 1762 16436 1768 16448
rect 1723 16408 1768 16436
rect 1762 16396 1768 16408
rect 1820 16396 1826 16448
rect 3605 16439 3663 16445
rect 3605 16405 3617 16439
rect 3651 16436 3663 16439
rect 3970 16436 3976 16448
rect 3651 16408 3976 16436
rect 3651 16405 3663 16408
rect 3605 16399 3663 16405
rect 3970 16396 3976 16408
rect 4028 16396 4034 16448
rect 4338 16396 4344 16448
rect 4396 16436 4402 16448
rect 4433 16439 4491 16445
rect 4433 16436 4445 16439
rect 4396 16408 4445 16436
rect 4396 16396 4402 16408
rect 4433 16405 4445 16408
rect 4479 16405 4491 16439
rect 4433 16399 4491 16405
rect 7653 16439 7711 16445
rect 7653 16405 7665 16439
rect 7699 16436 7711 16439
rect 7742 16436 7748 16448
rect 7699 16408 7748 16436
rect 7699 16405 7711 16408
rect 7653 16399 7711 16405
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 8478 16396 8484 16448
rect 8536 16436 8542 16448
rect 8757 16439 8815 16445
rect 8757 16436 8769 16439
rect 8536 16408 8769 16436
rect 8536 16396 8542 16408
rect 8757 16405 8769 16408
rect 8803 16405 8815 16439
rect 10870 16436 10876 16448
rect 10831 16408 10876 16436
rect 8757 16399 8815 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 18874 16436 18880 16448
rect 18835 16408 18880 16436
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 5353 16235 5411 16241
rect 5353 16201 5365 16235
rect 5399 16232 5411 16235
rect 5442 16232 5448 16244
rect 5399 16204 5448 16232
rect 5399 16201 5411 16204
rect 5353 16195 5411 16201
rect 5442 16192 5448 16204
rect 5500 16232 5506 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5500 16204 6193 16232
rect 5500 16192 5506 16204
rect 6181 16201 6193 16204
rect 6227 16201 6239 16235
rect 7926 16232 7932 16244
rect 7887 16204 7932 16232
rect 6181 16195 6239 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 9490 16232 9496 16244
rect 9451 16204 9496 16232
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10100 16204 11529 16232
rect 10100 16192 10106 16204
rect 11517 16201 11529 16204
rect 11563 16232 11575 16235
rect 11606 16232 11612 16244
rect 11563 16204 11612 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 13265 16235 13323 16241
rect 13265 16201 13277 16235
rect 13311 16232 13323 16235
rect 13446 16232 13452 16244
rect 13311 16204 13452 16232
rect 13311 16201 13323 16204
rect 13265 16195 13323 16201
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14921 16235 14979 16241
rect 14921 16232 14933 16235
rect 14323 16204 14933 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 14921 16201 14933 16204
rect 14967 16232 14979 16235
rect 15286 16232 15292 16244
rect 14967 16204 15292 16232
rect 14967 16201 14979 16204
rect 14921 16195 14979 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 18506 16232 18512 16244
rect 18371 16204 18512 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 19705 16235 19763 16241
rect 19705 16232 19717 16235
rect 19484 16204 19717 16232
rect 19484 16192 19490 16204
rect 19705 16201 19717 16204
rect 19751 16232 19763 16235
rect 19981 16235 20039 16241
rect 19981 16232 19993 16235
rect 19751 16204 19993 16232
rect 19751 16201 19763 16204
rect 19705 16195 19763 16201
rect 19981 16201 19993 16204
rect 20027 16201 20039 16235
rect 19981 16195 20039 16201
rect 21082 16192 21088 16244
rect 21140 16232 21146 16244
rect 21729 16235 21787 16241
rect 21729 16232 21741 16235
rect 21140 16204 21741 16232
rect 21140 16192 21146 16204
rect 21729 16201 21741 16204
rect 21775 16232 21787 16235
rect 22738 16232 22744 16244
rect 21775 16204 22744 16232
rect 21775 16201 21787 16204
rect 21729 16195 21787 16201
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 3605 16167 3663 16173
rect 3605 16133 3617 16167
rect 3651 16164 3663 16167
rect 7098 16164 7104 16176
rect 3651 16136 7104 16164
rect 3651 16133 3663 16136
rect 3605 16127 3663 16133
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 1670 16096 1676 16108
rect 1627 16068 1676 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 1912 16068 2881 16096
rect 1912 16056 1918 16068
rect 2869 16065 2881 16068
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 3120 16031 3178 16037
rect 3120 15997 3132 16031
rect 3166 16028 3178 16031
rect 3620 16028 3648 16127
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 10962 16164 10968 16176
rect 10923 16136 10968 16164
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 12897 16167 12955 16173
rect 12897 16133 12909 16167
rect 12943 16164 12955 16167
rect 13354 16164 13360 16176
rect 12943 16136 13360 16164
rect 12943 16133 12955 16136
rect 12897 16127 12955 16133
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 13998 16164 14004 16176
rect 13959 16136 14004 16164
rect 13998 16124 14004 16136
rect 14056 16124 14062 16176
rect 15151 16167 15209 16173
rect 15151 16133 15163 16167
rect 15197 16164 15209 16167
rect 18414 16164 18420 16176
rect 15197 16136 18420 16164
rect 15197 16133 15209 16136
rect 15151 16127 15209 16133
rect 18414 16124 18420 16136
rect 18472 16124 18478 16176
rect 18874 16164 18880 16176
rect 18787 16136 18880 16164
rect 3973 16099 4031 16105
rect 3973 16065 3985 16099
rect 4019 16096 4031 16099
rect 4798 16096 4804 16108
rect 4019 16068 4804 16096
rect 4019 16065 4031 16068
rect 3973 16059 4031 16065
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 7561 16099 7619 16105
rect 7561 16065 7573 16099
rect 7607 16096 7619 16099
rect 8110 16096 8116 16108
rect 7607 16068 8116 16096
rect 7607 16065 7619 16068
rect 7561 16059 7619 16065
rect 8110 16056 8116 16068
rect 8168 16096 8174 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 8168 16068 10425 16096
rect 8168 16056 8174 16068
rect 10413 16065 10425 16068
rect 10459 16096 10471 16099
rect 10870 16096 10876 16108
rect 10459 16068 10876 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 14366 16096 14372 16108
rect 13495 16068 14372 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 18800 16105 18828 16136
rect 18874 16124 18880 16136
rect 18932 16164 18938 16176
rect 21818 16164 21824 16176
rect 18932 16136 21824 16164
rect 18932 16124 18938 16136
rect 21818 16124 21824 16136
rect 21876 16124 21882 16176
rect 16761 16099 16819 16105
rect 16761 16096 16773 16099
rect 16724 16068 16773 16096
rect 16724 16056 16730 16068
rect 16761 16065 16773 16068
rect 16807 16096 16819 16099
rect 17405 16099 17463 16105
rect 17405 16096 17417 16099
rect 16807 16068 17417 16096
rect 16807 16065 16819 16068
rect 16761 16059 16819 16065
rect 17405 16065 17417 16068
rect 17451 16065 17463 16099
rect 17405 16059 17463 16065
rect 18785 16099 18843 16105
rect 18785 16065 18797 16099
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16096 20867 16099
rect 22189 16099 22247 16105
rect 22189 16096 22201 16099
rect 20855 16068 22201 16096
rect 20855 16065 20867 16068
rect 20809 16059 20867 16065
rect 22189 16065 22201 16068
rect 22235 16096 22247 16099
rect 22554 16096 22560 16108
rect 22235 16068 22560 16096
rect 22235 16065 22247 16068
rect 22189 16059 22247 16065
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 3166 16000 3648 16028
rect 3166 15997 3178 16000
rect 3120 15991 3178 15997
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 4396 16000 4445 16028
rect 4396 15988 4402 16000
rect 4433 15997 4445 16000
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 8478 15988 8484 16040
rect 8536 16028 8542 16040
rect 8573 16031 8631 16037
rect 8573 16028 8585 16031
rect 8536 16000 8585 16028
rect 8536 15988 8542 16000
rect 8573 15997 8585 16000
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 14918 15988 14924 16040
rect 14976 16028 14982 16040
rect 15048 16031 15106 16037
rect 15048 16028 15060 16031
rect 14976 16000 15060 16028
rect 14976 15988 14982 16000
rect 15048 15997 15060 16000
rect 15094 16028 15106 16031
rect 15473 16031 15531 16037
rect 15473 16028 15485 16031
rect 15094 16000 15485 16028
rect 15094 15997 15106 16000
rect 15048 15991 15106 15997
rect 15473 15997 15485 16000
rect 15519 15997 15531 16031
rect 16022 16028 16028 16040
rect 15983 16000 16028 16028
rect 15473 15991 15531 15997
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 16482 16028 16488 16040
rect 16443 16000 16488 16028
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 18966 15988 18972 16040
rect 19024 16028 19030 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 19024 16000 20545 16028
rect 19024 15988 19030 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 1673 15963 1731 15969
rect 1673 15929 1685 15963
rect 1719 15960 1731 15963
rect 1762 15960 1768 15972
rect 1719 15932 1768 15960
rect 1719 15929 1731 15932
rect 1673 15923 1731 15929
rect 1762 15920 1768 15932
rect 1820 15920 1826 15972
rect 2225 15963 2283 15969
rect 2225 15929 2237 15963
rect 2271 15960 2283 15963
rect 2406 15960 2412 15972
rect 2271 15932 2412 15960
rect 2271 15929 2283 15932
rect 2225 15923 2283 15929
rect 2406 15920 2412 15932
rect 2464 15920 2470 15972
rect 4522 15920 4528 15972
rect 4580 15960 4586 15972
rect 5813 15963 5871 15969
rect 5813 15960 5825 15963
rect 4580 15932 5825 15960
rect 4580 15920 4586 15932
rect 5813 15929 5825 15932
rect 5859 15960 5871 15963
rect 6917 15963 6975 15969
rect 6917 15960 6929 15963
rect 5859 15932 6929 15960
rect 5859 15929 5871 15932
rect 5813 15923 5871 15929
rect 6917 15929 6929 15932
rect 6963 15929 6975 15963
rect 6917 15923 6975 15929
rect 7009 15963 7067 15969
rect 7009 15929 7021 15963
rect 7055 15960 7067 15963
rect 7742 15960 7748 15972
rect 7055 15932 7748 15960
rect 7055 15929 7067 15932
rect 7009 15923 7067 15929
rect 1780 15892 1808 15920
rect 2501 15895 2559 15901
rect 2501 15892 2513 15895
rect 1780 15864 2513 15892
rect 2501 15861 2513 15864
rect 2547 15861 2559 15895
rect 2501 15855 2559 15861
rect 3191 15895 3249 15901
rect 3191 15861 3203 15895
rect 3237 15892 3249 15895
rect 3326 15892 3332 15904
rect 3237 15864 3332 15892
rect 3237 15861 3249 15864
rect 3191 15855 3249 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 4212 15864 4353 15892
rect 4212 15852 4218 15864
rect 4341 15861 4353 15864
rect 4387 15892 4399 15895
rect 4801 15895 4859 15901
rect 4801 15892 4813 15895
rect 4387 15864 4813 15892
rect 4387 15861 4399 15864
rect 4341 15855 4399 15861
rect 4801 15861 4813 15864
rect 4847 15861 4859 15895
rect 4801 15855 4859 15861
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7024 15892 7052 15923
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 8894 15963 8952 15969
rect 8894 15960 8906 15963
rect 8404 15932 8906 15960
rect 8404 15904 8432 15932
rect 8894 15929 8906 15932
rect 8940 15960 8952 15963
rect 9769 15963 9827 15969
rect 9769 15960 9781 15963
rect 8940 15932 9781 15960
rect 8940 15929 8952 15932
rect 8894 15923 8952 15929
rect 9769 15929 9781 15932
rect 9815 15960 9827 15963
rect 10042 15960 10048 15972
rect 9815 15932 10048 15960
rect 9815 15929 9827 15932
rect 9769 15923 9827 15929
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 10505 15963 10563 15969
rect 10505 15929 10517 15963
rect 10551 15929 10563 15963
rect 10505 15923 10563 15929
rect 13541 15963 13599 15969
rect 13541 15929 13553 15963
rect 13587 15960 13599 15963
rect 15654 15960 15660 15972
rect 13587 15932 15660 15960
rect 13587 15929 13599 15932
rect 13541 15923 13599 15929
rect 8386 15892 8392 15904
rect 6687 15864 7052 15892
rect 8347 15864 8392 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 10134 15892 10140 15904
rect 10095 15864 10140 15892
rect 10134 15852 10140 15864
rect 10192 15892 10198 15904
rect 10520 15892 10548 15923
rect 10192 15864 10548 15892
rect 11977 15895 12035 15901
rect 10192 15852 10198 15864
rect 11977 15861 11989 15895
rect 12023 15892 12035 15895
rect 12066 15892 12072 15904
rect 12023 15864 12072 15892
rect 12023 15861 12035 15864
rect 11977 15855 12035 15861
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13556 15892 13584 15923
rect 15654 15920 15660 15932
rect 15712 15920 15718 15972
rect 19106 15963 19164 15969
rect 19106 15960 19118 15963
rect 18616 15932 19118 15960
rect 13412 15864 13584 15892
rect 13412 15852 13418 15864
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13688 15864 14289 15892
rect 13688 15852 13694 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 14366 15852 14372 15904
rect 14424 15892 14430 15904
rect 14424 15864 14469 15892
rect 14424 15852 14430 15864
rect 15470 15852 15476 15904
rect 15528 15892 15534 15904
rect 15841 15895 15899 15901
rect 15841 15892 15853 15895
rect 15528 15864 15853 15892
rect 15528 15852 15534 15864
rect 15841 15861 15853 15864
rect 15887 15861 15899 15895
rect 17034 15892 17040 15904
rect 16995 15864 17040 15892
rect 15841 15855 15899 15861
rect 17034 15852 17040 15864
rect 17092 15892 17098 15904
rect 18616 15901 18644 15932
rect 19106 15929 19118 15932
rect 19152 15960 19164 15963
rect 19426 15960 19432 15972
rect 19152 15932 19432 15960
rect 19152 15929 19164 15932
rect 19106 15923 19164 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 20548 15960 20576 15991
rect 20901 15963 20959 15969
rect 20901 15960 20913 15963
rect 20548 15932 20913 15960
rect 20901 15929 20913 15932
rect 20947 15929 20959 15963
rect 20901 15923 20959 15929
rect 21082 15920 21088 15972
rect 21140 15960 21146 15972
rect 21453 15963 21511 15969
rect 21453 15960 21465 15963
rect 21140 15932 21465 15960
rect 21140 15920 21146 15932
rect 21453 15929 21465 15932
rect 21499 15960 21511 15963
rect 22186 15960 22192 15972
rect 21499 15932 22192 15960
rect 21499 15929 21511 15932
rect 21453 15923 21511 15929
rect 22186 15920 22192 15932
rect 22244 15960 22250 15972
rect 22922 15960 22928 15972
rect 22244 15932 22928 15960
rect 22244 15920 22250 15932
rect 22922 15920 22928 15932
rect 22980 15920 22986 15972
rect 18601 15895 18659 15901
rect 18601 15892 18613 15895
rect 17092 15864 18613 15892
rect 17092 15852 17098 15864
rect 18601 15861 18613 15864
rect 18647 15861 18659 15895
rect 22462 15892 22468 15904
rect 22423 15864 22468 15892
rect 18601 15855 18659 15861
rect 22462 15852 22468 15864
rect 22520 15852 22526 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2682 15688 2688 15700
rect 1780 15660 2688 15688
rect 1780 15629 1808 15660
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4706 15688 4712 15700
rect 3927 15660 4712 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 4985 15691 5043 15697
rect 4985 15688 4997 15691
rect 4856 15660 4997 15688
rect 4856 15648 4862 15660
rect 4985 15657 4997 15660
rect 5031 15657 5043 15691
rect 7006 15688 7012 15700
rect 6967 15660 7012 15688
rect 4985 15651 5043 15657
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7616 15660 7849 15688
rect 7616 15648 7622 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 8711 15691 8769 15697
rect 8711 15657 8723 15691
rect 8757 15688 8769 15691
rect 8846 15688 8852 15700
rect 8757 15660 8852 15688
rect 8757 15657 8769 15660
rect 8711 15651 8769 15657
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 9824 15660 10609 15688
rect 9824 15648 9830 15660
rect 10597 15657 10609 15660
rect 10643 15657 10655 15691
rect 10597 15651 10655 15657
rect 12345 15691 12403 15697
rect 12345 15657 12357 15691
rect 12391 15688 12403 15691
rect 13538 15688 13544 15700
rect 12391 15660 13544 15688
rect 12391 15657 12403 15660
rect 12345 15651 12403 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 14734 15688 14740 15700
rect 13740 15660 14740 15688
rect 1765 15623 1823 15629
rect 1765 15589 1777 15623
rect 1811 15589 1823 15623
rect 1765 15583 1823 15589
rect 1854 15580 1860 15632
rect 1912 15620 1918 15632
rect 2406 15620 2412 15632
rect 1912 15592 1957 15620
rect 2367 15592 2412 15620
rect 1912 15580 1918 15592
rect 2406 15580 2412 15592
rect 2464 15580 2470 15632
rect 3786 15580 3792 15632
rect 3844 15620 3850 15632
rect 4154 15620 4160 15632
rect 3844 15592 4160 15620
rect 3844 15580 3850 15592
rect 4154 15580 4160 15592
rect 4212 15620 4218 15632
rect 10042 15629 10048 15632
rect 4386 15623 4444 15629
rect 4386 15620 4398 15623
rect 4212 15592 4398 15620
rect 4212 15580 4218 15592
rect 4386 15589 4398 15592
rect 4432 15589 4444 15623
rect 10039 15620 10048 15629
rect 10003 15592 10048 15620
rect 4386 15583 4444 15589
rect 10039 15583 10048 15592
rect 10042 15580 10048 15583
rect 10100 15580 10106 15632
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 13740 15629 13768 15660
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15838 15648 15844 15700
rect 15896 15688 15902 15700
rect 16022 15688 16028 15700
rect 15896 15660 16028 15688
rect 15896 15648 15902 15660
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 17313 15691 17371 15697
rect 17313 15657 17325 15691
rect 17359 15688 17371 15691
rect 19150 15688 19156 15700
rect 17359 15660 19156 15688
rect 17359 15657 17371 15660
rect 17313 15651 17371 15657
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 19426 15688 19432 15700
rect 19387 15660 19432 15688
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19981 15691 20039 15697
rect 19981 15657 19993 15691
rect 20027 15688 20039 15691
rect 20070 15688 20076 15700
rect 20027 15660 20076 15688
rect 20027 15657 20039 15660
rect 19981 15651 20039 15657
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 20714 15688 20720 15700
rect 20675 15660 20720 15688
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 11746 15623 11804 15629
rect 11746 15620 11758 15623
rect 11664 15592 11758 15620
rect 11664 15580 11670 15592
rect 11746 15589 11758 15592
rect 11792 15589 11804 15623
rect 11746 15583 11804 15589
rect 13725 15623 13783 15629
rect 13725 15589 13737 15623
rect 13771 15589 13783 15623
rect 13725 15583 13783 15589
rect 13817 15623 13875 15629
rect 13817 15589 13829 15623
rect 13863 15620 13875 15623
rect 13906 15620 13912 15632
rect 13863 15592 13912 15620
rect 13863 15589 13875 15592
rect 13817 15583 13875 15589
rect 13906 15580 13912 15592
rect 13964 15580 13970 15632
rect 16206 15580 16212 15632
rect 16264 15620 16270 15632
rect 16714 15623 16772 15629
rect 16714 15620 16726 15623
rect 16264 15592 16726 15620
rect 16264 15580 16270 15592
rect 16714 15589 16726 15592
rect 16760 15620 16772 15623
rect 17034 15620 17040 15632
rect 16760 15592 17040 15620
rect 16760 15589 16772 15592
rect 16714 15583 16772 15589
rect 17034 15580 17040 15592
rect 17092 15580 17098 15632
rect 21174 15620 21180 15632
rect 21135 15592 21180 15620
rect 21174 15580 21180 15592
rect 21232 15580 21238 15632
rect 21726 15620 21732 15632
rect 21687 15592 21732 15620
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 22738 15620 22744 15632
rect 22699 15592 22744 15620
rect 22738 15580 22744 15592
rect 22796 15580 22802 15632
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15552 7619 15555
rect 7926 15552 7932 15564
rect 7607 15524 7932 15552
rect 7607 15521 7619 15524
rect 7561 15515 7619 15521
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 8570 15552 8576 15564
rect 8531 15524 8576 15552
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 15356 15555 15414 15561
rect 15356 15521 15368 15555
rect 15402 15552 15414 15555
rect 15746 15552 15752 15564
rect 15402 15524 15752 15552
rect 15402 15521 15414 15524
rect 15356 15515 15414 15521
rect 15746 15512 15752 15524
rect 15804 15512 15810 15564
rect 16298 15512 16304 15564
rect 16356 15552 16362 15564
rect 20162 15552 20168 15564
rect 16356 15524 20168 15552
rect 16356 15512 16362 15524
rect 20162 15512 20168 15524
rect 20220 15512 20226 15564
rect 24210 15512 24216 15564
rect 24268 15552 24274 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 24268 15524 24593 15552
rect 24268 15512 24274 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 24762 15512 24768 15564
rect 24820 15552 24826 15564
rect 27614 15552 27620 15564
rect 24820 15524 27620 15552
rect 24820 15512 24826 15524
rect 27614 15512 27620 15524
rect 27672 15512 27678 15564
rect 4062 15484 4068 15496
rect 4023 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 6641 15487 6699 15493
rect 6641 15453 6653 15487
rect 6687 15453 6699 15487
rect 9674 15484 9680 15496
rect 9635 15456 9680 15484
rect 6641 15447 6699 15453
rect 2958 15308 2964 15360
rect 3016 15348 3022 15360
rect 3053 15351 3111 15357
rect 3053 15348 3065 15351
rect 3016 15320 3065 15348
rect 3016 15308 3022 15320
rect 3053 15317 3065 15320
rect 3099 15348 3111 15351
rect 4890 15348 4896 15360
rect 3099 15320 4896 15348
rect 3099 15317 3111 15320
rect 3053 15311 3111 15317
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5534 15348 5540 15360
rect 5495 15320 5540 15348
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 6178 15348 6184 15360
rect 6139 15320 6184 15348
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 6656 15348 6684 15447
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 11422 15484 11428 15496
rect 11335 15456 11428 15484
rect 11422 15444 11428 15456
rect 11480 15484 11486 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 11480 15456 12633 15484
rect 11480 15444 11486 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 14366 15484 14372 15496
rect 14327 15456 14372 15484
rect 12621 15447 12679 15453
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 17402 15484 17408 15496
rect 16439 15456 17408 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 17402 15444 17408 15456
rect 17460 15444 17466 15496
rect 19061 15487 19119 15493
rect 19061 15453 19073 15487
rect 19107 15453 19119 15487
rect 19061 15447 19119 15453
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 21082 15484 21088 15496
rect 20395 15456 21088 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 12250 15376 12256 15428
rect 12308 15416 12314 15428
rect 12989 15419 13047 15425
rect 12989 15416 13001 15419
rect 12308 15388 13001 15416
rect 12308 15376 12314 15388
rect 12989 15385 13001 15388
rect 13035 15385 13047 15419
rect 12989 15379 13047 15385
rect 6914 15348 6920 15360
rect 6595 15320 6920 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 9030 15348 9036 15360
rect 8991 15320 9036 15348
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 9398 15348 9404 15360
rect 9359 15320 9404 15348
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 10962 15348 10968 15360
rect 10923 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11238 15348 11244 15360
rect 11199 15320 11244 15348
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 13354 15348 13360 15360
rect 13315 15320 13360 15348
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15427 15351 15485 15357
rect 15427 15348 15439 15351
rect 14792 15320 15439 15348
rect 14792 15308 14798 15320
rect 15427 15317 15439 15320
rect 15473 15317 15485 15351
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 15427 15311 15485 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 18969 15351 19027 15357
rect 18969 15317 18981 15351
rect 19015 15348 19027 15351
rect 19076 15348 19104 15447
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15484 22707 15487
rect 22738 15484 22744 15496
rect 22695 15456 22744 15484
rect 22695 15453 22707 15456
rect 22649 15447 22707 15453
rect 22738 15444 22744 15456
rect 22796 15444 22802 15496
rect 22922 15484 22928 15496
rect 22883 15456 22928 15484
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 19518 15348 19524 15360
rect 19015 15320 19524 15348
rect 19015 15317 19027 15320
rect 18969 15311 19027 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1854 15104 1860 15156
rect 1912 15144 1918 15156
rect 2685 15147 2743 15153
rect 2685 15144 2697 15147
rect 1912 15116 2697 15144
rect 1912 15104 1918 15116
rect 2685 15113 2697 15116
rect 2731 15144 2743 15147
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2731 15116 2973 15144
rect 2731 15113 2743 15116
rect 2685 15107 2743 15113
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 2961 15107 3019 15113
rect 4890 15104 4896 15156
rect 4948 15144 4954 15156
rect 5675 15147 5733 15153
rect 5675 15144 5687 15147
rect 4948 15116 5687 15144
rect 4948 15104 4954 15116
rect 5675 15113 5687 15116
rect 5721 15113 5733 15147
rect 7742 15144 7748 15156
rect 7703 15116 7748 15144
rect 5675 15107 5733 15113
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 8570 15144 8576 15156
rect 8531 15116 8576 15144
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 9769 15147 9827 15153
rect 9769 15113 9781 15147
rect 9815 15144 9827 15147
rect 10134 15144 10140 15156
rect 9815 15116 10140 15144
rect 9815 15113 9827 15116
rect 9769 15107 9827 15113
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 11606 15144 11612 15156
rect 11567 15116 11612 15144
rect 11606 15104 11612 15116
rect 11664 15144 11670 15156
rect 12158 15144 12164 15156
rect 11664 15116 12164 15144
rect 11664 15104 11670 15116
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 13354 15144 13360 15156
rect 13315 15116 13360 15144
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 15381 15147 15439 15153
rect 15381 15113 15393 15147
rect 15427 15144 15439 15147
rect 15746 15144 15752 15156
rect 15427 15116 15752 15144
rect 15427 15113 15439 15116
rect 15381 15107 15439 15113
rect 15746 15104 15752 15116
rect 15804 15144 15810 15156
rect 16850 15144 16856 15156
rect 15804 15116 16856 15144
rect 15804 15104 15810 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17402 15144 17408 15156
rect 17363 15116 17408 15144
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 18966 15144 18972 15156
rect 18927 15116 18972 15144
rect 18966 15104 18972 15116
rect 19024 15104 19030 15156
rect 20901 15147 20959 15153
rect 20901 15113 20913 15147
rect 20947 15144 20959 15147
rect 21174 15144 21180 15156
rect 20947 15116 21180 15144
rect 20947 15113 20959 15116
rect 20901 15107 20959 15113
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 22830 15144 22836 15156
rect 22791 15116 22836 15144
rect 22830 15104 22836 15116
rect 22888 15104 22894 15156
rect 4062 15036 4068 15088
rect 4120 15076 4126 15088
rect 5353 15079 5411 15085
rect 5353 15076 5365 15079
rect 4120 15048 5365 15076
rect 4120 15036 4126 15048
rect 5353 15045 5365 15048
rect 5399 15045 5411 15079
rect 15838 15076 15844 15088
rect 5353 15039 5411 15045
rect 13786 15048 15844 15076
rect 3970 15008 3976 15020
rect 3931 14980 3976 15008
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4798 15008 4804 15020
rect 4632 14980 4804 15008
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 1811 14912 3341 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 3329 14909 3341 14912
rect 3375 14940 3387 14943
rect 3418 14940 3424 14952
rect 3375 14912 3424 14940
rect 3375 14909 3387 14912
rect 3329 14903 3387 14909
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 4632 14949 4660 14980
rect 4798 14968 4804 14980
rect 4856 15008 4862 15020
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4856 14980 4997 15008
rect 4856 14968 4862 14980
rect 4985 14977 4997 14980
rect 5031 14977 5043 15011
rect 4985 14971 5043 14977
rect 6178 14968 6184 15020
rect 6236 15008 6242 15020
rect 6730 15008 6736 15020
rect 6236 14980 6736 15008
rect 6236 14968 6242 14980
rect 6730 14968 6736 14980
rect 6788 15008 6794 15020
rect 6825 15011 6883 15017
rect 6825 15008 6837 15011
rect 6788 14980 6837 15008
rect 6788 14968 6794 14980
rect 6825 14977 6837 14980
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 8754 14968 8760 15020
rect 8812 15008 8818 15020
rect 8849 15011 8907 15017
rect 8849 15008 8861 15011
rect 8812 14980 8861 15008
rect 8812 14968 8818 14980
rect 8849 14977 8861 14980
rect 8895 15008 8907 15011
rect 9030 15008 9036 15020
rect 8895 14980 9036 15008
rect 8895 14977 8907 14980
rect 8849 14971 8907 14977
rect 9030 14968 9036 14980
rect 9088 14968 9094 15020
rect 13786 15008 13814 15048
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 19242 15076 19248 15088
rect 15948 15048 19248 15076
rect 14274 15008 14280 15020
rect 10888 14980 13814 15008
rect 14235 14980 14280 15008
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 5534 14940 5540 14952
rect 5495 14912 5540 14940
rect 4617 14903 4675 14909
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 10888 14949 10916 14980
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14424 14980 14565 15008
rect 14424 14968 14430 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 14642 14968 14648 15020
rect 14700 15008 14706 15020
rect 15948 15008 15976 15048
rect 19242 15036 19248 15048
rect 19300 15076 19306 15088
rect 24765 15079 24823 15085
rect 19300 15048 23474 15076
rect 19300 15036 19306 15048
rect 14700 14980 15976 15008
rect 17129 15011 17187 15017
rect 14700 14968 14706 14980
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 18046 15008 18052 15020
rect 17175 14980 18052 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 20990 14968 20996 15020
rect 21048 15008 21054 15020
rect 22738 15008 22744 15020
rect 21048 14980 22744 15008
rect 21048 14968 21054 14980
rect 22738 14968 22744 14980
rect 22796 15008 22802 15020
rect 23109 15011 23167 15017
rect 23109 15008 23121 15011
rect 22796 14980 23121 15008
rect 22796 14968 22802 14980
rect 23109 14977 23121 14980
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 9185 14912 10057 14940
rect 2086 14875 2144 14881
rect 2086 14872 2098 14875
rect 1688 14844 2098 14872
rect 1688 14816 1716 14844
rect 2086 14841 2098 14844
rect 2132 14872 2144 14875
rect 3786 14872 3792 14884
rect 2132 14844 3792 14872
rect 2132 14841 2144 14844
rect 2086 14835 2144 14841
rect 3786 14832 3792 14844
rect 3844 14872 3850 14884
rect 6181 14875 6239 14881
rect 6181 14872 6193 14875
rect 3844 14844 6193 14872
rect 3844 14832 3850 14844
rect 6181 14841 6193 14844
rect 6227 14872 6239 14875
rect 6549 14875 6607 14881
rect 6549 14872 6561 14875
rect 6227 14844 6561 14872
rect 6227 14841 6239 14844
rect 6181 14835 6239 14841
rect 6549 14841 6561 14844
rect 6595 14872 6607 14875
rect 7006 14872 7012 14884
rect 6595 14844 7012 14872
rect 6595 14841 6607 14844
rect 6549 14835 6607 14841
rect 7006 14832 7012 14844
rect 7064 14872 7070 14884
rect 7146 14875 7204 14881
rect 7146 14872 7158 14875
rect 7064 14844 7158 14872
rect 7064 14832 7070 14844
rect 7146 14841 7158 14844
rect 7192 14872 7204 14875
rect 7282 14872 7288 14884
rect 7192 14844 7288 14872
rect 7192 14841 7204 14844
rect 7146 14835 7204 14841
rect 7282 14832 7288 14844
rect 7340 14872 7346 14884
rect 8205 14875 8263 14881
rect 8205 14872 8217 14875
rect 7340 14844 8217 14872
rect 7340 14832 7346 14844
rect 8205 14841 8217 14844
rect 8251 14872 8263 14875
rect 8386 14872 8392 14884
rect 8251 14844 8392 14872
rect 8251 14841 8263 14844
rect 8205 14835 8263 14841
rect 8386 14832 8392 14844
rect 8444 14872 8450 14884
rect 9185 14881 9213 14912
rect 10045 14909 10057 14912
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 10505 14943 10563 14949
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10873 14943 10931 14949
rect 10873 14940 10885 14943
rect 10551 14912 10885 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10873 14909 10885 14912
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 11238 14940 11244 14952
rect 11195 14912 11244 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 9170 14875 9228 14881
rect 9170 14872 9182 14875
rect 8444 14844 9182 14872
rect 8444 14832 8450 14844
rect 9170 14841 9182 14844
rect 9216 14841 9228 14875
rect 9170 14835 9228 14841
rect 9306 14832 9312 14884
rect 9364 14872 9370 14884
rect 11164 14872 11192 14903
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 12250 14900 12256 14952
rect 12308 14940 12314 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12308 14912 12449 14940
rect 12308 14900 12314 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 16393 14943 16451 14949
rect 16393 14940 16405 14943
rect 12437 14903 12495 14909
rect 15856 14912 16405 14940
rect 9364 14844 11192 14872
rect 9364 14832 9370 14844
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 12802 14881 12808 14884
rect 12758 14875 12808 14881
rect 12758 14872 12770 14875
rect 12216 14844 12770 14872
rect 12216 14832 12222 14844
rect 12758 14841 12770 14844
rect 12804 14841 12808 14875
rect 12758 14835 12808 14841
rect 12802 14832 12808 14835
rect 12860 14832 12866 14884
rect 12986 14832 12992 14884
rect 13044 14872 13050 14884
rect 13630 14872 13636 14884
rect 13044 14844 13636 14872
rect 13044 14832 13050 14844
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 14369 14875 14427 14881
rect 14369 14841 14381 14875
rect 14415 14841 14427 14875
rect 14369 14835 14427 14841
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 10686 14804 10692 14816
rect 10647 14776 10692 14804
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 13906 14804 13912 14816
rect 13771 14776 13912 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14090 14804 14096 14816
rect 14051 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14804 14154 14816
rect 14384 14804 14412 14835
rect 14148 14776 14412 14804
rect 14148 14764 14154 14776
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 15856 14813 15884 14912
rect 16393 14909 16405 14912
rect 16439 14909 16451 14943
rect 16393 14903 16451 14909
rect 16482 14900 16488 14952
rect 16540 14940 16546 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16540 14912 16865 14940
rect 16540 14900 16546 14912
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 19978 14940 19984 14952
rect 19939 14912 19984 14940
rect 16853 14903 16911 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 21729 14943 21787 14949
rect 21729 14940 21741 14943
rect 21652 14912 21741 14940
rect 20346 14881 20352 14884
rect 18370 14875 18428 14881
rect 18370 14841 18382 14875
rect 18416 14872 18428 14875
rect 19245 14875 19303 14881
rect 19245 14872 19257 14875
rect 18416 14844 19257 14872
rect 18416 14841 18428 14844
rect 18370 14835 18428 14841
rect 19245 14841 19257 14844
rect 19291 14872 19303 14875
rect 19797 14875 19855 14881
rect 19797 14872 19809 14875
rect 19291 14844 19809 14872
rect 19291 14841 19303 14844
rect 19245 14835 19303 14841
rect 19797 14841 19809 14844
rect 19843 14872 19855 14875
rect 20302 14875 20352 14881
rect 20302 14872 20314 14875
rect 19843 14844 20314 14872
rect 19843 14841 19855 14844
rect 19797 14835 19855 14841
rect 20302 14841 20314 14844
rect 20348 14841 20352 14875
rect 20302 14835 20352 14841
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15712 14776 15853 14804
rect 15712 14764 15718 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 15841 14767 15899 14773
rect 16206 14764 16212 14776
rect 16264 14804 16270 14816
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 16264 14776 17785 14804
rect 16264 14764 16270 14776
rect 17773 14773 17785 14776
rect 17819 14804 17831 14807
rect 18385 14804 18413 14835
rect 20346 14832 20352 14835
rect 20404 14832 20410 14884
rect 21652 14816 21680 14912
rect 21729 14909 21741 14912
rect 21775 14909 21787 14943
rect 22186 14940 22192 14952
rect 22147 14912 22192 14940
rect 21729 14903 21787 14909
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 23446 14940 23474 15048
rect 24765 15045 24777 15079
rect 24811 15076 24823 15079
rect 27614 15076 27620 15088
rect 24811 15048 27620 15076
rect 24811 15045 24823 15048
rect 24765 15039 24823 15045
rect 27614 15036 27620 15048
rect 27672 15036 27678 15088
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 23446 14912 24593 14940
rect 24581 14909 24593 14912
rect 24627 14940 24639 14943
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24627 14912 25145 14940
rect 24627 14909 24639 14912
rect 24581 14903 24639 14909
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 17819 14776 18413 14804
rect 17819 14773 17831 14776
rect 17773 14767 17831 14773
rect 21082 14764 21088 14816
rect 21140 14804 21146 14816
rect 21177 14807 21235 14813
rect 21177 14804 21189 14807
rect 21140 14776 21189 14804
rect 21140 14764 21146 14776
rect 21177 14773 21189 14776
rect 21223 14773 21235 14807
rect 21634 14804 21640 14816
rect 21595 14776 21640 14804
rect 21177 14767 21235 14773
rect 21634 14764 21640 14776
rect 21692 14764 21698 14816
rect 21818 14804 21824 14816
rect 21779 14776 21824 14804
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 24397 14807 24455 14813
rect 24397 14804 24409 14807
rect 24268 14776 24409 14804
rect 24268 14764 24274 14776
rect 24397 14773 24409 14776
rect 24443 14773 24455 14807
rect 24397 14767 24455 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 2593 14603 2651 14609
rect 2593 14600 2605 14603
rect 1544 14572 2605 14600
rect 1544 14560 1550 14572
rect 2593 14569 2605 14572
rect 2639 14569 2651 14603
rect 2593 14563 2651 14569
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 4120 14572 4169 14600
rect 4120 14560 4126 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 6730 14600 6736 14612
rect 6691 14572 6736 14600
rect 4157 14563 4215 14569
rect 6730 14560 6736 14572
rect 6788 14560 6794 14612
rect 8846 14600 8852 14612
rect 8588 14572 8852 14600
rect 1765 14535 1823 14541
rect 1765 14501 1777 14535
rect 1811 14532 1823 14535
rect 2314 14532 2320 14544
rect 1811 14504 2320 14532
rect 1811 14501 1823 14504
rect 1765 14495 1823 14501
rect 2314 14492 2320 14504
rect 2372 14492 2378 14544
rect 7561 14535 7619 14541
rect 7561 14501 7573 14535
rect 7607 14532 7619 14535
rect 7929 14535 7987 14541
rect 7929 14532 7941 14535
rect 7607 14504 7941 14532
rect 7607 14501 7619 14504
rect 7561 14495 7619 14501
rect 7929 14501 7941 14504
rect 7975 14532 7987 14535
rect 8588 14532 8616 14572
rect 8846 14560 8852 14572
rect 8904 14600 8910 14612
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8904 14572 9137 14600
rect 8904 14560 8910 14572
rect 9125 14569 9137 14572
rect 9171 14600 9183 14603
rect 9306 14600 9312 14612
rect 9171 14572 9312 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9674 14600 9680 14612
rect 9539 14572 9680 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9674 14560 9680 14572
rect 9732 14600 9738 14612
rect 10686 14600 10692 14612
rect 9732 14572 10692 14600
rect 9732 14560 9738 14572
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 11624 14572 12909 14600
rect 7975 14504 8616 14532
rect 7975 14501 7987 14504
rect 7929 14495 7987 14501
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2424 14436 2973 14464
rect 2424 14408 2452 14436
rect 2961 14433 2973 14436
rect 3007 14433 3019 14467
rect 4246 14464 4252 14476
rect 4207 14436 4252 14464
rect 2961 14427 3019 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4706 14464 4712 14476
rect 4667 14436 4712 14464
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 5074 14464 5080 14476
rect 5035 14436 5080 14464
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5442 14464 5448 14476
rect 5403 14436 5448 14464
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 6546 14464 6552 14476
rect 6507 14436 6552 14464
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7374 14464 7380 14476
rect 7055 14436 7380 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 2406 14396 2412 14408
rect 1719 14368 2412 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2866 14356 2872 14408
rect 2924 14396 2930 14408
rect 3513 14399 3571 14405
rect 3513 14396 3525 14399
rect 2924 14368 3525 14396
rect 2924 14356 2930 14368
rect 3513 14365 3525 14368
rect 3559 14396 3571 14399
rect 5092 14396 5120 14424
rect 3559 14368 5120 14396
rect 6365 14399 6423 14405
rect 3559 14365 3571 14368
rect 3513 14359 3571 14365
rect 6365 14365 6377 14399
rect 6411 14396 6423 14399
rect 7024 14396 7052 14427
rect 7374 14424 7380 14436
rect 7432 14464 7438 14476
rect 7576 14464 7604 14495
rect 8018 14464 8024 14476
rect 7432 14436 7604 14464
rect 7979 14436 8024 14464
rect 7432 14424 7438 14436
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8588 14473 8616 14504
rect 8757 14535 8815 14541
rect 8757 14501 8769 14535
rect 8803 14532 8815 14535
rect 9398 14532 9404 14544
rect 8803 14504 9404 14532
rect 8803 14501 8815 14504
rect 8757 14495 8815 14501
rect 9398 14492 9404 14504
rect 9456 14492 9462 14544
rect 10962 14492 10968 14544
rect 11020 14532 11026 14544
rect 11624 14532 11652 14572
rect 12897 14569 12909 14572
rect 12943 14600 12955 14603
rect 13262 14600 13268 14612
rect 12943 14572 13268 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 14274 14600 14280 14612
rect 14235 14572 14280 14600
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 14734 14600 14740 14612
rect 14695 14572 14740 14600
rect 14734 14560 14740 14572
rect 14792 14560 14798 14612
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 16761 14603 16819 14609
rect 16761 14600 16773 14603
rect 16540 14572 16773 14600
rect 16540 14560 16546 14572
rect 16761 14569 16773 14572
rect 16807 14569 16819 14603
rect 17402 14600 17408 14612
rect 17363 14572 17408 14600
rect 16761 14563 16819 14569
rect 12250 14532 12256 14544
rect 11020 14504 11652 14532
rect 12211 14504 12256 14532
rect 11020 14492 11026 14504
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 9836 14467 9894 14473
rect 9836 14433 9848 14467
rect 9882 14464 9894 14467
rect 10686 14464 10692 14476
rect 9882 14436 10088 14464
rect 10599 14436 10692 14464
rect 9882 14433 9894 14436
rect 9836 14427 9894 14433
rect 10060 14408 10088 14436
rect 10686 14424 10692 14436
rect 10744 14464 10750 14476
rect 10781 14467 10839 14473
rect 10781 14464 10793 14467
rect 10744 14436 10793 14464
rect 10744 14424 10750 14436
rect 10781 14433 10793 14436
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 6411 14368 7052 14396
rect 6411 14365 6423 14368
rect 6365 14359 6423 14365
rect 10042 14356 10048 14408
rect 10100 14356 10106 14408
rect 2130 14288 2136 14340
rect 2188 14328 2194 14340
rect 2225 14331 2283 14337
rect 2225 14328 2237 14331
rect 2188 14300 2237 14328
rect 2188 14288 2194 14300
rect 2225 14297 2237 14300
rect 2271 14328 2283 14331
rect 5534 14328 5540 14340
rect 2271 14300 5540 14328
rect 2271 14297 2283 14300
rect 2225 14291 2283 14297
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 8662 14288 8668 14340
rect 8720 14328 8726 14340
rect 11164 14328 11192 14504
rect 11514 14464 11520 14476
rect 11475 14436 11520 14464
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11624 14473 11652 14504
rect 12250 14492 12256 14504
rect 12308 14492 12314 14544
rect 12802 14492 12808 14544
rect 12860 14532 12866 14544
rect 13402 14535 13460 14541
rect 13402 14532 13414 14535
rect 12860 14504 13414 14532
rect 12860 14492 12866 14504
rect 13402 14501 13414 14504
rect 13448 14501 13460 14535
rect 15930 14532 15936 14544
rect 15891 14504 15936 14532
rect 13402 14495 13460 14501
rect 15930 14492 15936 14504
rect 15988 14492 15994 14544
rect 16776 14532 16804 14563
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 20717 14603 20775 14609
rect 20717 14569 20729 14603
rect 20763 14600 20775 14603
rect 21174 14600 21180 14612
rect 20763 14572 21180 14600
rect 20763 14569 20775 14572
rect 20717 14563 20775 14569
rect 21174 14560 21180 14572
rect 21232 14560 21238 14612
rect 22646 14600 22652 14612
rect 22607 14572 22652 14600
rect 22646 14560 22652 14572
rect 22704 14560 22710 14612
rect 23750 14600 23756 14612
rect 23711 14572 23756 14600
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 19705 14535 19763 14541
rect 16776 14504 19472 14532
rect 17788 14476 17816 14504
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14433 11667 14467
rect 11609 14427 11667 14433
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14433 12035 14467
rect 17310 14464 17316 14476
rect 17271 14436 17316 14464
rect 11977 14427 12035 14433
rect 11992 14396 12020 14427
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17770 14464 17776 14476
rect 17683 14436 17776 14464
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 18966 14464 18972 14476
rect 18927 14436 18972 14464
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 19444 14473 19472 14504
rect 19705 14501 19717 14535
rect 19751 14532 19763 14535
rect 19978 14532 19984 14544
rect 19751 14504 19984 14532
rect 19751 14501 19763 14504
rect 19705 14495 19763 14501
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 21082 14532 21088 14544
rect 20732 14504 21088 14532
rect 19429 14467 19487 14473
rect 19429 14433 19441 14467
rect 19475 14464 19487 14467
rect 20732 14464 20760 14504
rect 21082 14492 21088 14504
rect 21140 14532 21146 14544
rect 22186 14532 22192 14544
rect 21140 14504 22192 14532
rect 21140 14492 21146 14504
rect 19475 14436 20760 14464
rect 19475 14433 19487 14436
rect 19429 14427 19487 14433
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 21376 14473 21404 14504
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20864 14436 20913 14464
rect 20864 14424 20870 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 21361 14467 21419 14473
rect 21361 14433 21373 14467
rect 21407 14433 21419 14467
rect 21361 14427 21419 14433
rect 22465 14467 22523 14473
rect 22465 14433 22477 14467
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 13078 14396 13084 14408
rect 8720 14300 11192 14328
rect 11256 14368 12020 14396
rect 13039 14368 13084 14396
rect 8720 14288 8726 14300
rect 11256 14272 11284 14368
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14396 15899 14399
rect 16758 14396 16764 14408
rect 15887 14368 16764 14396
rect 15887 14365 15899 14368
rect 15841 14359 15899 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 21453 14399 21511 14405
rect 21453 14396 21465 14399
rect 19576 14368 21465 14396
rect 19576 14356 19582 14368
rect 21453 14365 21465 14368
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 14001 14331 14059 14337
rect 14001 14297 14013 14331
rect 14047 14328 14059 14331
rect 14090 14328 14096 14340
rect 14047 14300 14096 14328
rect 14047 14297 14059 14300
rect 14001 14291 14059 14297
rect 14090 14288 14096 14300
rect 14148 14328 14154 14340
rect 15286 14328 15292 14340
rect 14148 14300 15292 14328
rect 14148 14288 14154 14300
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 16390 14328 16396 14340
rect 16351 14300 16396 14328
rect 16390 14288 16396 14300
rect 16448 14288 16454 14340
rect 20162 14288 20168 14340
rect 20220 14328 20226 14340
rect 22480 14328 22508 14427
rect 23474 14424 23480 14476
rect 23532 14464 23538 14476
rect 23569 14467 23627 14473
rect 23569 14464 23581 14467
rect 23532 14436 23581 14464
rect 23532 14424 23538 14436
rect 23569 14433 23581 14436
rect 23615 14433 23627 14467
rect 23569 14427 23627 14433
rect 22646 14328 22652 14340
rect 20220 14300 22652 14328
rect 20220 14288 20226 14300
rect 22646 14288 22652 14300
rect 22704 14288 22710 14340
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4246 14260 4252 14272
rect 3927 14232 4252 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 9907 14263 9965 14269
rect 9907 14229 9919 14263
rect 9953 14260 9965 14263
rect 10134 14260 10140 14272
rect 9953 14232 10140 14260
rect 9953 14229 9965 14232
rect 9907 14223 9965 14229
rect 10134 14220 10140 14232
rect 10192 14220 10198 14272
rect 10321 14263 10379 14269
rect 10321 14229 10333 14263
rect 10367 14260 10379 14263
rect 11238 14260 11244 14272
rect 10367 14232 11244 14260
rect 10367 14229 10379 14232
rect 10321 14223 10379 14229
rect 11238 14220 11244 14232
rect 11296 14220 11302 14272
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 12529 14263 12587 14269
rect 12529 14260 12541 14263
rect 11664 14232 12541 14260
rect 11664 14220 11670 14232
rect 12529 14229 12541 14232
rect 12575 14229 12587 14263
rect 12529 14223 12587 14229
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 21913 14263 21971 14269
rect 21913 14260 21925 14263
rect 21876 14232 21925 14260
rect 21876 14220 21882 14232
rect 21913 14229 21925 14232
rect 21959 14229 21971 14263
rect 21913 14223 21971 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2866 14056 2872 14068
rect 2827 14028 2872 14056
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 9585 14059 9643 14065
rect 9585 14025 9597 14059
rect 9631 14056 9643 14059
rect 10042 14056 10048 14068
rect 9631 14028 10048 14056
rect 9631 14025 9643 14028
rect 9585 14019 9643 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 15930 14056 15936 14068
rect 15611 14028 15936 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 16758 14056 16764 14068
rect 16719 14028 16764 14056
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 17310 14056 17316 14068
rect 17271 14028 17316 14056
rect 17310 14016 17316 14028
rect 17368 14016 17374 14068
rect 17770 14056 17776 14068
rect 17731 14028 17776 14056
rect 17770 14016 17776 14028
rect 17828 14056 17834 14068
rect 18417 14059 18475 14065
rect 18417 14056 18429 14059
rect 17828 14028 18429 14056
rect 17828 14016 17834 14028
rect 18417 14025 18429 14028
rect 18463 14025 18475 14059
rect 18417 14019 18475 14025
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 21140 14028 21373 14056
rect 21140 14016 21146 14028
rect 21361 14025 21373 14028
rect 21407 14025 21419 14059
rect 22646 14056 22652 14068
rect 22607 14028 22652 14056
rect 21361 14019 21419 14025
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 23474 14056 23480 14068
rect 23446 14016 23480 14056
rect 23532 14056 23538 14068
rect 24121 14059 24179 14065
rect 24121 14056 24133 14059
rect 23532 14028 24133 14056
rect 23532 14016 23538 14028
rect 24121 14025 24133 14028
rect 24167 14025 24179 14059
rect 24121 14019 24179 14025
rect 106 13948 112 14000
rect 164 13988 170 14000
rect 3145 13991 3203 13997
rect 3145 13988 3157 13991
rect 164 13960 3157 13988
rect 164 13948 170 13960
rect 3145 13957 3157 13960
rect 3191 13957 3203 13991
rect 3145 13951 3203 13957
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 4157 13991 4215 13997
rect 4157 13988 4169 13991
rect 3568 13960 4169 13988
rect 3568 13948 3574 13960
rect 4157 13957 4169 13960
rect 4203 13988 4215 13991
rect 5442 13988 5448 14000
rect 4203 13960 5448 13988
rect 4203 13957 4215 13960
rect 4157 13951 4215 13957
rect 5442 13948 5448 13960
rect 5500 13948 5506 14000
rect 11422 13988 11428 14000
rect 11383 13960 11428 13988
rect 11422 13948 11428 13960
rect 11480 13948 11486 14000
rect 17862 13988 17868 14000
rect 12912 13960 15148 13988
rect 1486 13920 1492 13932
rect 1447 13892 1492 13920
rect 1486 13880 1492 13892
rect 1544 13880 1550 13932
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 6546 13920 6552 13932
rect 6507 13892 6552 13920
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 11606 13920 11612 13932
rect 9876 13892 11612 13920
rect 9876 13864 9904 13892
rect 2958 13852 2964 13864
rect 2919 13824 2964 13852
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 4246 13852 4252 13864
rect 4207 13824 4252 13852
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4706 13852 4712 13864
rect 4667 13824 4712 13852
rect 4706 13812 4712 13824
rect 4764 13852 4770 13864
rect 4764 13824 5028 13852
rect 4764 13812 4770 13824
rect 1578 13784 1584 13796
rect 1539 13756 1584 13784
rect 1578 13744 1584 13756
rect 1636 13784 1642 13796
rect 2409 13787 2467 13793
rect 2409 13784 2421 13787
rect 1636 13756 2421 13784
rect 1636 13744 1642 13756
rect 2409 13753 2421 13756
rect 2455 13753 2467 13787
rect 2409 13747 2467 13753
rect 3789 13787 3847 13793
rect 3789 13753 3801 13787
rect 3835 13784 3847 13787
rect 5000 13784 5028 13824
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 5132 13824 5177 13852
rect 5132 13812 5138 13824
rect 5350 13812 5356 13864
rect 5408 13852 5414 13864
rect 5445 13855 5503 13861
rect 5445 13852 5457 13855
rect 5408 13824 5457 13852
rect 5408 13812 5414 13824
rect 5445 13821 5457 13824
rect 5491 13821 5503 13855
rect 5445 13815 5503 13821
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7190 13852 7196 13864
rect 7147 13824 7196 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7374 13852 7380 13864
rect 7335 13824 7380 13852
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 8665 13855 8723 13861
rect 8496 13824 8616 13852
rect 6089 13787 6147 13793
rect 6089 13784 6101 13787
rect 3835 13756 6101 13784
rect 3835 13753 3847 13756
rect 3789 13747 3847 13753
rect 6089 13753 6101 13756
rect 6135 13784 6147 13787
rect 8110 13784 8116 13796
rect 6135 13756 8116 13784
rect 6135 13753 6147 13756
rect 6089 13747 6147 13753
rect 8110 13744 8116 13756
rect 8168 13784 8174 13796
rect 8496 13784 8524 13824
rect 8168 13756 8524 13784
rect 8168 13744 8174 13756
rect 4338 13716 4344 13728
rect 4299 13688 4344 13716
rect 4338 13676 4344 13688
rect 4396 13676 4402 13728
rect 6914 13716 6920 13728
rect 6875 13688 6920 13716
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 8018 13716 8024 13728
rect 7979 13688 8024 13716
rect 8018 13676 8024 13688
rect 8076 13676 8082 13728
rect 8478 13716 8484 13728
rect 8439 13688 8484 13716
rect 8478 13676 8484 13688
rect 8536 13676 8542 13728
rect 8588 13716 8616 13824
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 8846 13852 8852 13864
rect 8711 13824 8745 13852
rect 8807 13824 8852 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 8680 13784 8708 13815
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9858 13852 9864 13864
rect 9819 13824 9864 13852
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 10520 13861 10548 13892
rect 11606 13880 11612 13892
rect 11664 13920 11670 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11664 13892 11805 13920
rect 11664 13880 11670 13892
rect 11793 13889 11805 13892
rect 11839 13920 11851 13923
rect 12912 13920 12940 13960
rect 11839 13892 12940 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 10008 13824 10057 13852
rect 10008 13812 10014 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13821 10563 13855
rect 11054 13852 11060 13864
rect 11015 13824 11060 13852
rect 10505 13815 10563 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11238 13852 11244 13864
rect 11199 13824 11244 13852
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 12434 13852 12440 13864
rect 12395 13824 12440 13852
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12912 13861 12940 13892
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 15120 13920 15148 13960
rect 15304 13960 17868 13988
rect 15304 13920 15332 13960
rect 17862 13948 17868 13960
rect 17920 13948 17926 14000
rect 19168 13960 19334 13988
rect 13136 13892 13814 13920
rect 15120 13892 15332 13920
rect 13136 13880 13142 13892
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 13262 13852 13268 13864
rect 13223 13824 13268 13852
rect 12897 13815 12955 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13630 13852 13636 13864
rect 13591 13824 13636 13852
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13786 13852 13814 13892
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15930 13920 15936 13932
rect 15436 13892 15936 13920
rect 15436 13880 15442 13892
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16390 13920 16396 13932
rect 16080 13892 16396 13920
rect 16080 13880 16086 13892
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13786 13824 13921 13852
rect 13909 13821 13921 13824
rect 13955 13852 13967 13855
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13955 13824 14197 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 14424 13824 15209 13852
rect 14424 13812 14430 13824
rect 15197 13821 15209 13824
rect 15243 13852 15255 13855
rect 15396 13852 15424 13880
rect 19168 13861 19196 13960
rect 19306 13920 19334 13960
rect 22002 13948 22008 14000
rect 22060 13988 22066 14000
rect 23446 13988 23474 14016
rect 22060 13960 23474 13988
rect 22060 13948 22066 13960
rect 23566 13948 23572 14000
rect 23624 13988 23630 14000
rect 24489 13991 24547 13997
rect 24489 13988 24501 13991
rect 23624 13960 24501 13988
rect 23624 13948 23630 13960
rect 24489 13957 24501 13960
rect 24535 13957 24547 13991
rect 24489 13951 24547 13957
rect 20070 13920 20076 13932
rect 19306 13892 20076 13920
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 23799 13923 23857 13929
rect 23799 13920 23811 13923
rect 20180 13892 23811 13920
rect 15243 13824 15424 13852
rect 18877 13855 18935 13861
rect 15243 13821 15255 13824
rect 15197 13815 15255 13821
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 19153 13855 19211 13861
rect 19153 13852 19165 13855
rect 18923 13824 19165 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 19153 13821 19165 13824
rect 19199 13821 19211 13855
rect 19426 13852 19432 13864
rect 19387 13824 19432 13852
rect 19153 13815 19211 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20180 13852 20208 13892
rect 23799 13889 23811 13892
rect 23845 13889 23857 13923
rect 23799 13883 23857 13889
rect 19628 13824 20208 13852
rect 9030 13784 9036 13796
rect 8680 13756 9036 13784
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 14829 13787 14887 13793
rect 14829 13753 14841 13787
rect 14875 13784 14887 13787
rect 15749 13787 15807 13793
rect 15749 13784 15761 13787
rect 14875 13756 15761 13784
rect 14875 13753 14887 13756
rect 14829 13747 14887 13753
rect 15749 13753 15761 13756
rect 15795 13753 15807 13787
rect 15749 13747 15807 13753
rect 15841 13787 15899 13793
rect 15841 13753 15853 13787
rect 15887 13784 15899 13787
rect 15930 13784 15936 13796
rect 15887 13756 15936 13784
rect 15887 13753 15899 13756
rect 15841 13747 15899 13753
rect 9858 13716 9864 13728
rect 8588 13688 9864 13716
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 12250 13716 12256 13728
rect 12211 13688 12256 13716
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 15764 13716 15792 13747
rect 15930 13744 15936 13756
rect 15988 13744 15994 13796
rect 19628 13784 19656 13824
rect 22738 13812 22744 13864
rect 22796 13852 22802 13864
rect 23566 13852 23572 13864
rect 22796 13824 23572 13852
rect 22796 13812 22802 13824
rect 23566 13812 23572 13824
rect 23624 13852 23630 13864
rect 23696 13855 23754 13861
rect 23696 13852 23708 13855
rect 23624 13824 23708 13852
rect 23624 13812 23630 13824
rect 23696 13821 23708 13824
rect 23742 13821 23754 13855
rect 23696 13815 23754 13821
rect 18202 13756 19656 13784
rect 19705 13787 19763 13793
rect 18202 13716 18230 13756
rect 19705 13753 19717 13787
rect 19751 13784 19763 13787
rect 19886 13784 19892 13796
rect 19751 13756 19892 13784
rect 19751 13753 19763 13756
rect 19705 13747 19763 13753
rect 19886 13744 19892 13756
rect 19944 13744 19950 13796
rect 20070 13744 20076 13796
rect 20128 13784 20134 13796
rect 21729 13787 21787 13793
rect 20128 13756 20852 13784
rect 20128 13744 20134 13756
rect 20824 13728 20852 13756
rect 21729 13753 21741 13787
rect 21775 13753 21787 13787
rect 21729 13747 21787 13753
rect 20530 13716 20536 13728
rect 15764 13688 18230 13716
rect 20491 13688 20536 13716
rect 20530 13676 20536 13688
rect 20588 13676 20594 13728
rect 20806 13676 20812 13728
rect 20864 13716 20870 13728
rect 20993 13719 21051 13725
rect 20993 13716 21005 13719
rect 20864 13688 21005 13716
rect 20864 13676 20870 13688
rect 20993 13685 21005 13688
rect 21039 13685 21051 13719
rect 21744 13716 21772 13747
rect 21818 13744 21824 13796
rect 21876 13784 21882 13796
rect 21876 13756 21921 13784
rect 21876 13744 21882 13756
rect 22186 13744 22192 13796
rect 22244 13784 22250 13796
rect 22373 13787 22431 13793
rect 22373 13784 22385 13787
rect 22244 13756 22385 13784
rect 22244 13744 22250 13756
rect 22373 13753 22385 13756
rect 22419 13753 22431 13787
rect 22373 13747 22431 13753
rect 22278 13716 22284 13728
rect 21744 13688 22284 13716
rect 20993 13679 21051 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2409 13515 2467 13521
rect 2409 13512 2421 13515
rect 2372 13484 2421 13512
rect 2372 13472 2378 13484
rect 2409 13481 2421 13484
rect 2455 13512 2467 13515
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2455 13484 2697 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 4157 13515 4215 13521
rect 4157 13512 4169 13515
rect 3476 13484 4169 13512
rect 3476 13472 3482 13484
rect 4157 13481 4169 13484
rect 4203 13481 4215 13515
rect 4157 13475 4215 13481
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7432 13484 7849 13512
rect 7432 13472 7438 13484
rect 7837 13481 7849 13484
rect 7883 13481 7895 13515
rect 9030 13512 9036 13524
rect 8991 13484 9036 13512
rect 7837 13475 7895 13481
rect 1670 13404 1676 13456
rect 1728 13444 1734 13456
rect 1810 13447 1868 13453
rect 1810 13444 1822 13447
rect 1728 13416 1822 13444
rect 1728 13404 1734 13416
rect 1810 13413 1822 13416
rect 1856 13413 1868 13447
rect 1810 13407 1868 13413
rect 6454 13404 6460 13456
rect 6512 13444 6518 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 6512 13416 6561 13444
rect 6512 13404 6518 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 7098 13444 7104 13456
rect 7059 13416 7104 13444
rect 6549 13407 6607 13413
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 7852 13444 7880 13475
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 9364 13484 10793 13512
rect 9364 13472 9370 13484
rect 10781 13481 10793 13484
rect 10827 13512 10839 13515
rect 11422 13512 11428 13524
rect 10827 13484 11428 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 12066 13512 12072 13524
rect 12027 13484 12072 13512
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12621 13515 12679 13521
rect 12621 13512 12633 13515
rect 12492 13484 12633 13512
rect 12492 13472 12498 13484
rect 12621 13481 12633 13484
rect 12667 13481 12679 13515
rect 12621 13475 12679 13481
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 12860 13484 13093 13512
rect 12860 13472 12866 13484
rect 13081 13481 13093 13484
rect 13127 13481 13139 13515
rect 14366 13512 14372 13524
rect 14327 13484 14372 13512
rect 13081 13475 13139 13481
rect 8754 13444 8760 13456
rect 7852 13416 8524 13444
rect 8715 13416 8760 13444
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13376 3571 13379
rect 4338 13376 4344 13388
rect 3559 13348 4344 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 4338 13336 4344 13348
rect 4396 13336 4402 13388
rect 4522 13376 4528 13388
rect 4483 13348 4528 13376
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 5074 13376 5080 13388
rect 5035 13348 5080 13376
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 5534 13376 5540 13388
rect 5491 13348 5540 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 8496 13385 8524 13416
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 12452 13444 12480 13472
rect 11164 13416 12480 13444
rect 13096 13444 13124 13475
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 19426 13512 19432 13524
rect 19387 13484 19432 13512
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 13814 13453 13820 13456
rect 13770 13447 13820 13453
rect 13770 13444 13782 13447
rect 13096 13416 13782 13444
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 8481 13379 8539 13385
rect 8343 13348 8432 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13308 1547 13311
rect 3053 13311 3111 13317
rect 3053 13308 3065 13311
rect 1535 13280 3065 13308
rect 1535 13277 1547 13280
rect 1489 13271 1547 13277
rect 3053 13277 3065 13280
rect 3099 13308 3111 13311
rect 3694 13308 3700 13320
rect 3099 13280 3700 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3694 13268 3700 13280
rect 3752 13268 3758 13320
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 8404 13308 8432 13348
rect 8481 13345 8493 13379
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10008 13348 10425 13376
rect 10008 13336 10014 13348
rect 10413 13345 10425 13348
rect 10459 13376 10471 13379
rect 10686 13376 10692 13388
rect 10459 13348 10692 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 10686 13336 10692 13348
rect 10744 13376 10750 13388
rect 10962 13376 10968 13388
rect 10744 13348 10968 13376
rect 10744 13336 10750 13348
rect 10962 13336 10968 13348
rect 11020 13376 11026 13388
rect 11164 13385 11192 13416
rect 13770 13413 13782 13416
rect 13816 13413 13820 13447
rect 13770 13407 13820 13413
rect 13814 13404 13820 13407
rect 13872 13404 13878 13456
rect 13906 13404 13912 13456
rect 13964 13444 13970 13456
rect 15289 13447 15347 13453
rect 15289 13444 15301 13447
rect 13964 13416 15301 13444
rect 13964 13404 13970 13416
rect 15289 13413 15301 13416
rect 15335 13413 15347 13447
rect 18138 13444 18144 13456
rect 18099 13416 18144 13444
rect 15289 13407 15347 13413
rect 18138 13404 18144 13416
rect 18196 13404 18202 13456
rect 21450 13444 21456 13456
rect 21411 13416 21456 13444
rect 21450 13404 21456 13416
rect 21508 13404 21514 13456
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 11020 13348 11161 13376
rect 11020 13336 11026 13348
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 11606 13376 11612 13388
rect 11567 13348 11612 13376
rect 11149 13339 11207 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13345 11759 13379
rect 12250 13376 12256 13388
rect 12211 13348 12256 13376
rect 11701 13339 11759 13345
rect 9398 13308 9404 13320
rect 8404 13280 9404 13308
rect 6457 13271 6515 13277
rect 5905 13243 5963 13249
rect 5905 13209 5917 13243
rect 5951 13240 5963 13243
rect 6472 13240 6500 13271
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 11514 13308 11520 13320
rect 9907 13280 11520 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 7006 13240 7012 13252
rect 5951 13212 6408 13240
rect 6472 13212 7012 13240
rect 5951 13209 5963 13212
rect 5905 13203 5963 13209
rect 3786 13172 3792 13184
rect 3747 13144 3792 13172
rect 3786 13132 3792 13144
rect 3844 13172 3850 13184
rect 5350 13172 5356 13184
rect 3844 13144 5356 13172
rect 3844 13132 3850 13144
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 6270 13172 6276 13184
rect 6231 13144 6276 13172
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 6380 13172 6408 13212
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 11054 13240 11060 13252
rect 9416 13212 11060 13240
rect 6914 13172 6920 13184
rect 6380 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 7248 13144 7481 13172
rect 7248 13132 7254 13144
rect 7469 13141 7481 13144
rect 7515 13172 7527 13175
rect 7742 13172 7748 13184
rect 7515 13144 7748 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 9416 13181 9444 13212
rect 11054 13200 11060 13212
rect 11112 13240 11118 13252
rect 11710 13240 11738 13339
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 15378 13376 15384 13388
rect 15339 13348 15384 13376
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 16850 13376 16856 13388
rect 16811 13348 16856 13376
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 19518 13376 19524 13388
rect 18748 13348 19524 13376
rect 18748 13336 18754 13348
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 24670 13385 24676 13388
rect 24648 13379 24676 13385
rect 24648 13376 24660 13379
rect 24583 13348 24660 13376
rect 24648 13345 24660 13348
rect 24728 13376 24734 13388
rect 26234 13376 26240 13388
rect 24728 13348 26240 13376
rect 24648 13339 24676 13345
rect 24670 13336 24676 13339
rect 24728 13336 24734 13348
rect 26234 13336 26240 13348
rect 26292 13336 26298 13388
rect 13446 13308 13452 13320
rect 13407 13280 13452 13308
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 18049 13311 18107 13317
rect 18049 13277 18061 13311
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 21361 13311 21419 13317
rect 21361 13277 21373 13311
rect 21407 13308 21419 13311
rect 22462 13308 22468 13320
rect 21407 13280 22468 13308
rect 21407 13277 21419 13280
rect 21361 13271 21419 13277
rect 11112 13212 11738 13240
rect 11112 13200 11118 13212
rect 16206 13200 16212 13252
rect 16264 13240 16270 13252
rect 17773 13243 17831 13249
rect 17773 13240 17785 13243
rect 16264 13212 17785 13240
rect 16264 13200 16270 13212
rect 17773 13209 17785 13212
rect 17819 13240 17831 13243
rect 18064 13240 18092 13271
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 18414 13240 18420 13252
rect 17819 13212 18420 13240
rect 17819 13209 17831 13212
rect 17773 13203 17831 13209
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 18598 13240 18604 13252
rect 18559 13212 18604 13240
rect 18598 13200 18604 13212
rect 18656 13240 18662 13252
rect 21910 13240 21916 13252
rect 18656 13212 21916 13240
rect 18656 13200 18662 13212
rect 21910 13200 21916 13212
rect 21968 13200 21974 13252
rect 9401 13175 9459 13181
rect 9401 13172 9413 13175
rect 9272 13144 9413 13172
rect 9272 13132 9278 13144
rect 9401 13141 9413 13144
rect 9447 13141 9459 13175
rect 9401 13135 9459 13141
rect 16991 13175 17049 13181
rect 16991 13141 17003 13175
rect 17037 13172 17049 13175
rect 17126 13172 17132 13184
rect 17037 13144 17132 13172
rect 17037 13141 17049 13144
rect 16991 13135 17049 13141
rect 17126 13132 17132 13144
rect 17184 13132 17190 13184
rect 19058 13172 19064 13184
rect 19019 13144 19064 13172
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 19702 13172 19708 13184
rect 19663 13144 19708 13172
rect 19702 13132 19708 13144
rect 19760 13132 19766 13184
rect 22278 13172 22284 13184
rect 22239 13144 22284 13172
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 22370 13132 22376 13184
rect 22428 13172 22434 13184
rect 24719 13175 24777 13181
rect 24719 13172 24731 13175
rect 22428 13144 24731 13172
rect 22428 13132 22434 13144
rect 24719 13141 24731 13144
rect 24765 13141 24777 13175
rect 24719 13135 24777 13141
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 1673 12971 1731 12977
rect 1673 12968 1685 12971
rect 1636 12940 1685 12968
rect 1636 12928 1642 12940
rect 1673 12937 1685 12940
rect 1719 12937 1731 12971
rect 3510 12968 3516 12980
rect 3471 12940 3516 12968
rect 1673 12931 1731 12937
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5132 12940 5825 12968
rect 5132 12928 5138 12940
rect 5813 12937 5825 12940
rect 5859 12968 5871 12971
rect 6178 12968 6184 12980
rect 5859 12940 6184 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 6178 12928 6184 12940
rect 6236 12968 6242 12980
rect 8662 12968 8668 12980
rect 6236 12940 8668 12968
rect 6236 12928 6242 12940
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11606 12968 11612 12980
rect 11563 12940 11612 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 14185 12971 14243 12977
rect 14185 12968 14197 12971
rect 13872 12940 14197 12968
rect 13872 12928 13878 12940
rect 14185 12937 14197 12940
rect 14231 12968 14243 12971
rect 14734 12968 14740 12980
rect 14231 12940 14740 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 15378 12968 15384 12980
rect 15339 12940 15384 12968
rect 15378 12928 15384 12940
rect 15436 12928 15442 12980
rect 16850 12968 16856 12980
rect 16811 12940 16856 12968
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17497 12971 17555 12977
rect 17497 12937 17509 12971
rect 17543 12968 17555 12971
rect 18138 12968 18144 12980
rect 17543 12940 18144 12968
rect 17543 12937 17555 12940
rect 17497 12931 17555 12937
rect 18138 12928 18144 12940
rect 18196 12968 18202 12980
rect 18969 12971 19027 12977
rect 18969 12968 18981 12971
rect 18196 12940 18981 12968
rect 18196 12928 18202 12940
rect 18969 12937 18981 12940
rect 19015 12937 19027 12971
rect 18969 12931 19027 12937
rect 20993 12971 21051 12977
rect 20993 12937 21005 12971
rect 21039 12968 21051 12971
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 21039 12940 21373 12968
rect 21039 12937 21051 12940
rect 20993 12931 21051 12937
rect 21361 12937 21373 12940
rect 21407 12968 21419 12971
rect 21450 12968 21456 12980
rect 21407 12940 21456 12968
rect 21407 12937 21419 12940
rect 21361 12931 21419 12937
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24670 12968 24676 12980
rect 24535 12940 24676 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 24765 12971 24823 12977
rect 24765 12937 24777 12971
rect 24811 12968 24823 12971
rect 24854 12968 24860 12980
rect 24811 12940 24860 12968
rect 24811 12937 24823 12940
rect 24765 12931 24823 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 4522 12832 4528 12844
rect 2823 12804 4528 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 2038 12764 2044 12776
rect 1951 12736 2044 12764
rect 2038 12724 2044 12736
rect 2096 12764 2102 12776
rect 2314 12764 2320 12776
rect 2096 12736 2320 12764
rect 2096 12724 2102 12736
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 4172 12773 4200 12804
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 5092 12832 5120 12928
rect 5718 12860 5724 12912
rect 5776 12900 5782 12912
rect 7837 12903 7895 12909
rect 7837 12900 7849 12903
rect 5776 12872 7849 12900
rect 5776 12860 5782 12872
rect 7837 12869 7849 12872
rect 7883 12900 7895 12903
rect 8386 12900 8392 12912
rect 7883 12872 8392 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8386 12860 8392 12872
rect 8444 12900 8450 12912
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 8444 12872 8493 12900
rect 8444 12860 8450 12872
rect 8481 12869 8493 12872
rect 8527 12869 8539 12903
rect 8754 12900 8760 12912
rect 8481 12863 8539 12869
rect 8588 12872 8760 12900
rect 6914 12832 6920 12844
rect 4632 12804 5120 12832
rect 6875 12804 6920 12832
rect 4632 12776 4660 12804
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 7156 12804 7205 12832
rect 7156 12792 7162 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4614 12764 4620 12776
rect 4527 12736 4620 12764
rect 4157 12727 4215 12733
rect 3145 12699 3203 12705
rect 3145 12665 3157 12699
rect 3191 12696 3203 12699
rect 3896 12696 3924 12727
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5350 12764 5356 12776
rect 5031 12736 5356 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 8588 12764 8616 12872
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 11149 12903 11207 12909
rect 11149 12900 11161 12903
rect 8996 12872 11161 12900
rect 8996 12860 9002 12872
rect 11149 12869 11161 12872
rect 11195 12900 11207 12903
rect 12250 12900 12256 12912
rect 11195 12872 12256 12900
rect 11195 12869 11207 12872
rect 11149 12863 11207 12869
rect 12250 12860 12256 12872
rect 12308 12900 12314 12912
rect 13630 12900 13636 12912
rect 12308 12872 13636 12900
rect 12308 12860 12314 12872
rect 13630 12860 13636 12872
rect 13688 12860 13694 12912
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 21818 12900 21824 12912
rect 15988 12872 21824 12900
rect 15988 12860 15994 12872
rect 21818 12860 21824 12872
rect 21876 12860 21882 12912
rect 8846 12832 8852 12844
rect 8807 12804 8852 12832
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13044 12804 13308 12832
rect 13044 12792 13050 12804
rect 8435 12736 8616 12764
rect 8665 12767 8723 12773
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8665 12733 8677 12767
rect 8711 12733 8723 12767
rect 10686 12764 10692 12776
rect 10647 12736 10692 12764
rect 8665 12727 8723 12733
rect 3191 12668 3924 12696
rect 3191 12665 3203 12668
rect 3145 12659 3203 12665
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2866 12628 2872 12640
rect 2464 12600 2872 12628
rect 2464 12588 2470 12600
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3694 12628 3700 12640
rect 3655 12600 3700 12628
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 3896 12628 3924 12668
rect 6270 12656 6276 12708
rect 6328 12696 6334 12708
rect 7009 12699 7067 12705
rect 7009 12696 7021 12699
rect 6328 12668 7021 12696
rect 6328 12656 6334 12668
rect 7009 12665 7021 12668
rect 7055 12696 7067 12699
rect 7098 12696 7104 12708
rect 7055 12668 7104 12696
rect 7055 12665 7067 12668
rect 7009 12659 7067 12665
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 4338 12628 4344 12640
rect 3896 12600 4344 12628
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 5353 12631 5411 12637
rect 5353 12628 5365 12631
rect 4580 12600 5365 12628
rect 4580 12588 4586 12600
rect 5353 12597 5365 12600
rect 5399 12628 5411 12631
rect 5718 12628 5724 12640
rect 5399 12600 5724 12628
rect 5399 12597 5411 12600
rect 5353 12591 5411 12597
rect 5718 12588 5724 12600
rect 5776 12588 5782 12640
rect 6362 12628 6368 12640
rect 6323 12600 6368 12628
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 8018 12588 8024 12640
rect 8076 12628 8082 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 8076 12600 8217 12628
rect 8076 12588 8082 12600
rect 8205 12597 8217 12600
rect 8251 12628 8263 12631
rect 8680 12628 8708 12727
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 12434 12764 12440 12776
rect 12395 12736 12440 12764
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 13078 12764 13084 12776
rect 13039 12736 13084 12764
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13280 12773 13308 12804
rect 13446 12792 13452 12844
rect 13504 12832 13510 12844
rect 15565 12835 15623 12841
rect 13504 12804 13814 12832
rect 13504 12792 13510 12804
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12733 13323 12767
rect 13630 12764 13636 12776
rect 13591 12736 13636 12764
rect 13265 12727 13323 12733
rect 13630 12724 13636 12736
rect 13688 12724 13694 12776
rect 9214 12656 9220 12708
rect 9272 12696 9278 12708
rect 9861 12699 9919 12705
rect 9861 12696 9873 12699
rect 9272 12668 9873 12696
rect 9272 12656 9278 12668
rect 9861 12665 9873 12668
rect 9907 12665 9919 12699
rect 10042 12696 10048 12708
rect 10003 12668 10048 12696
rect 9861 12659 9919 12665
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 11885 12699 11943 12705
rect 11885 12696 11897 12699
rect 10836 12668 11897 12696
rect 10836 12656 10842 12668
rect 11885 12665 11897 12668
rect 11931 12696 11943 12699
rect 13096 12696 13124 12724
rect 11931 12668 13124 12696
rect 13786 12696 13814 12804
rect 15565 12801 15577 12835
rect 15611 12832 15623 12835
rect 16485 12835 16543 12841
rect 16485 12832 16497 12835
rect 15611 12804 16497 12832
rect 15611 12801 15623 12804
rect 15565 12795 15623 12801
rect 16485 12801 16497 12804
rect 16531 12832 16543 12835
rect 16574 12832 16580 12844
rect 16531 12804 16580 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12832 19855 12835
rect 20346 12832 20352 12844
rect 19843 12804 20352 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 20346 12792 20352 12804
rect 20404 12832 20410 12844
rect 20404 12792 20437 12832
rect 18049 12767 18107 12773
rect 18049 12733 18061 12767
rect 18095 12764 18107 12767
rect 18598 12764 18604 12776
rect 18095 12736 18604 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 18598 12724 18604 12736
rect 18656 12724 18662 12776
rect 20070 12764 20076 12776
rect 20031 12736 20076 12764
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 13909 12699 13967 12705
rect 13909 12696 13921 12699
rect 13786 12668 13921 12696
rect 11931 12665 11943 12668
rect 11885 12659 11943 12665
rect 13909 12665 13921 12668
rect 13955 12696 13967 12699
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 13955 12668 14565 12696
rect 13955 12665 13967 12668
rect 13909 12659 13967 12665
rect 14553 12665 14565 12668
rect 14599 12665 14611 12699
rect 14553 12659 14611 12665
rect 15013 12699 15071 12705
rect 15013 12665 15025 12699
rect 15059 12696 15071 12699
rect 15657 12699 15715 12705
rect 15657 12696 15669 12699
rect 15059 12668 15669 12696
rect 15059 12665 15071 12668
rect 15013 12659 15071 12665
rect 15657 12665 15669 12668
rect 15703 12696 15715 12699
rect 15930 12696 15936 12708
rect 15703 12668 15936 12696
rect 15703 12665 15715 12668
rect 15657 12659 15715 12665
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 16206 12696 16212 12708
rect 16167 12668 16212 12696
rect 16206 12656 16212 12668
rect 16264 12656 16270 12708
rect 18370 12699 18428 12705
rect 18370 12665 18382 12699
rect 18416 12665 18428 12699
rect 18370 12659 18428 12665
rect 8251 12600 8708 12628
rect 8251 12597 8263 12600
rect 8205 12591 8263 12597
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17460 12600 17785 12628
rect 17460 12588 17466 12600
rect 17773 12597 17785 12600
rect 17819 12628 17831 12631
rect 18385 12628 18413 12659
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 20409 12705 20437 12792
rect 19613 12699 19671 12705
rect 19613 12696 19625 12699
rect 19576 12668 19625 12696
rect 19576 12656 19582 12668
rect 19613 12665 19625 12668
rect 19659 12696 19671 12699
rect 20394 12699 20452 12705
rect 19659 12668 20024 12696
rect 19659 12665 19671 12668
rect 19613 12659 19671 12665
rect 19334 12628 19340 12640
rect 17819 12600 19340 12628
rect 17819 12597 17831 12600
rect 17773 12591 17831 12597
rect 19334 12588 19340 12600
rect 19392 12628 19398 12640
rect 19797 12631 19855 12637
rect 19797 12628 19809 12631
rect 19392 12600 19809 12628
rect 19392 12588 19398 12600
rect 19797 12597 19809 12600
rect 19843 12628 19855 12631
rect 19889 12631 19947 12637
rect 19889 12628 19901 12631
rect 19843 12600 19901 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 19889 12597 19901 12600
rect 19935 12597 19947 12631
rect 19996 12628 20024 12668
rect 20394 12665 20406 12699
rect 20440 12665 20452 12699
rect 21836 12696 21864 12860
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12832 22155 12835
rect 22370 12832 22376 12844
rect 22143 12804 22376 12832
rect 22143 12801 22155 12804
rect 22097 12795 22155 12801
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 22462 12792 22468 12844
rect 22520 12832 22526 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 22520 12804 23029 12832
rect 22520 12792 22526 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 23106 12724 23112 12776
rect 23164 12764 23170 12776
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 23164 12736 24593 12764
rect 23164 12724 23170 12736
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 22189 12699 22247 12705
rect 22189 12696 22201 12699
rect 21836 12668 22201 12696
rect 20394 12659 20452 12665
rect 22189 12665 22201 12668
rect 22235 12665 22247 12699
rect 24596 12696 24624 12727
rect 25222 12696 25228 12708
rect 24596 12668 25228 12696
rect 22189 12659 22247 12665
rect 25222 12656 25228 12668
rect 25280 12656 25286 12708
rect 22646 12628 22652 12640
rect 19996 12600 22652 12628
rect 19889 12591 19947 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 106 12384 112 12436
rect 164 12424 170 12436
rect 3697 12427 3755 12433
rect 164 12396 2636 12424
rect 164 12384 170 12396
rect 1670 12356 1676 12368
rect 1631 12328 1676 12356
rect 1670 12316 1676 12328
rect 1728 12316 1734 12368
rect 2038 12356 2044 12368
rect 1999 12328 2044 12356
rect 2038 12316 2044 12328
rect 2096 12316 2102 12368
rect 2498 12356 2504 12368
rect 2459 12328 2504 12356
rect 2498 12316 2504 12328
rect 2556 12316 2562 12368
rect 2608 12356 2636 12396
rect 3697 12393 3709 12427
rect 3743 12424 3755 12427
rect 3786 12424 3792 12436
rect 3743 12396 3792 12424
rect 3743 12393 3755 12396
rect 3697 12387 3755 12393
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 3896 12396 4261 12424
rect 3896 12356 3924 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 12434 12424 12440 12436
rect 4249 12387 4307 12393
rect 9876 12396 11468 12424
rect 12395 12396 12440 12424
rect 2608 12328 3924 12356
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 9876 12365 9904 12396
rect 11440 12368 11468 12396
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12897 12427 12955 12433
rect 12897 12393 12909 12427
rect 12943 12424 12955 12427
rect 12986 12424 12992 12436
rect 12943 12396 12992 12424
rect 12943 12393 12955 12396
rect 12897 12387 12955 12393
rect 12986 12384 12992 12396
rect 13044 12424 13050 12436
rect 13170 12424 13176 12436
rect 13044 12396 13176 12424
rect 13044 12384 13050 12396
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16209 12427 16267 12433
rect 16209 12424 16221 12427
rect 15988 12396 16221 12424
rect 15988 12384 15994 12396
rect 16209 12393 16221 12396
rect 16255 12393 16267 12427
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 16209 12387 16267 12393
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 18598 12424 18604 12436
rect 18559 12396 18604 12424
rect 18598 12384 18604 12396
rect 18656 12424 18662 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 18656 12396 18889 12424
rect 18656 12384 18662 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 21634 12424 21640 12436
rect 18877 12387 18935 12393
rect 18984 12396 21640 12424
rect 7882 12359 7940 12365
rect 7882 12356 7894 12359
rect 7340 12328 7894 12356
rect 7340 12316 7346 12328
rect 7882 12325 7894 12328
rect 7928 12325 7940 12359
rect 7882 12319 7940 12325
rect 9861 12359 9919 12365
rect 9861 12325 9873 12359
rect 9907 12325 9919 12359
rect 9861 12319 9919 12325
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 11330 12356 11336 12368
rect 10192 12328 11336 12356
rect 10192 12316 10198 12328
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 11422 12316 11428 12368
rect 11480 12356 11486 12368
rect 14458 12356 14464 12368
rect 11480 12328 11525 12356
rect 13740 12328 14464 12356
rect 11480 12316 11486 12328
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3568 12260 4077 12288
rect 3568 12248 3574 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 5537 12291 5595 12297
rect 5537 12257 5549 12291
rect 5583 12257 5595 12291
rect 5718 12288 5724 12300
rect 5679 12260 5724 12288
rect 5537 12251 5595 12257
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2455 12192 3280 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2958 12152 2964 12164
rect 2919 12124 2964 12152
rect 2958 12112 2964 12124
rect 3016 12112 3022 12164
rect 3252 12152 3280 12192
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4396 12192 4721 12220
rect 4396 12180 4402 12192
rect 4709 12189 4721 12192
rect 4755 12220 4767 12223
rect 5552 12220 5580 12251
rect 5718 12248 5724 12260
rect 5776 12288 5782 12300
rect 5994 12288 6000 12300
rect 5776 12260 6000 12288
rect 5776 12248 5782 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12288 6699 12291
rect 6914 12288 6920 12300
rect 6687 12260 6920 12288
rect 6687 12257 6699 12260
rect 6641 12251 6699 12257
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 7469 12291 7527 12297
rect 7469 12257 7481 12291
rect 7515 12288 7527 12291
rect 9214 12288 9220 12300
rect 7515 12260 9220 12288
rect 7515 12257 7527 12260
rect 7469 12251 7527 12257
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 10962 12288 10968 12300
rect 10923 12260 10968 12288
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 13740 12297 13768 12328
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 14734 12316 14740 12368
rect 14792 12356 14798 12368
rect 15610 12359 15668 12365
rect 15610 12356 15622 12359
rect 14792 12328 15622 12356
rect 14792 12316 14798 12328
rect 15610 12325 15622 12328
rect 15656 12325 15668 12359
rect 15610 12319 15668 12325
rect 18984 12300 19012 12396
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 22281 12427 22339 12433
rect 22281 12393 22293 12427
rect 22327 12424 22339 12427
rect 22370 12424 22376 12436
rect 22327 12396 22376 12424
rect 22327 12393 22339 12396
rect 22281 12387 22339 12393
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 21358 12356 21364 12368
rect 21319 12328 21364 12356
rect 21358 12316 21364 12328
rect 21416 12316 21422 12368
rect 21910 12356 21916 12368
rect 21871 12328 21916 12356
rect 21910 12316 21916 12328
rect 21968 12316 21974 12368
rect 22922 12356 22928 12368
rect 22883 12328 22928 12356
rect 22922 12316 22928 12328
rect 22980 12316 22986 12368
rect 24210 12316 24216 12368
rect 24268 12356 24274 12368
rect 24489 12359 24547 12365
rect 24489 12356 24501 12359
rect 24268 12328 24501 12356
rect 24268 12316 24274 12328
rect 24489 12325 24501 12328
rect 24535 12325 24547 12359
rect 24489 12319 24547 12325
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12257 13783 12291
rect 13725 12251 13783 12257
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12288 14243 12291
rect 17586 12288 17592 12300
rect 14231 12260 17592 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 6086 12220 6092 12232
rect 4755 12192 6092 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12220 6791 12223
rect 7561 12223 7619 12229
rect 7561 12220 7573 12223
rect 6779 12192 7573 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 7561 12189 7573 12192
rect 7607 12220 7619 12223
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 7607 12192 9137 12220
rect 7607 12189 7619 12192
rect 7561 12183 7619 12189
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12189 9827 12223
rect 10134 12220 10140 12232
rect 10095 12192 10140 12220
rect 9769 12183 9827 12189
rect 3326 12152 3332 12164
rect 3252 12124 3332 12152
rect 3326 12112 3332 12124
rect 3384 12112 3390 12164
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4126 12124 4997 12152
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 4126 12084 4154 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 4985 12115 5043 12121
rect 8202 12112 8208 12164
rect 8260 12152 8266 12164
rect 9784 12152 9812 12183
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12802 12220 12808 12232
rect 12023 12192 12808 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 14200 12220 14228 12251
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 18966 12288 18972 12300
rect 18927 12260 18972 12288
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 19337 12291 19395 12297
rect 19337 12257 19349 12291
rect 19383 12288 19395 12291
rect 19426 12288 19432 12300
rect 19383 12260 19432 12288
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 13786 12192 14228 12220
rect 14369 12223 14427 12229
rect 13786 12164 13814 12192
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 15289 12223 15347 12229
rect 15289 12220 15301 12223
rect 14415 12192 15301 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 15289 12189 15301 12192
rect 15335 12220 15347 12223
rect 16482 12220 16488 12232
rect 15335 12192 16488 12220
rect 15335 12189 15347 12192
rect 15289 12183 15347 12189
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 17034 12220 17040 12232
rect 16995 12192 17040 12220
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 21082 12180 21088 12232
rect 21140 12220 21146 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21140 12192 21281 12220
rect 21140 12180 21146 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 22830 12220 22836 12232
rect 22791 12192 22836 12220
rect 21269 12183 21327 12189
rect 10962 12152 10968 12164
rect 8260 12124 10968 12152
rect 8260 12112 8266 12124
rect 10962 12112 10968 12124
rect 11020 12112 11026 12164
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 13357 12155 13415 12161
rect 13357 12152 13369 12155
rect 12768 12124 13369 12152
rect 12768 12112 12774 12124
rect 13357 12121 13369 12124
rect 13403 12152 13415 12155
rect 13786 12152 13820 12164
rect 13403 12124 13820 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 21284 12152 21312 12183
rect 22830 12180 22836 12192
rect 22888 12180 22894 12232
rect 23109 12223 23167 12229
rect 23109 12189 23121 12223
rect 23155 12189 23167 12223
rect 23109 12183 23167 12189
rect 22186 12152 22192 12164
rect 21284 12124 22192 12152
rect 22186 12112 22192 12124
rect 22244 12152 22250 12164
rect 23124 12152 23152 12183
rect 24026 12180 24032 12232
rect 24084 12220 24090 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 24084 12192 24409 12220
rect 24084 12180 24090 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24673 12223 24731 12229
rect 24673 12220 24685 12223
rect 24397 12183 24455 12189
rect 24504 12192 24685 12220
rect 24504 12152 24532 12192
rect 24673 12189 24685 12192
rect 24719 12189 24731 12223
rect 24673 12183 24731 12189
rect 22244 12124 24532 12152
rect 22244 12112 22250 12124
rect 7006 12084 7012 12096
rect 1452 12056 4154 12084
rect 6967 12056 7012 12084
rect 1452 12044 1458 12056
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 8478 12084 8484 12096
rect 8439 12056 8484 12084
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 8846 12084 8852 12096
rect 8807 12056 8852 12084
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 16666 12084 16672 12096
rect 15712 12056 16672 12084
rect 15712 12044 15718 12056
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18230 12084 18236 12096
rect 18003 12056 18236 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 20070 12084 20076 12096
rect 20031 12056 20076 12084
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2133 11883 2191 11889
rect 2133 11849 2145 11883
rect 2179 11880 2191 11883
rect 2498 11880 2504 11892
rect 2179 11852 2504 11880
rect 2179 11849 2191 11852
rect 2133 11843 2191 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 4614 11880 4620 11892
rect 3743 11852 4620 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 7653 11883 7711 11889
rect 7653 11880 7665 11883
rect 5592 11852 7665 11880
rect 5592 11840 5598 11852
rect 7653 11849 7665 11852
rect 7699 11880 7711 11883
rect 8938 11880 8944 11892
rect 7699 11852 8944 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 10778 11880 10784 11892
rect 9447 11852 10784 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 11330 11840 11336 11892
rect 11388 11880 11394 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11388 11852 11989 11880
rect 11388 11840 11394 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 11977 11843 12035 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16482 11880 16488 11892
rect 16443 11852 16488 11880
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 20530 11880 20536 11892
rect 18156 11852 20536 11880
rect 2516 11812 2544 11840
rect 3973 11815 4031 11821
rect 3973 11812 3985 11815
rect 2516 11784 3985 11812
rect 3973 11781 3985 11784
rect 4019 11812 4031 11815
rect 4019 11784 4154 11812
rect 4019 11781 4031 11784
rect 3973 11775 4031 11781
rect 2958 11744 2964 11756
rect 2919 11716 2964 11744
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 4126 11676 4154 11784
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 6641 11815 6699 11821
rect 6641 11812 6653 11815
rect 6328 11784 6653 11812
rect 6328 11772 6334 11784
rect 6641 11781 6653 11784
rect 6687 11812 6699 11815
rect 13170 11812 13176 11824
rect 6687 11784 13176 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 13170 11772 13176 11784
rect 13228 11772 13234 11824
rect 15838 11812 15844 11824
rect 13648 11784 15844 11812
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 7006 11744 7012 11756
rect 5767 11716 7012 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7282 11744 7288 11756
rect 7243 11716 7288 11744
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 8404 11716 9413 11744
rect 8404 11688 8432 11716
rect 9401 11713 9413 11716
rect 9447 11744 9459 11747
rect 9493 11747 9551 11753
rect 9493 11744 9505 11747
rect 9447 11716 9505 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9493 11713 9505 11716
rect 9539 11713 9551 11747
rect 9493 11707 9551 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9861 11747 9919 11753
rect 9861 11744 9873 11747
rect 9732 11716 9873 11744
rect 9732 11704 9738 11716
rect 9861 11713 9873 11716
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 4126 11648 4261 11676
rect 4249 11645 4261 11648
rect 4295 11645 4307 11679
rect 8018 11676 8024 11688
rect 7979 11648 8024 11676
rect 4249 11639 4307 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8386 11676 8392 11688
rect 8347 11648 8392 11676
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11645 8815 11679
rect 8938 11676 8944 11688
rect 8899 11648 8944 11676
rect 8757 11639 8815 11645
rect 2682 11608 2688 11620
rect 2643 11580 2688 11608
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 2777 11611 2835 11617
rect 2777 11577 2789 11611
rect 2823 11577 2835 11611
rect 4157 11611 4215 11617
rect 4157 11608 4169 11611
rect 2777 11571 2835 11577
rect 3436 11580 4169 11608
rect 106 11500 112 11552
rect 164 11540 170 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 164 11512 1593 11540
rect 164 11500 170 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1581 11503 1639 11509
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2792 11540 2820 11571
rect 3436 11540 3464 11580
rect 4157 11577 4169 11580
rect 4203 11577 4215 11611
rect 4157 11571 4215 11577
rect 2547 11512 3464 11540
rect 5353 11543 5411 11549
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 5442 11540 5448 11552
rect 5399 11512 5448 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 6273 11543 6331 11549
rect 6273 11540 6285 11543
rect 6144 11512 6285 11540
rect 6144 11500 6150 11512
rect 6273 11509 6285 11512
rect 6319 11540 6331 11543
rect 8662 11540 8668 11552
rect 6319 11512 8668 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 8772 11540 8800 11639
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 9263 11648 10057 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 10045 11645 10057 11648
rect 10091 11676 10103 11679
rect 10870 11676 10876 11688
rect 10091 11648 10876 11676
rect 10091 11645 10103 11648
rect 10045 11639 10103 11645
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 13648 11685 13676 11784
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 18156 11756 18184 11852
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21269 11883 21327 11889
rect 21269 11880 21281 11883
rect 20947 11852 21281 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 21269 11849 21281 11852
rect 21315 11880 21327 11883
rect 21358 11880 21364 11892
rect 21315 11852 21364 11880
rect 21315 11849 21327 11852
rect 21269 11843 21327 11849
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 23382 11880 23388 11892
rect 22888 11852 23388 11880
rect 22888 11840 22894 11852
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 24026 11880 24032 11892
rect 23987 11852 24032 11880
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 24210 11840 24216 11892
rect 24268 11880 24274 11892
rect 24305 11883 24363 11889
rect 24305 11880 24317 11883
rect 24268 11852 24317 11880
rect 24268 11840 24274 11852
rect 24305 11849 24317 11852
rect 24351 11849 24363 11883
rect 24762 11880 24768 11892
rect 24723 11852 24768 11880
rect 24305 11843 24363 11849
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 18230 11772 18236 11824
rect 18288 11812 18294 11824
rect 21821 11815 21879 11821
rect 21821 11812 21833 11815
rect 18288 11784 21833 11812
rect 18288 11772 18294 11784
rect 21821 11781 21833 11784
rect 21867 11781 21879 11815
rect 21821 11775 21879 11781
rect 14458 11744 14464 11756
rect 14371 11716 14464 11744
rect 14458 11704 14464 11716
rect 14516 11744 14522 11756
rect 15930 11744 15936 11756
rect 14516 11716 15936 11744
rect 14516 11704 14522 11716
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 16807 11747 16865 11753
rect 16807 11744 16819 11747
rect 16632 11716 16819 11744
rect 16632 11704 16638 11716
rect 16807 11713 16819 11716
rect 16853 11713 16865 11747
rect 18138 11744 18144 11756
rect 18051 11716 18144 11744
rect 16807 11707 16865 11713
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 18414 11744 18420 11756
rect 18375 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 19426 11744 19432 11756
rect 19387 11716 19432 11744
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11676 13323 11679
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13311 11648 13645 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14093 11679 14151 11685
rect 13872 11648 13917 11676
rect 13872 11636 13878 11648
rect 14093 11645 14105 11679
rect 14139 11676 14151 11679
rect 14918 11676 14924 11688
rect 14139 11648 14924 11676
rect 14139 11645 14151 11648
rect 14093 11639 14151 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 16704 11679 16762 11685
rect 16704 11676 16716 11679
rect 15120 11648 16716 11676
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10366 11611 10424 11617
rect 10366 11608 10378 11611
rect 9732 11580 10378 11608
rect 9732 11568 9738 11580
rect 10366 11577 10378 11580
rect 10412 11577 10424 11611
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 10366 11571 10424 11577
rect 10980 11580 11345 11608
rect 9214 11540 9220 11552
rect 8772 11512 9220 11540
rect 9214 11500 9220 11512
rect 9272 11500 9278 11552
rect 10980 11549 11008 11580
rect 11333 11577 11345 11580
rect 11379 11608 11391 11611
rect 11422 11608 11428 11620
rect 11379 11580 11428 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 11422 11568 11428 11580
rect 11480 11608 11486 11620
rect 11701 11611 11759 11617
rect 11701 11608 11713 11611
rect 11480 11580 11713 11608
rect 11480 11568 11486 11580
rect 11701 11577 11713 11580
rect 11747 11608 11759 11611
rect 13446 11608 13452 11620
rect 11747 11580 13452 11608
rect 11747 11577 11759 11580
rect 11701 11571 11759 11577
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 13538 11568 13544 11620
rect 13596 11608 13602 11620
rect 15120 11608 15148 11648
rect 16704 11645 16716 11648
rect 16750 11676 16762 11679
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 16750 11648 17141 11676
rect 16750 11645 16762 11648
rect 16704 11639 16762 11645
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19797 11679 19855 11685
rect 19797 11676 19809 11679
rect 19392 11648 19809 11676
rect 19392 11636 19398 11648
rect 19797 11645 19809 11648
rect 19843 11645 19855 11679
rect 19797 11639 19855 11645
rect 13596 11580 15148 11608
rect 15242 11611 15300 11617
rect 13596 11568 13602 11580
rect 15242 11577 15254 11611
rect 15288 11608 15300 11611
rect 16022 11608 16028 11620
rect 15288 11580 16028 11608
rect 15288 11577 15300 11580
rect 15242 11571 15300 11577
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11509 11023 11543
rect 10965 11503 11023 11509
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12768 11512 12817 11540
rect 12768 11500 12774 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 15257 11540 15285 11571
rect 16022 11568 16028 11580
rect 16080 11608 16086 11620
rect 16117 11611 16175 11617
rect 16117 11608 16129 11611
rect 16080 11580 16129 11608
rect 16080 11568 16086 11580
rect 16117 11577 16129 11580
rect 16163 11608 16175 11611
rect 17402 11608 17408 11620
rect 16163 11580 17408 11608
rect 16163 11577 16175 11580
rect 16117 11571 16175 11577
rect 17402 11568 17408 11580
rect 17460 11608 17466 11620
rect 17497 11611 17555 11617
rect 17497 11608 17509 11611
rect 17460 11580 17509 11608
rect 17460 11568 17466 11580
rect 17497 11577 17509 11580
rect 17543 11577 17555 11611
rect 17497 11571 17555 11577
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 19812 11608 19840 11639
rect 20302 11611 20360 11617
rect 20302 11608 20314 11611
rect 18288 11580 18333 11608
rect 19812 11580 20314 11608
rect 18288 11568 18294 11580
rect 20302 11577 20314 11580
rect 20348 11577 20360 11611
rect 21836 11608 21864 11775
rect 22370 11772 22376 11824
rect 22428 11812 22434 11824
rect 24228 11812 24256 11840
rect 22428 11784 24256 11812
rect 22428 11772 22434 11784
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11744 22155 11747
rect 22186 11744 22192 11756
rect 22143 11716 22192 11744
rect 22143 11713 22155 11716
rect 22097 11707 22155 11713
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 22462 11744 22468 11756
rect 22423 11716 22468 11744
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 22922 11676 22928 11688
rect 22756 11648 22928 11676
rect 22189 11611 22247 11617
rect 22189 11608 22201 11611
rect 21836 11580 22201 11608
rect 20302 11571 20360 11577
rect 22189 11577 22201 11580
rect 22235 11608 22247 11611
rect 22756 11608 22784 11648
rect 22922 11636 22928 11648
rect 22980 11676 22986 11688
rect 23017 11679 23075 11685
rect 23017 11676 23029 11679
rect 22980 11648 23029 11676
rect 22980 11636 22986 11648
rect 23017 11645 23029 11648
rect 23063 11645 23075 11679
rect 24578 11676 24584 11688
rect 24491 11648 24584 11676
rect 23017 11639 23075 11645
rect 24578 11636 24584 11648
rect 24636 11676 24642 11688
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24636 11648 25145 11676
rect 24636 11636 24642 11648
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 22235 11580 22784 11608
rect 22235 11577 22247 11580
rect 22189 11571 22247 11577
rect 22830 11568 22836 11620
rect 22888 11608 22894 11620
rect 24026 11608 24032 11620
rect 22888 11580 24032 11608
rect 22888 11568 22894 11580
rect 24026 11568 24032 11580
rect 24084 11568 24090 11620
rect 14792 11512 15285 11540
rect 14792 11500 14798 11512
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 15841 11543 15899 11549
rect 15841 11540 15853 11543
rect 15712 11512 15853 11540
rect 15712 11500 15718 11512
rect 15841 11509 15853 11512
rect 15887 11509 15899 11543
rect 15841 11503 15899 11509
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 18966 11540 18972 11552
rect 18472 11512 18972 11540
rect 18472 11500 18478 11512
rect 18966 11500 18972 11512
rect 19024 11540 19030 11552
rect 19061 11543 19119 11549
rect 19061 11540 19073 11543
rect 19024 11512 19073 11540
rect 19024 11500 19030 11512
rect 19061 11509 19073 11512
rect 19107 11509 19119 11543
rect 19061 11503 19119 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 5905 11339 5963 11345
rect 4212 11308 4257 11336
rect 4212 11296 4218 11308
rect 5905 11305 5917 11339
rect 5951 11336 5963 11339
rect 5994 11336 6000 11348
rect 5951 11308 6000 11336
rect 5951 11305 5963 11308
rect 5905 11299 5963 11305
rect 1670 11228 1676 11280
rect 1728 11268 1734 11280
rect 2406 11268 2412 11280
rect 1728 11240 2412 11268
rect 1728 11228 1734 11240
rect 2406 11228 2412 11240
rect 2464 11268 2470 11280
rect 2546 11271 2604 11277
rect 2546 11268 2558 11271
rect 2464 11240 2558 11268
rect 2464 11228 2470 11240
rect 2546 11237 2558 11240
rect 2592 11237 2604 11271
rect 2546 11231 2604 11237
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 5920 11268 5948 11299
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6178 11336 6184 11348
rect 6139 11308 6184 11336
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 9033 11339 9091 11345
rect 9033 11305 9045 11339
rect 9079 11336 9091 11339
rect 9306 11336 9312 11348
rect 9079 11308 9312 11336
rect 9079 11305 9091 11308
rect 9033 11299 9091 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 10597 11339 10655 11345
rect 9732 11308 10063 11336
rect 9732 11296 9738 11308
rect 6362 11268 6368 11280
rect 3936 11240 5948 11268
rect 6323 11240 6368 11268
rect 3936 11228 3942 11240
rect 4816 11212 4844 11240
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 7098 11268 7104 11280
rect 7011 11240 7104 11268
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4798 11200 4804 11212
rect 4711 11172 4804 11200
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 4982 11200 4988 11212
rect 4943 11172 4988 11200
rect 4982 11160 4988 11172
rect 5040 11160 5046 11212
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11200 5503 11203
rect 5534 11200 5540 11212
rect 5491 11172 5540 11200
rect 5491 11169 5503 11172
rect 5445 11163 5503 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 7024 11209 7052 11240
rect 7098 11228 7104 11240
rect 7156 11268 7162 11280
rect 8478 11268 8484 11280
rect 7156 11240 8484 11268
rect 7156 11228 7162 11240
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 8662 11268 8668 11280
rect 8575 11240 8668 11268
rect 8662 11228 8668 11240
rect 8720 11268 8726 11280
rect 9858 11268 9864 11280
rect 8720 11240 9864 11268
rect 8720 11228 8726 11240
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 10035 11277 10063 11308
rect 10597 11305 10609 11339
rect 10643 11336 10655 11339
rect 10686 11336 10692 11348
rect 10643 11308 10692 11336
rect 10643 11305 10655 11308
rect 10597 11299 10655 11305
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 10870 11336 10876 11348
rect 10831 11308 10876 11336
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 11020 11308 12817 11336
rect 11020 11296 11026 11308
rect 12805 11305 12817 11308
rect 12851 11305 12863 11339
rect 14918 11336 14924 11348
rect 14879 11308 14924 11336
rect 12805 11299 12863 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16945 11339 17003 11345
rect 16945 11305 16957 11339
rect 16991 11336 17003 11339
rect 17034 11336 17040 11348
rect 16991 11308 17040 11336
rect 16991 11305 17003 11308
rect 16945 11299 17003 11305
rect 17034 11296 17040 11308
rect 17092 11336 17098 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 17092 11308 17141 11336
rect 17092 11296 17098 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 17129 11299 17187 11305
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 20441 11339 20499 11345
rect 20441 11336 20453 11339
rect 20036 11308 20453 11336
rect 20036 11296 20042 11308
rect 20441 11305 20453 11308
rect 20487 11305 20499 11339
rect 21082 11336 21088 11348
rect 21043 11308 21088 11336
rect 20441 11299 20499 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21407 11339 21465 11345
rect 21407 11305 21419 11339
rect 21453 11336 21465 11339
rect 22278 11336 22284 11348
rect 21453 11308 22284 11336
rect 21453 11305 21465 11308
rect 21407 11299 21465 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 23983 11339 24041 11345
rect 23983 11305 23995 11339
rect 24029 11336 24041 11339
rect 24578 11336 24584 11348
rect 24029 11308 24584 11336
rect 24029 11305 24041 11308
rect 23983 11299 24041 11305
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 10018 11271 10076 11277
rect 10018 11237 10030 11271
rect 10064 11237 10076 11271
rect 10704 11268 10732 11296
rect 11241 11271 11299 11277
rect 11241 11268 11253 11271
rect 10704 11240 11253 11268
rect 10018 11231 10076 11237
rect 11241 11237 11253 11240
rect 11287 11237 11299 11271
rect 11606 11268 11612 11280
rect 11567 11240 11612 11268
rect 11241 11231 11299 11237
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 15654 11268 15660 11280
rect 15615 11240 15660 11268
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 16206 11268 16212 11280
rect 16167 11240 16212 11268
rect 16206 11228 16212 11240
rect 16264 11228 16270 11280
rect 19797 11271 19855 11277
rect 17604 11240 19472 11268
rect 17604 11212 17632 11240
rect 19444 11212 19472 11240
rect 19797 11237 19809 11271
rect 19843 11268 19855 11271
rect 20070 11268 20076 11280
rect 19843 11240 20076 11268
rect 19843 11237 19855 11240
rect 19797 11231 19855 11237
rect 20070 11228 20076 11240
rect 20128 11228 20134 11280
rect 22370 11228 22376 11280
rect 22428 11268 22434 11280
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22428 11240 22477 11268
rect 22428 11228 22434 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11169 7067 11203
rect 8018 11200 8024 11212
rect 7009 11163 7067 11169
rect 7760 11172 8024 11200
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11132 2283 11135
rect 2774 11132 2780 11144
rect 2271 11104 2780 11132
rect 2271 11101 2283 11104
rect 2225 11095 2283 11101
rect 2774 11092 2780 11104
rect 2832 11092 2838 11144
rect 3881 11135 3939 11141
rect 3881 11101 3893 11135
rect 3927 11132 3939 11135
rect 5000 11132 5028 11160
rect 3927 11104 5028 11132
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 2498 11024 2504 11076
rect 2556 11064 2562 11076
rect 3145 11067 3203 11073
rect 3145 11064 3157 11067
rect 2556 11036 3157 11064
rect 2556 11024 2562 11036
rect 3145 11033 3157 11036
rect 3191 11033 3203 11067
rect 3145 11027 3203 11033
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 1946 10996 1952 11008
rect 1907 10968 1952 10996
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3384 10968 3433 10996
rect 3384 10956 3390 10968
rect 3421 10965 3433 10968
rect 3467 10965 3479 10999
rect 7466 10996 7472 11008
rect 7427 10968 7472 10996
rect 3421 10959 3479 10965
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 7760 11005 7788 11172
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 13446 11200 13452 11212
rect 13407 11172 13452 11200
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 17037 11203 17095 11209
rect 17037 11200 17049 11203
rect 16724 11172 17049 11200
rect 16724 11160 16730 11172
rect 17037 11169 17049 11172
rect 17083 11169 17095 11203
rect 17586 11200 17592 11212
rect 17499 11172 17592 11200
rect 17037 11163 17095 11169
rect 17586 11160 17592 11172
rect 17644 11160 17650 11212
rect 19058 11200 19064 11212
rect 19019 11172 19064 11200
rect 19058 11160 19064 11172
rect 19116 11160 19122 11212
rect 19426 11160 19432 11212
rect 19484 11200 19490 11212
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 19484 11172 19533 11200
rect 19484 11160 19490 11172
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 21082 11160 21088 11212
rect 21140 11200 21146 11212
rect 21304 11203 21362 11209
rect 21304 11200 21316 11203
rect 21140 11172 21316 11200
rect 21140 11160 21146 11172
rect 21304 11169 21316 11172
rect 21350 11169 21362 11203
rect 21304 11163 21362 11169
rect 23014 11160 23020 11212
rect 23072 11200 23078 11212
rect 23566 11200 23572 11212
rect 23072 11172 23572 11200
rect 23072 11160 23078 11172
rect 23566 11160 23572 11172
rect 23624 11200 23630 11212
rect 23880 11203 23938 11209
rect 23880 11200 23892 11203
rect 23624 11172 23892 11200
rect 23624 11160 23630 11172
rect 23880 11169 23892 11172
rect 23926 11169 23938 11203
rect 23880 11163 23938 11169
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 11793 11095 11851 11101
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 11808 11064 11836 11095
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11132 14703 11135
rect 15562 11132 15568 11144
rect 14691 11104 15568 11132
rect 14691 11101 14703 11104
rect 14645 11095 14703 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11101 22431 11135
rect 22373 11095 22431 11101
rect 11974 11064 11980 11076
rect 10192 11036 11980 11064
rect 10192 11024 10198 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22388 11064 22416 11095
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 22649 11135 22707 11141
rect 22649 11132 22661 11135
rect 22520 11104 22661 11132
rect 22520 11092 22526 11104
rect 22649 11101 22661 11104
rect 22695 11101 22707 11135
rect 22649 11095 22707 11101
rect 22336 11036 22416 11064
rect 22336 11024 22342 11036
rect 7745 10999 7803 11005
rect 7745 10996 7757 10999
rect 7616 10968 7757 10996
rect 7616 10956 7622 10968
rect 7745 10965 7757 10968
rect 7791 10965 7803 10999
rect 7745 10959 7803 10965
rect 9214 10956 9220 11008
rect 9272 10996 9278 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 9272 10968 9321 10996
rect 9272 10956 9278 10968
rect 9309 10965 9321 10968
rect 9355 10965 9367 10999
rect 12526 10996 12532 11008
rect 12487 10968 12532 10996
rect 9309 10959 9367 10965
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 16482 10956 16488 11008
rect 16540 10996 16546 11008
rect 17310 10996 17316 11008
rect 16540 10968 17316 10996
rect 16540 10956 16546 10968
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 19610 10956 19616 11008
rect 19668 10996 19674 11008
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 19668 10968 20085 10996
rect 19668 10956 19674 10968
rect 20073 10965 20085 10968
rect 20119 10965 20131 10999
rect 20073 10959 20131 10965
rect 22097 10999 22155 11005
rect 22097 10965 22109 10999
rect 22143 10996 22155 10999
rect 22186 10996 22192 11008
rect 22143 10968 22192 10996
rect 22143 10965 22155 10968
rect 22097 10959 22155 10965
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2406 10792 2412 10804
rect 2367 10764 2412 10792
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 2774 10792 2780 10804
rect 2735 10764 2780 10792
rect 2774 10752 2780 10764
rect 2832 10792 2838 10804
rect 4154 10792 4160 10804
rect 2832 10764 4160 10792
rect 2832 10752 2838 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 4396 10764 4445 10792
rect 4396 10752 4402 10764
rect 4433 10761 4445 10764
rect 4479 10761 4491 10795
rect 4433 10755 4491 10761
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9824 10764 9965 10792
rect 9824 10752 9830 10764
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10100 10764 10333 10792
rect 10100 10752 10106 10764
rect 10321 10761 10333 10764
rect 10367 10792 10379 10795
rect 10686 10792 10692 10804
rect 10367 10764 10692 10792
rect 10367 10761 10379 10764
rect 10321 10755 10379 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 13446 10792 13452 10804
rect 13407 10764 13452 10792
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 17083 10795 17141 10801
rect 17083 10792 17095 10795
rect 15620 10764 17095 10792
rect 15620 10752 15626 10764
rect 17083 10761 17095 10764
rect 17129 10761 17141 10795
rect 17083 10755 17141 10761
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 22002 10792 22008 10804
rect 21140 10764 22008 10792
rect 21140 10752 21146 10764
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22695 10795 22753 10801
rect 22695 10761 22707 10795
rect 22741 10792 22753 10795
rect 22830 10792 22836 10804
rect 22741 10764 22836 10792
rect 22741 10761 22753 10764
rect 22695 10755 22753 10761
rect 22830 10752 22836 10764
rect 22888 10752 22894 10804
rect 23382 10752 23388 10804
rect 23440 10792 23446 10804
rect 23799 10795 23857 10801
rect 23799 10792 23811 10795
rect 23440 10764 23811 10792
rect 23440 10752 23446 10764
rect 23799 10761 23811 10764
rect 23845 10761 23857 10795
rect 23799 10755 23857 10761
rect 2958 10684 2964 10736
rect 3016 10724 3022 10736
rect 4065 10727 4123 10733
rect 3016 10696 3096 10724
rect 3016 10684 3022 10696
rect 1486 10656 1492 10668
rect 1399 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10656 1550 10668
rect 1946 10656 1952 10668
rect 1544 10628 1952 10656
rect 1544 10616 1550 10628
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 3068 10665 3096 10696
rect 4065 10693 4077 10727
rect 4111 10724 4123 10727
rect 5534 10724 5540 10736
rect 4111 10696 5540 10724
rect 4111 10693 4123 10696
rect 4065 10687 4123 10693
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 6270 10724 6276 10736
rect 5920 10696 6276 10724
rect 5920 10665 5948 10696
rect 6270 10684 6276 10696
rect 6328 10684 6334 10736
rect 12710 10724 12716 10736
rect 8173 10696 12716 10724
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3053 10619 3111 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 7377 10659 7435 10665
rect 6236 10628 6868 10656
rect 6236 10616 6242 10628
rect 6840 10600 6868 10628
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 8173 10656 8201 10696
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 15654 10684 15660 10736
rect 15712 10724 15718 10736
rect 22370 10724 22376 10736
rect 15712 10696 22376 10724
rect 15712 10684 15718 10696
rect 22370 10684 22376 10696
rect 22428 10684 22434 10736
rect 7423 10628 8201 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10192 10628 10609 10656
rect 10192 10616 10198 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 10962 10656 10968 10668
rect 10923 10628 10968 10656
rect 10597 10619 10655 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 12802 10656 12808 10668
rect 12763 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 14921 10659 14979 10665
rect 14921 10656 14933 10659
rect 14200 10628 14933 10656
rect 5166 10588 5172 10600
rect 5127 10560 5172 10588
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 6822 10588 6828 10600
rect 5491 10560 6224 10588
rect 6735 10560 6828 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 1670 10520 1676 10532
rect 1627 10492 1676 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10489 2191 10523
rect 3142 10520 3148 10532
rect 3103 10492 3148 10520
rect 2133 10483 2191 10489
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 2148 10452 2176 10483
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 3697 10523 3755 10529
rect 3697 10520 3709 10523
rect 3574 10492 3709 10520
rect 3574 10452 3602 10492
rect 3697 10489 3709 10492
rect 3743 10489 3755 10523
rect 3697 10483 3755 10489
rect 4982 10452 4988 10464
rect 1820 10424 3602 10452
rect 4943 10424 4988 10452
rect 1820 10412 1826 10424
rect 4982 10412 4988 10424
rect 5040 10452 5046 10464
rect 5276 10452 5304 10551
rect 6196 10464 6224 10560
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 7466 10588 7472 10600
rect 7055 10560 7472 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 8036 10560 8217 10588
rect 6178 10452 6184 10464
rect 5040 10424 5304 10452
rect 6139 10424 6184 10452
rect 5040 10412 5046 10424
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 8036 10461 8064 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8205 10551 8263 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 9364 10560 9413 10588
rect 9364 10548 9370 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 14001 10591 14059 10597
rect 14001 10588 14013 10591
rect 13872 10560 14013 10588
rect 13872 10548 13878 10560
rect 14001 10557 14013 10560
rect 14047 10557 14059 10591
rect 14001 10551 14059 10557
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14200 10597 14228 10628
rect 14921 10625 14933 10628
rect 14967 10656 14979 10659
rect 15470 10656 15476 10668
rect 14967 10628 15476 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 15470 10616 15476 10628
rect 15528 10656 15534 10668
rect 18509 10659 18567 10665
rect 18509 10656 18521 10659
rect 15528 10628 18521 10656
rect 15528 10616 15534 10628
rect 18509 10625 18521 10628
rect 18555 10625 18567 10659
rect 18509 10619 18567 10625
rect 20165 10659 20223 10665
rect 20165 10625 20177 10659
rect 20211 10656 20223 10659
rect 23014 10656 23020 10668
rect 20211 10628 23020 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23566 10616 23572 10668
rect 23624 10656 23630 10668
rect 24489 10659 24547 10665
rect 24489 10656 24501 10659
rect 23624 10628 24501 10656
rect 23624 10616 23630 10628
rect 24489 10625 24501 10628
rect 24535 10625 24547 10659
rect 24489 10619 24547 10625
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 14148 10560 14197 10588
rect 14148 10548 14154 10560
rect 14185 10557 14197 10560
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14599 10560 15301 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 15289 10557 15301 10560
rect 15335 10588 15347 10591
rect 15562 10588 15568 10600
rect 15335 10560 15568 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 15930 10588 15936 10600
rect 15891 10560 15936 10588
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16850 10588 16856 10600
rect 16163 10560 16856 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 16980 10591 17038 10597
rect 16980 10557 16992 10591
rect 17026 10557 17038 10591
rect 16980 10551 17038 10557
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18230 10588 18236 10600
rect 17911 10560 18236 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 9674 10520 9680 10532
rect 9635 10492 9680 10520
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 12526 10520 12532 10532
rect 10744 10492 10789 10520
rect 12487 10492 12532 10520
rect 10744 10480 10750 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10520 12679 10523
rect 12986 10520 12992 10532
rect 12667 10492 12992 10520
rect 12667 10489 12679 10492
rect 12621 10483 12679 10489
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7616 10424 7665 10452
rect 7616 10412 7622 10424
rect 7653 10421 7665 10424
rect 7699 10452 7711 10455
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7699 10424 8033 10452
rect 7699 10421 7711 10424
rect 7653 10415 7711 10421
rect 8021 10421 8033 10424
rect 8067 10421 8079 10455
rect 11606 10452 11612 10464
rect 11519 10424 11612 10452
rect 8021 10415 8079 10421
rect 11606 10412 11612 10424
rect 11664 10452 11670 10464
rect 12253 10455 12311 10461
rect 12253 10452 12265 10455
rect 11664 10424 12265 10452
rect 11664 10412 11670 10424
rect 12253 10421 12265 10424
rect 12299 10452 12311 10455
rect 12636 10452 12664 10483
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 16995 10520 17023 10551
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 22002 10548 22008 10600
rect 22060 10588 22066 10600
rect 22592 10591 22650 10597
rect 22592 10588 22604 10591
rect 22060 10560 22604 10588
rect 22060 10548 22066 10560
rect 22592 10557 22604 10560
rect 22638 10588 22650 10591
rect 23106 10588 23112 10600
rect 22638 10560 23112 10588
rect 22638 10557 22650 10560
rect 22592 10551 22650 10557
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 23728 10591 23786 10597
rect 23728 10557 23740 10591
rect 23774 10588 23786 10591
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23774 10560 23949 10588
rect 23774 10557 23786 10560
rect 23728 10551 23786 10557
rect 23937 10557 23949 10560
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 24118 10548 24124 10600
rect 24176 10588 24182 10600
rect 24708 10591 24766 10597
rect 24708 10588 24720 10591
rect 24176 10560 24720 10588
rect 24176 10548 24182 10560
rect 24708 10557 24720 10560
rect 24754 10588 24766 10591
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24754 10560 25145 10588
rect 24754 10557 24766 10560
rect 24708 10551 24766 10557
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 17405 10523 17463 10529
rect 17405 10520 17417 10523
rect 13786 10492 17417 10520
rect 12299 10424 12664 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13786 10452 13814 10492
rect 17405 10489 17417 10492
rect 17451 10489 17463 10523
rect 17405 10483 17463 10489
rect 18049 10523 18107 10529
rect 18049 10489 18061 10523
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 12768 10424 13814 10452
rect 12768 10412 12774 10424
rect 15930 10412 15936 10464
rect 15988 10452 15994 10464
rect 16482 10452 16488 10464
rect 15988 10424 16488 10452
rect 15988 10412 15994 10424
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16724 10424 16773 10452
rect 16724 10412 16730 10424
rect 16761 10421 16773 10424
rect 16807 10421 16819 10455
rect 16761 10415 16819 10421
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18064 10452 18092 10483
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 19058 10520 19064 10532
rect 18656 10492 19064 10520
rect 18656 10480 18662 10492
rect 19058 10480 19064 10492
rect 19116 10520 19122 10532
rect 19245 10523 19303 10529
rect 19245 10520 19257 10523
rect 19116 10492 19257 10520
rect 19116 10480 19122 10492
rect 19245 10489 19257 10492
rect 19291 10489 19303 10523
rect 19245 10483 19303 10489
rect 19334 10480 19340 10532
rect 19392 10520 19398 10532
rect 19521 10523 19579 10529
rect 19521 10520 19533 10523
rect 19392 10492 19533 10520
rect 19392 10480 19398 10492
rect 19521 10489 19533 10492
rect 19567 10489 19579 10523
rect 19521 10483 19579 10489
rect 19610 10480 19616 10532
rect 19668 10520 19674 10532
rect 21085 10523 21143 10529
rect 19668 10492 19713 10520
rect 19668 10480 19674 10492
rect 21085 10489 21097 10523
rect 21131 10489 21143 10523
rect 21085 10483 21143 10489
rect 18966 10452 18972 10464
rect 17920 10424 18972 10452
rect 17920 10412 17926 10424
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 20438 10452 20444 10464
rect 20399 10424 20444 10452
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 20901 10455 20959 10461
rect 20901 10421 20913 10455
rect 20947 10452 20959 10455
rect 21100 10452 21128 10483
rect 21174 10480 21180 10532
rect 21232 10520 21238 10532
rect 21726 10520 21732 10532
rect 21232 10492 21277 10520
rect 21687 10492 21732 10520
rect 21232 10480 21238 10492
rect 21726 10480 21732 10492
rect 21784 10480 21790 10532
rect 21818 10480 21824 10532
rect 21876 10520 21882 10532
rect 24811 10523 24869 10529
rect 24811 10520 24823 10523
rect 21876 10492 24823 10520
rect 21876 10480 21882 10492
rect 24811 10489 24823 10492
rect 24857 10489 24869 10523
rect 24811 10483 24869 10489
rect 21542 10452 21548 10464
rect 20947 10424 21548 10452
rect 20947 10421 20959 10424
rect 20901 10415 20959 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 23937 10455 23995 10461
rect 23937 10421 23949 10455
rect 23983 10452 23995 10455
rect 24210 10452 24216 10464
rect 23983 10424 24216 10452
rect 23983 10421 23995 10424
rect 23937 10415 23995 10421
rect 24210 10412 24216 10424
rect 24268 10412 24274 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2590 10248 2596 10260
rect 2503 10220 2596 10248
rect 2590 10208 2596 10220
rect 2648 10248 2654 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 2648 10220 3065 10248
rect 2648 10208 2654 10220
rect 3053 10217 3065 10220
rect 3099 10248 3111 10251
rect 3142 10248 3148 10260
rect 3099 10220 3148 10248
rect 3099 10217 3111 10220
rect 3053 10211 3111 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3878 10248 3884 10260
rect 3839 10220 3884 10248
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 4341 10251 4399 10257
rect 4341 10217 4353 10251
rect 4387 10248 4399 10251
rect 4522 10248 4528 10260
rect 4387 10220 4528 10248
rect 4387 10217 4399 10220
rect 4341 10211 4399 10217
rect 4522 10208 4528 10220
rect 4580 10208 4586 10260
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6052 10220 6776 10248
rect 6052 10208 6058 10220
rect 2035 10183 2093 10189
rect 2035 10149 2047 10183
rect 2081 10180 2093 10183
rect 2406 10180 2412 10192
rect 2081 10152 2412 10180
rect 2081 10149 2093 10152
rect 2035 10143 2093 10149
rect 2406 10140 2412 10152
rect 2464 10140 2470 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 6236 10152 6684 10180
rect 6236 10140 6242 10152
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4798 10112 4804 10124
rect 4759 10084 4804 10112
rect 4798 10072 4804 10084
rect 4856 10072 4862 10124
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6365 10115 6423 10121
rect 6365 10112 6377 10115
rect 6135 10084 6377 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6365 10081 6377 10084
rect 6411 10112 6423 10115
rect 6546 10112 6552 10124
rect 6411 10084 6552 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6656 10121 6684 10152
rect 6641 10115 6699 10121
rect 6641 10081 6653 10115
rect 6687 10081 6699 10115
rect 6748 10112 6776 10220
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7745 10251 7803 10257
rect 7745 10248 7757 10251
rect 6880 10220 7757 10248
rect 6880 10208 6886 10220
rect 7745 10217 7757 10220
rect 7791 10248 7803 10251
rect 8018 10248 8024 10260
rect 7791 10220 8024 10248
rect 7791 10217 7803 10220
rect 7745 10211 7803 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 8478 10208 8484 10260
rect 8536 10248 8542 10260
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 8536 10220 9413 10248
rect 8536 10208 8542 10220
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9401 10211 9459 10217
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9732 10220 9873 10248
rect 9732 10208 9738 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 9968 10220 10916 10248
rect 7101 10183 7159 10189
rect 7101 10149 7113 10183
rect 7147 10180 7159 10183
rect 9214 10180 9220 10192
rect 7147 10152 9220 10180
rect 7147 10149 7159 10152
rect 7101 10143 7159 10149
rect 9214 10140 9220 10152
rect 9272 10180 9278 10192
rect 9968 10180 9996 10220
rect 10778 10180 10784 10192
rect 9272 10152 9996 10180
rect 10739 10152 10784 10180
rect 9272 10140 9278 10152
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 10888 10180 10916 10220
rect 11514 10208 11520 10260
rect 11572 10248 11578 10260
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 11572 10220 11621 10248
rect 11572 10208 11578 10220
rect 11609 10217 11621 10220
rect 11655 10217 11667 10251
rect 11974 10248 11980 10260
rect 11935 10220 11980 10248
rect 11609 10211 11667 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 14458 10248 14464 10260
rect 12216 10220 14464 10248
rect 12216 10208 12222 10220
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15105 10251 15163 10257
rect 15105 10217 15117 10251
rect 15151 10248 15163 10251
rect 15654 10248 15660 10260
rect 15151 10220 15660 10248
rect 15151 10217 15163 10220
rect 15105 10211 15163 10217
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 16945 10251 17003 10257
rect 16945 10217 16957 10251
rect 16991 10248 17003 10251
rect 17586 10248 17592 10260
rect 16991 10220 17592 10248
rect 16991 10217 17003 10220
rect 16945 10211 17003 10217
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19613 10251 19671 10257
rect 19613 10248 19625 10251
rect 19576 10220 19625 10248
rect 19576 10208 19582 10220
rect 19613 10217 19625 10220
rect 19659 10217 19671 10251
rect 19613 10211 19671 10217
rect 21821 10251 21879 10257
rect 21821 10217 21833 10251
rect 21867 10248 21879 10251
rect 22646 10248 22652 10260
rect 21867 10220 22652 10248
rect 21867 10217 21879 10220
rect 21821 10211 21879 10217
rect 22646 10208 22652 10220
rect 22704 10248 22710 10260
rect 22704 10220 22876 10248
rect 22704 10208 22710 10220
rect 17126 10180 17132 10192
rect 10888 10152 13400 10180
rect 17087 10152 17132 10180
rect 13372 10124 13400 10152
rect 17126 10140 17132 10152
rect 17184 10140 17190 10192
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 19055 10183 19113 10189
rect 17276 10152 17321 10180
rect 17276 10140 17282 10152
rect 19055 10149 19067 10183
rect 19101 10180 19113 10183
rect 19242 10180 19248 10192
rect 19101 10152 19248 10180
rect 19101 10149 19113 10152
rect 19055 10143 19113 10149
rect 19242 10140 19248 10152
rect 19300 10140 19306 10192
rect 19426 10140 19432 10192
rect 19484 10180 19490 10192
rect 19889 10183 19947 10189
rect 19889 10180 19901 10183
rect 19484 10152 19901 10180
rect 19484 10140 19490 10152
rect 19889 10149 19901 10152
rect 19935 10149 19947 10183
rect 19889 10143 19947 10149
rect 20898 10140 20904 10192
rect 20956 10180 20962 10192
rect 22848 10189 22876 10220
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 24305 10251 24363 10257
rect 24305 10248 24317 10251
rect 22980 10220 24317 10248
rect 22980 10208 22986 10220
rect 24305 10217 24317 10220
rect 24351 10217 24363 10251
rect 24305 10211 24363 10217
rect 21222 10183 21280 10189
rect 21222 10180 21234 10183
rect 20956 10152 21234 10180
rect 20956 10140 20962 10152
rect 21222 10149 21234 10152
rect 21268 10149 21280 10183
rect 21222 10143 21280 10149
rect 22833 10183 22891 10189
rect 22833 10149 22845 10183
rect 22879 10149 22891 10183
rect 22833 10143 22891 10149
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 6748 10084 7389 10112
rect 6641 10075 6699 10081
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 8110 10112 8116 10124
rect 8071 10084 8116 10112
rect 7377 10075 7435 10081
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 2314 10044 2320 10056
rect 1719 10016 2320 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 2314 10004 2320 10016
rect 2372 10044 2378 10056
rect 2372 10016 3740 10044
rect 2372 10004 2378 10016
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 3418 9908 3424 9920
rect 2740 9880 3424 9908
rect 2740 9868 2746 9880
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 3712 9908 3740 10016
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 7392 10044 7420 10075
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 12158 10112 12164 10124
rect 12119 10084 12164 10112
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12710 10112 12716 10124
rect 12623 10084 12716 10112
rect 12710 10072 12716 10084
rect 12768 10112 12774 10124
rect 12768 10084 13032 10112
rect 12768 10072 12774 10084
rect 7834 10044 7840 10056
rect 4396 10016 6592 10044
rect 7392 10016 7840 10044
rect 4396 10004 4402 10016
rect 3970 9936 3976 9988
rect 4028 9976 4034 9988
rect 4982 9976 4988 9988
rect 4028 9948 4988 9976
rect 4028 9936 4034 9948
rect 4982 9936 4988 9948
rect 5040 9936 5046 9988
rect 5905 9979 5963 9985
rect 5905 9945 5917 9979
rect 5951 9976 5963 9979
rect 6362 9976 6368 9988
rect 5951 9948 6368 9976
rect 5951 9945 5963 9948
rect 5905 9939 5963 9945
rect 6362 9936 6368 9948
rect 6420 9976 6426 9988
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 6420 9948 6469 9976
rect 6420 9936 6426 9948
rect 6457 9945 6469 9948
rect 6503 9945 6515 9979
rect 6564 9976 6592 10016
rect 7834 10004 7840 10016
rect 7892 10044 7898 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7892 10016 8033 10044
rect 7892 10004 7898 10016
rect 8021 10013 8033 10016
rect 8067 10044 8079 10047
rect 8662 10044 8668 10056
rect 8067 10016 8668 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8662 10004 8668 10016
rect 8720 10044 8726 10056
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 8720 10016 9045 10044
rect 8720 10004 8726 10016
rect 9033 10013 9045 10016
rect 9079 10013 9091 10047
rect 10686 10044 10692 10056
rect 10647 10016 10692 10044
rect 9033 10007 9091 10013
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 10962 10044 10968 10056
rect 10875 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13004 10044 13032 10084
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13412 10084 13737 10112
rect 13412 10072 13418 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 14090 10112 14096 10124
rect 13955 10084 14096 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 15654 10112 15660 10124
rect 15615 10084 15660 10112
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 18138 10112 18144 10124
rect 18051 10084 18144 10112
rect 18138 10072 18144 10084
rect 18196 10112 18202 10124
rect 21818 10112 21824 10124
rect 18196 10084 21824 10112
rect 18196 10072 18202 10084
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 24213 10115 24271 10121
rect 24213 10112 24225 10115
rect 23446 10084 24225 10112
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13004 10016 14197 10044
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 16114 10044 16120 10056
rect 16075 10016 16120 10044
rect 14185 10007 14243 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19150 10044 19156 10056
rect 18739 10016 19156 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19150 10004 19156 10016
rect 19208 10044 19214 10056
rect 19208 10016 20392 10044
rect 19208 10004 19214 10016
rect 10980 9976 11008 10004
rect 6564 9948 11008 9976
rect 6457 9939 6515 9945
rect 12986 9936 12992 9988
rect 13044 9976 13050 9988
rect 13630 9976 13636 9988
rect 13044 9948 13636 9976
rect 13044 9936 13050 9948
rect 13630 9936 13636 9948
rect 13688 9976 13694 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 13688 9948 14565 9976
rect 13688 9936 13694 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 17678 9976 17684 9988
rect 17639 9948 17684 9976
rect 14553 9939 14611 9945
rect 17678 9936 17684 9948
rect 17736 9936 17742 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 20257 9979 20315 9985
rect 20257 9976 20269 9979
rect 19392 9948 20269 9976
rect 19392 9936 19398 9948
rect 20257 9945 20269 9948
rect 20303 9945 20315 9979
rect 20364 9976 20392 10016
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20772 10016 20913 10044
rect 20772 10004 20778 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 22738 10044 22744 10056
rect 22699 10016 22744 10044
rect 20901 10007 20959 10013
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 23014 10044 23020 10056
rect 22975 10016 23020 10044
rect 23014 10004 23020 10016
rect 23072 10004 23078 10056
rect 22922 9976 22928 9988
rect 20364 9948 22928 9976
rect 20257 9939 20315 9945
rect 22922 9936 22928 9948
rect 22980 9936 22986 9988
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 23446 9976 23474 10084
rect 24213 10081 24225 10084
rect 24259 10081 24271 10115
rect 24762 10112 24768 10124
rect 24723 10084 24768 10112
rect 24213 10075 24271 10081
rect 24762 10072 24768 10084
rect 24820 10072 24826 10124
rect 23348 9948 23474 9976
rect 23348 9936 23354 9948
rect 4522 9908 4528 9920
rect 3712 9880 4528 9908
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 5224 9880 6101 9908
rect 5224 9868 5230 9880
rect 6089 9877 6101 9880
rect 6135 9908 6147 9911
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 6135 9880 6193 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 6181 9877 6193 9880
rect 6227 9877 6239 9911
rect 6181 9871 6239 9877
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 10229 9911 10287 9917
rect 10229 9908 10241 9911
rect 9916 9880 10241 9908
rect 9916 9868 9922 9880
rect 10229 9877 10241 9880
rect 10275 9877 10287 9911
rect 10229 9871 10287 9877
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 16393 9911 16451 9917
rect 16393 9908 16405 9911
rect 16356 9880 16405 9908
rect 16356 9868 16362 9880
rect 16393 9877 16405 9880
rect 16439 9877 16451 9911
rect 22278 9908 22284 9920
rect 22239 9880 22284 9908
rect 16393 9871 16451 9877
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 23198 9868 23204 9920
rect 23256 9908 23262 9920
rect 24762 9908 24768 9920
rect 23256 9880 24768 9908
rect 23256 9868 23262 9880
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1670 9704 1676 9716
rect 1631 9676 1676 9704
rect 1670 9664 1676 9676
rect 1728 9664 1734 9716
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2958 9704 2964 9716
rect 2919 9676 2964 9704
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 4065 9707 4123 9713
rect 4065 9673 4077 9707
rect 4111 9704 4123 9707
rect 6178 9704 6184 9716
rect 4111 9676 6184 9704
rect 4111 9673 4123 9676
rect 4065 9667 4123 9673
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8168 9676 8953 9704
rect 8168 9664 8174 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 10778 9704 10784 9716
rect 10739 9676 10784 9704
rect 8941 9667 8999 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 11471 9707 11529 9713
rect 11471 9673 11483 9707
rect 11517 9704 11529 9707
rect 12986 9704 12992 9716
rect 11517 9676 12992 9704
rect 11517 9673 11529 9676
rect 11471 9667 11529 9673
rect 12986 9664 12992 9676
rect 13044 9664 13050 9716
rect 13081 9707 13139 9713
rect 13081 9673 13093 9707
rect 13127 9704 13139 9707
rect 13265 9707 13323 9713
rect 13265 9704 13277 9707
rect 13127 9676 13277 9704
rect 13127 9673 13139 9676
rect 13081 9667 13139 9673
rect 13265 9673 13277 9676
rect 13311 9704 13323 9707
rect 13446 9704 13452 9716
rect 13311 9676 13452 9704
rect 13311 9673 13323 9676
rect 13265 9667 13323 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 13633 9707 13691 9713
rect 13633 9673 13645 9707
rect 13679 9704 13691 9707
rect 13722 9704 13728 9716
rect 13679 9676 13728 9704
rect 13679 9673 13691 9676
rect 13633 9667 13691 9673
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 15105 9707 15163 9713
rect 15105 9673 15117 9707
rect 15151 9704 15163 9707
rect 15838 9704 15844 9716
rect 15151 9676 15844 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 7800 9608 10609 9636
rect 7800 9596 7806 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 10597 9599 10655 9605
rect 10686 9596 10692 9648
rect 10744 9636 10750 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 10744 9608 11253 9636
rect 10744 9596 10750 9608
rect 11241 9605 11253 9608
rect 11287 9636 11299 9639
rect 12802 9636 12808 9648
rect 11287 9608 12808 9636
rect 11287 9605 11299 9608
rect 11241 9599 11299 9605
rect 12802 9596 12808 9608
rect 12860 9596 12866 9648
rect 15120 9636 15148 9667
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 16022 9704 16028 9716
rect 15983 9676 16028 9704
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 19153 9707 19211 9713
rect 19153 9673 19165 9707
rect 19199 9704 19211 9707
rect 19242 9704 19248 9716
rect 19199 9676 19248 9704
rect 19199 9673 19211 9676
rect 19153 9667 19211 9673
rect 19242 9664 19248 9676
rect 19300 9704 19306 9716
rect 19429 9707 19487 9713
rect 19429 9704 19441 9707
rect 19300 9676 19441 9704
rect 19300 9664 19306 9676
rect 19429 9673 19441 9676
rect 19475 9673 19487 9707
rect 19429 9667 19487 9673
rect 21634 9664 21640 9716
rect 21692 9704 21698 9716
rect 22646 9704 22652 9716
rect 21692 9676 22508 9704
rect 22607 9676 22652 9704
rect 21692 9664 21698 9676
rect 13233 9608 15148 9636
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9568 5319 9571
rect 6362 9568 6368 9580
rect 5307 9540 6368 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6687 9540 7512 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2041 9503 2099 9509
rect 2041 9500 2053 9503
rect 2004 9472 2053 9500
rect 2004 9460 2010 9472
rect 2041 9469 2053 9472
rect 2087 9500 2099 9503
rect 2590 9500 2596 9512
rect 2087 9472 2596 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 2740 9472 3525 9500
rect 2740 9460 2746 9472
rect 3513 9469 3525 9472
rect 3559 9500 3571 9503
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 3559 9472 4261 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 4249 9469 4261 9472
rect 4295 9500 4307 9503
rect 5166 9500 5172 9512
rect 4295 9472 4844 9500
rect 5127 9472 5172 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 4430 9432 4436 9444
rect 1912 9404 4436 9432
rect 1912 9392 1918 9404
rect 4430 9392 4436 9404
rect 4488 9392 4494 9444
rect 4816 9432 4844 9472
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5445 9503 5503 9509
rect 5445 9469 5457 9503
rect 5491 9500 5503 9503
rect 6730 9500 6736 9512
rect 5491 9472 6736 9500
rect 5491 9469 5503 9472
rect 5445 9463 5503 9469
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4816 9404 5089 9432
rect 5077 9401 5089 9404
rect 5123 9432 5135 9435
rect 5460 9432 5488 9463
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7484 9509 7512 9540
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8352 9540 11427 9568
rect 8352 9528 8358 9540
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 7558 9500 7564 9512
rect 7515 9472 7564 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7834 9500 7840 9512
rect 7795 9472 7840 9500
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8018 9500 8024 9512
rect 7979 9472 8024 9500
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 8938 9500 8944 9512
rect 8619 9472 8944 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 5123 9404 5488 9432
rect 5905 9435 5963 9441
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 6086 9432 6092 9444
rect 5951 9404 6092 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 6086 9392 6092 9404
rect 6144 9392 6150 9444
rect 6178 9392 6184 9444
rect 6236 9432 6242 9444
rect 7101 9435 7159 9441
rect 7101 9432 7113 9435
rect 6236 9404 7113 9432
rect 6236 9392 6242 9404
rect 7101 9401 7113 9404
rect 7147 9432 7159 9435
rect 8588 9432 8616 9463
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 11399 9509 11427 9540
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 13233 9568 13261 9608
rect 11848 9540 13261 9568
rect 11848 9528 11854 9540
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13688 9540 13829 9568
rect 13688 9528 13694 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 11384 9503 11442 9509
rect 11384 9469 11396 9503
rect 11430 9500 11442 9503
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11430 9472 11897 9500
rect 11430 9469 11442 9472
rect 11384 9463 11442 9469
rect 11885 9469 11897 9472
rect 11931 9500 11943 9503
rect 12618 9500 12624 9512
rect 11931 9472 12624 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12764 9503 12822 9509
rect 12764 9469 12776 9503
rect 12810 9500 12822 9503
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 12810 9472 13093 9500
rect 12810 9469 12822 9472
rect 12764 9463 12822 9469
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 9858 9432 9864 9444
rect 7147 9404 8616 9432
rect 9819 9404 9864 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 9953 9435 10011 9441
rect 9953 9401 9965 9435
rect 9999 9401 10011 9435
rect 9953 9395 10011 9401
rect 10505 9435 10563 9441
rect 10505 9401 10517 9435
rect 10551 9432 10563 9435
rect 10686 9432 10692 9444
rect 10551 9404 10692 9432
rect 10551 9401 10563 9404
rect 10505 9395 10563 9401
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4522 9364 4528 9376
rect 4212 9336 4528 9364
rect 4212 9324 4218 9336
rect 4522 9324 4528 9336
rect 4580 9324 4586 9376
rect 4709 9367 4767 9373
rect 4709 9333 4721 9367
rect 4755 9364 4767 9367
rect 5442 9364 5448 9376
rect 4755 9336 5448 9364
rect 4755 9333 4767 9336
rect 4709 9327 4767 9333
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9364 9646 9376
rect 9968 9364 9996 9395
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 13906 9392 13912 9444
rect 13964 9432 13970 9444
rect 14461 9435 14519 9441
rect 13964 9404 14009 9432
rect 13964 9392 13970 9404
rect 14461 9401 14473 9435
rect 14507 9432 14519 9435
rect 14826 9432 14832 9444
rect 14507 9404 14832 9432
rect 14507 9401 14519 9404
rect 14461 9395 14519 9401
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 9640 9336 9996 9364
rect 10597 9367 10655 9373
rect 9640 9324 9646 9336
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 12158 9364 12164 9376
rect 10643 9336 12164 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 12158 9324 12164 9336
rect 12216 9324 12222 9376
rect 12851 9367 12909 9373
rect 12851 9333 12863 9367
rect 12897 9364 12909 9367
rect 13630 9364 13636 9376
rect 12897 9336 13636 9364
rect 12897 9333 12909 9336
rect 12851 9327 12909 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 15473 9367 15531 9373
rect 15473 9333 15485 9367
rect 15519 9364 15531 9367
rect 15654 9364 15660 9376
rect 15519 9336 15660 9364
rect 15519 9333 15531 9336
rect 15473 9327 15531 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 16040 9364 16068 9664
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 20438 9636 20444 9648
rect 17460 9608 20444 9636
rect 17460 9596 17466 9608
rect 20438 9596 20444 9608
rect 20496 9636 20502 9648
rect 21174 9636 21180 9648
rect 20496 9608 21180 9636
rect 20496 9596 20502 9608
rect 21174 9596 21180 9608
rect 21232 9636 21238 9648
rect 21361 9639 21419 9645
rect 21361 9636 21373 9639
rect 21232 9608 21373 9636
rect 21232 9596 21238 9608
rect 21361 9605 21373 9608
rect 21407 9636 21419 9639
rect 21818 9636 21824 9648
rect 21407 9608 21824 9636
rect 21407 9605 21419 9608
rect 21361 9599 21419 9605
rect 21818 9596 21824 9608
rect 21876 9596 21882 9648
rect 22480 9636 22508 9676
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 24762 9664 24768 9716
rect 24820 9704 24826 9716
rect 25041 9707 25099 9713
rect 25041 9704 25053 9707
rect 24820 9676 25053 9704
rect 24820 9664 24826 9676
rect 25041 9673 25053 9676
rect 25087 9673 25099 9707
rect 25774 9704 25780 9716
rect 25735 9676 25780 9704
rect 25041 9667 25099 9673
rect 25774 9664 25780 9676
rect 25832 9664 25838 9716
rect 22480 9608 23244 9636
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 17736 9540 18429 9568
rect 17736 9528 17742 9540
rect 18417 9537 18429 9540
rect 18463 9568 18475 9571
rect 19334 9568 19340 9580
rect 18463 9540 19340 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 21634 9528 21640 9580
rect 21692 9568 21698 9580
rect 21913 9571 21971 9577
rect 21913 9568 21925 9571
rect 21692 9540 21925 9568
rect 21692 9528 21698 9540
rect 21913 9537 21925 9540
rect 21959 9568 21971 9571
rect 22738 9568 22744 9580
rect 21959 9540 22744 9568
rect 21959 9537 21971 9540
rect 21913 9531 21971 9537
rect 22738 9528 22744 9540
rect 22796 9568 22802 9580
rect 23017 9571 23075 9577
rect 23017 9568 23029 9571
rect 22796 9540 23029 9568
rect 22796 9528 22802 9540
rect 23017 9537 23029 9540
rect 23063 9537 23075 9571
rect 23216 9568 23244 9608
rect 23385 9571 23443 9577
rect 23385 9568 23397 9571
rect 23216 9540 23397 9568
rect 23017 9531 23075 9537
rect 23385 9537 23397 9540
rect 23431 9568 23443 9571
rect 23431 9540 23704 9568
rect 23431 9537 23443 9540
rect 23385 9531 23443 9537
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9500 16175 9503
rect 16298 9500 16304 9512
rect 16163 9472 16304 9500
rect 16163 9469 16175 9472
rect 16117 9463 16175 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 17218 9500 17224 9512
rect 17092 9472 17224 9500
rect 17092 9460 17098 9472
rect 17218 9460 17224 9472
rect 17276 9500 17282 9512
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 17276 9472 17325 9500
rect 17276 9460 17282 9472
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 17313 9463 17371 9469
rect 19518 9460 19524 9512
rect 19576 9500 19582 9512
rect 23676 9509 23704 9540
rect 19613 9503 19671 9509
rect 19613 9500 19625 9503
rect 19576 9472 19625 9500
rect 19576 9460 19582 9472
rect 19613 9469 19625 9472
rect 19659 9469 19671 9503
rect 19613 9463 19671 9469
rect 23661 9503 23719 9509
rect 23661 9469 23673 9503
rect 23707 9469 23719 9503
rect 23661 9463 23719 9469
rect 24213 9503 24271 9509
rect 24213 9469 24225 9503
rect 24259 9500 24271 9503
rect 24673 9503 24731 9509
rect 24673 9500 24685 9503
rect 24259 9472 24685 9500
rect 24259 9469 24271 9472
rect 24213 9463 24271 9469
rect 24673 9469 24685 9472
rect 24719 9469 24731 9503
rect 24673 9463 24731 9469
rect 25292 9503 25350 9509
rect 25292 9469 25304 9503
rect 25338 9500 25350 9503
rect 25774 9500 25780 9512
rect 25338 9472 25780 9500
rect 25338 9469 25350 9472
rect 25292 9463 25350 9469
rect 18138 9432 18144 9444
rect 18099 9404 18144 9432
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18233 9435 18291 9441
rect 18233 9401 18245 9435
rect 18279 9401 18291 9435
rect 18233 9395 18291 9401
rect 16485 9367 16543 9373
rect 16485 9364 16497 9367
rect 16040 9336 16497 9364
rect 16485 9333 16497 9336
rect 16531 9333 16543 9367
rect 16485 9327 16543 9333
rect 17037 9367 17095 9373
rect 17037 9333 17049 9367
rect 17083 9364 17095 9367
rect 17402 9364 17408 9376
rect 17083 9336 17408 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 17402 9324 17408 9336
rect 17460 9324 17466 9376
rect 17865 9367 17923 9373
rect 17865 9333 17877 9367
rect 17911 9364 17923 9367
rect 18248 9364 18276 9395
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 19934 9435 19992 9441
rect 19934 9432 19946 9435
rect 19300 9404 19946 9432
rect 19300 9392 19306 9404
rect 19934 9401 19946 9404
rect 19980 9432 19992 9435
rect 20898 9432 20904 9444
rect 19980 9404 20904 9432
rect 19980 9401 19992 9404
rect 19934 9395 19992 9401
rect 20898 9392 20904 9404
rect 20956 9392 20962 9444
rect 21266 9392 21272 9444
rect 21324 9432 21330 9444
rect 21637 9435 21695 9441
rect 21637 9432 21649 9435
rect 21324 9404 21649 9432
rect 21324 9392 21330 9404
rect 21637 9401 21649 9404
rect 21683 9401 21695 9435
rect 21637 9395 21695 9401
rect 21729 9435 21787 9441
rect 21729 9401 21741 9435
rect 21775 9432 21787 9435
rect 21818 9432 21824 9444
rect 21775 9404 21824 9432
rect 21775 9401 21787 9404
rect 21729 9395 21787 9401
rect 21818 9392 21824 9404
rect 21876 9392 21882 9444
rect 23290 9392 23296 9444
rect 23348 9432 23354 9444
rect 24228 9432 24256 9463
rect 25774 9460 25780 9472
rect 25832 9460 25838 9512
rect 23348 9404 24256 9432
rect 23348 9392 23354 9404
rect 18782 9364 18788 9376
rect 17911 9336 18788 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 20530 9364 20536 9376
rect 20491 9336 20536 9364
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 21450 9324 21456 9376
rect 21508 9364 21514 9376
rect 23753 9367 23811 9373
rect 23753 9364 23765 9367
rect 21508 9336 23765 9364
rect 21508 9324 21514 9336
rect 23753 9333 23765 9336
rect 23799 9333 23811 9367
rect 23753 9327 23811 9333
rect 23934 9324 23940 9376
rect 23992 9364 23998 9376
rect 25363 9367 25421 9373
rect 25363 9364 25375 9367
rect 23992 9336 25375 9364
rect 23992 9324 23998 9336
rect 25363 9333 25375 9336
rect 25409 9333 25421 9367
rect 25363 9327 25421 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 1486 9160 1492 9172
rect 1443 9132 1492 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 1486 9120 1492 9132
rect 1544 9120 1550 9172
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2314 9160 2320 9172
rect 2275 9132 2320 9160
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 3510 9160 3516 9172
rect 3471 9132 3516 9160
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 5074 9160 5080 9172
rect 3804 9132 5080 9160
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 8993 2467 9027
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2409 8987 2467 8993
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2424 8956 2452 8987
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3804 8965 3832 9132
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 6362 9160 6368 9172
rect 5828 9132 6368 9160
rect 5166 9092 5172 9104
rect 3896 9064 5172 9092
rect 3145 8959 3203 8965
rect 2188 8928 2636 8956
rect 2188 8916 2194 8928
rect 198 8848 204 8900
rect 256 8888 262 8900
rect 2501 8891 2559 8897
rect 2501 8888 2513 8891
rect 256 8860 2513 8888
rect 256 8848 262 8860
rect 2501 8857 2513 8860
rect 2547 8857 2559 8891
rect 2608 8888 2636 8928
rect 3145 8925 3157 8959
rect 3191 8956 3203 8959
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3191 8928 3801 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 3896 8888 3924 9064
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5828 9101 5856 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 6604 9132 6745 9160
rect 6604 9120 6610 9132
rect 6733 9129 6745 9132
rect 6779 9129 6791 9163
rect 6733 9123 6791 9129
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 7282 9160 7288 9172
rect 7239 9132 7288 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12710 9160 12716 9172
rect 12575 9132 12716 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 5813 9095 5871 9101
rect 5813 9061 5825 9095
rect 5859 9061 5871 9095
rect 5813 9055 5871 9061
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 9582 9092 9588 9104
rect 9180 9064 9588 9092
rect 9180 9052 9186 9064
rect 9582 9052 9588 9064
rect 9640 9092 9646 9104
rect 9861 9095 9919 9101
rect 9861 9092 9873 9095
rect 9640 9064 9873 9092
rect 9640 9052 9646 9064
rect 9861 9061 9873 9064
rect 9907 9061 9919 9095
rect 9861 9055 9919 9061
rect 4132 9027 4190 9033
rect 4132 8993 4144 9027
rect 4178 9024 4190 9027
rect 4246 9024 4252 9036
rect 4178 8996 4252 9024
rect 4178 8993 4190 8996
rect 4132 8987 4190 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 4522 9024 4528 9036
rect 4483 8996 4528 9024
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 5534 9024 5540 9036
rect 5495 8996 5540 9024
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 7558 9024 7564 9036
rect 7519 8996 7564 9024
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 7834 9024 7840 9036
rect 7795 8996 7840 9024
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 8113 9027 8171 9033
rect 8113 9024 8125 9027
rect 8076 8996 8125 9024
rect 8076 8984 8082 8996
rect 8113 8993 8125 8996
rect 8159 8993 8171 9027
rect 8665 9027 8723 9033
rect 8665 9024 8677 9027
rect 8113 8987 8171 8993
rect 8220 8996 8677 9024
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 5552 8956 5580 8984
rect 4028 8928 5580 8956
rect 4028 8916 4034 8928
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 8220 8956 8248 8996
rect 8665 8993 8677 8996
rect 8711 9024 8723 9027
rect 9306 9024 9312 9036
rect 8711 8996 9312 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 11790 9024 11796 9036
rect 11747 8996 11796 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 11790 8984 11796 8996
rect 11848 8984 11854 9036
rect 11977 9027 12035 9033
rect 11977 8993 11989 9027
rect 12023 9024 12035 9027
rect 12544 9024 12572 9123
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13320 9132 13369 9160
rect 13320 9120 13326 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 13504 9132 14197 9160
rect 13504 9120 13510 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 14185 9123 14243 9129
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 17184 9132 17325 9160
rect 17184 9120 17190 9132
rect 17313 9129 17325 9132
rect 17359 9129 17371 9163
rect 18782 9160 18788 9172
rect 18743 9132 18788 9160
rect 17313 9123 17371 9129
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 19150 9160 19156 9172
rect 19111 9132 19156 9160
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 20588 9132 22692 9160
rect 20588 9120 20594 9132
rect 16022 9052 16028 9104
rect 16080 9092 16086 9104
rect 16438 9095 16496 9101
rect 16438 9092 16450 9095
rect 16080 9064 16450 9092
rect 16080 9052 16086 9064
rect 16438 9061 16450 9064
rect 16484 9061 16496 9095
rect 16438 9055 16496 9061
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 18186 9095 18244 9101
rect 18186 9092 18198 9095
rect 17828 9064 18198 9092
rect 17828 9052 17834 9064
rect 18186 9061 18198 9064
rect 18232 9061 18244 9095
rect 18800 9092 18828 9120
rect 22664 9104 22692 9132
rect 23290 9120 23296 9172
rect 23348 9160 23354 9172
rect 23661 9163 23719 9169
rect 23661 9160 23673 9163
rect 23348 9132 23673 9160
rect 23348 9120 23354 9132
rect 23661 9129 23673 9132
rect 23707 9129 23719 9163
rect 23661 9123 23719 9129
rect 21082 9092 21088 9104
rect 18800 9064 21088 9092
rect 18186 9055 18244 9061
rect 21082 9052 21088 9064
rect 21140 9052 21146 9104
rect 21266 9052 21272 9104
rect 21324 9092 21330 9104
rect 21913 9095 21971 9101
rect 21913 9092 21925 9095
rect 21324 9064 21925 9092
rect 21324 9052 21330 9064
rect 21913 9061 21925 9064
rect 21959 9061 21971 9095
rect 22646 9092 22652 9104
rect 22559 9064 22652 9092
rect 21913 9055 21971 9061
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 23201 9095 23259 9101
rect 23201 9061 23213 9095
rect 23247 9092 23259 9095
rect 23566 9092 23572 9104
rect 23247 9064 23572 9092
rect 23247 9061 23259 9064
rect 23201 9055 23259 9061
rect 23566 9052 23572 9064
rect 23624 9052 23630 9104
rect 13906 9024 13912 9036
rect 12023 8996 12572 9024
rect 13867 8996 13912 9024
rect 12023 8993 12035 8996
rect 11977 8987 12035 8993
rect 8754 8956 8760 8968
rect 7524 8928 8248 8956
rect 8715 8928 8760 8956
rect 7524 8916 7530 8928
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 10778 8956 10784 8968
rect 9815 8928 10784 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11992 8956 12020 8987
rect 13906 8984 13912 8996
rect 13964 9024 13970 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 13964 8996 14565 9024
rect 13964 8984 13970 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 16114 9024 16120 9036
rect 16075 8996 16120 9024
rect 14553 8987 14611 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 16908 8996 17877 9024
rect 16908 8984 16914 8996
rect 17865 8993 17877 8996
rect 17911 9024 17923 9027
rect 18506 9024 18512 9036
rect 17911 8996 18512 9024
rect 17911 8993 17923 8996
rect 17865 8987 17923 8993
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 19848 9027 19906 9033
rect 19848 8993 19860 9027
rect 19894 9024 19906 9027
rect 20070 9024 20076 9036
rect 19894 8996 20076 9024
rect 19894 8993 19906 8996
rect 19848 8987 19906 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 25041 9027 25099 9033
rect 25041 8993 25053 9027
rect 25087 9024 25099 9027
rect 25130 9024 25136 9036
rect 25087 8996 25136 9024
rect 25087 8993 25099 8996
rect 25041 8987 25099 8993
rect 25130 8984 25136 8996
rect 25188 8984 25194 9036
rect 11296 8928 12020 8956
rect 12161 8959 12219 8965
rect 11296 8916 11302 8928
rect 12161 8925 12173 8959
rect 12207 8956 12219 8959
rect 12802 8956 12808 8968
rect 12207 8928 12808 8956
rect 12207 8925 12219 8928
rect 12161 8919 12219 8925
rect 12802 8916 12808 8928
rect 12860 8956 12866 8968
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12860 8928 13001 8956
rect 12860 8916 12866 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 19935 8959 19993 8965
rect 19935 8925 19947 8959
rect 19981 8956 19993 8959
rect 20622 8956 20628 8968
rect 19981 8928 20628 8956
rect 19981 8925 19993 8928
rect 19935 8919 19993 8925
rect 20622 8916 20628 8928
rect 20680 8956 20686 8968
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20680 8928 21005 8956
rect 20680 8916 20686 8928
rect 20993 8925 21005 8928
rect 21039 8925 21051 8959
rect 21266 8956 21272 8968
rect 21227 8928 21272 8956
rect 20993 8919 21051 8925
rect 21266 8916 21272 8928
rect 21324 8956 21330 8968
rect 21726 8956 21732 8968
rect 21324 8928 21732 8956
rect 21324 8916 21330 8928
rect 21726 8916 21732 8928
rect 21784 8956 21790 8968
rect 22557 8959 22615 8965
rect 22557 8956 22569 8959
rect 21784 8928 22569 8956
rect 21784 8916 21790 8928
rect 22557 8925 22569 8928
rect 22603 8956 22615 8959
rect 22922 8956 22928 8968
rect 22603 8928 22928 8956
rect 22603 8925 22615 8928
rect 22557 8919 22615 8925
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 24029 8959 24087 8965
rect 24029 8956 24041 8959
rect 23446 8928 24041 8956
rect 2608 8860 3924 8888
rect 2501 8851 2559 8857
rect 2516 8820 2544 8851
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 9916 8860 10333 8888
rect 9916 8848 9922 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 10321 8851 10379 8857
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 19705 8891 19763 8897
rect 19705 8888 19717 8891
rect 19576 8860 19717 8888
rect 19576 8848 19582 8860
rect 19705 8857 19717 8860
rect 19751 8888 19763 8891
rect 21450 8888 21456 8900
rect 19751 8860 21456 8888
rect 19751 8857 19763 8860
rect 19705 8851 19763 8857
rect 21450 8848 21456 8860
rect 21508 8848 21514 8900
rect 21542 8848 21548 8900
rect 21600 8888 21606 8900
rect 23446 8888 23474 8928
rect 24029 8925 24041 8928
rect 24075 8925 24087 8959
rect 24029 8919 24087 8925
rect 21600 8860 23474 8888
rect 21600 8848 21606 8860
rect 2774 8820 2780 8832
rect 2516 8792 2780 8820
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4203 8823 4261 8829
rect 4203 8820 4215 8823
rect 3844 8792 4215 8820
rect 3844 8780 3850 8792
rect 4203 8789 4215 8792
rect 4249 8789 4261 8823
rect 4203 8783 4261 8789
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5994 8820 6000 8832
rect 5031 8792 6000 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17276 8792 17693 8820
rect 17276 8780 17282 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 17681 8783 17739 8789
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 20625 8823 20683 8829
rect 20625 8820 20637 8823
rect 19484 8792 20637 8820
rect 19484 8780 19490 8792
rect 20625 8789 20637 8792
rect 20671 8820 20683 8823
rect 20714 8820 20720 8832
rect 20671 8792 20720 8820
rect 20671 8789 20683 8792
rect 20625 8783 20683 8789
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 20990 8780 20996 8832
rect 21048 8820 21054 8832
rect 21266 8820 21272 8832
rect 21048 8792 21272 8820
rect 21048 8780 21054 8792
rect 21266 8780 21272 8792
rect 21324 8780 21330 8832
rect 24026 8780 24032 8832
rect 24084 8820 24090 8832
rect 25179 8823 25237 8829
rect 25179 8820 25191 8823
rect 24084 8792 25191 8820
rect 24084 8780 24090 8792
rect 25179 8789 25191 8792
rect 25225 8789 25237 8823
rect 25179 8783 25237 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2501 8619 2559 8625
rect 2501 8585 2513 8619
rect 2547 8616 2559 8619
rect 2682 8616 2688 8628
rect 2547 8588 2688 8616
rect 2547 8585 2559 8588
rect 2501 8579 2559 8585
rect 2682 8576 2688 8588
rect 2740 8576 2746 8628
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 3970 8616 3976 8628
rect 2832 8588 3976 8616
rect 2832 8576 2838 8588
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 5442 8616 5448 8628
rect 4126 8588 5448 8616
rect 106 8508 112 8560
rect 164 8548 170 8560
rect 3145 8551 3203 8557
rect 3145 8548 3157 8551
rect 164 8520 3157 8548
rect 164 8508 170 8520
rect 3145 8517 3157 8520
rect 3191 8517 3203 8551
rect 3145 8511 3203 8517
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 4126 8480 4154 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5592 8588 5825 8616
rect 5592 8576 5598 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 6052 8588 6653 8616
rect 6052 8576 6058 8588
rect 6641 8585 6653 8588
rect 6687 8616 6699 8619
rect 7834 8616 7840 8628
rect 6687 8588 7840 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8720 8588 9413 8616
rect 8720 8576 8726 8588
rect 9401 8585 9413 8588
rect 9447 8616 9459 8619
rect 9766 8616 9772 8628
rect 9447 8588 9772 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10778 8616 10784 8628
rect 10739 8588 10784 8616
rect 10778 8576 10784 8588
rect 10836 8616 10842 8628
rect 17770 8616 17776 8628
rect 10836 8588 11376 8616
rect 10836 8576 10842 8588
rect 5350 8548 5356 8560
rect 5000 8520 5356 8548
rect 5000 8480 5028 8520
rect 5350 8508 5356 8520
rect 5408 8548 5414 8560
rect 8110 8548 8116 8560
rect 5408 8520 8116 8548
rect 5408 8508 5414 8520
rect 8110 8508 8116 8520
rect 8168 8508 8174 8560
rect 11238 8548 11244 8560
rect 11199 8520 11244 8548
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 3651 8452 4154 8480
rect 4816 8452 5028 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8412 3019 8415
rect 3786 8412 3792 8424
rect 3007 8384 3792 8412
rect 3007 8381 3019 8384
rect 2961 8375 3019 8381
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8412 4399 8415
rect 4522 8412 4528 8424
rect 4387 8384 4528 8412
rect 4387 8381 4399 8384
rect 4341 8375 4399 8381
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4816 8421 4844 8452
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 7340 8452 7849 8480
rect 7340 8440 7346 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8754 8440 8760 8492
rect 8812 8480 8818 8492
rect 9398 8480 9404 8492
rect 8812 8452 9404 8480
rect 8812 8440 8818 8452
rect 9398 8440 9404 8452
rect 9456 8480 9462 8492
rect 11348 8489 11376 8588
rect 16040 8588 17776 8616
rect 16040 8560 16068 8588
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 21082 8616 21088 8628
rect 21043 8588 21088 8616
rect 21082 8576 21088 8588
rect 21140 8576 21146 8628
rect 22646 8616 22652 8628
rect 22607 8588 22652 8616
rect 22646 8576 22652 8588
rect 22704 8576 22710 8628
rect 22922 8616 22928 8628
rect 22883 8588 22928 8616
rect 22922 8576 22928 8588
rect 22980 8576 22986 8628
rect 25130 8616 25136 8628
rect 25091 8588 25136 8616
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 16022 8548 16028 8560
rect 13320 8520 16028 8548
rect 13320 8508 13326 8520
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 17494 8548 17500 8560
rect 17407 8520 17500 8548
rect 17494 8508 17500 8520
rect 17552 8548 17558 8560
rect 17552 8520 18644 8548
rect 17552 8508 17558 8520
rect 9585 8483 9643 8489
rect 9585 8480 9597 8483
rect 9456 8452 9597 8480
rect 9456 8440 9462 8452
rect 9585 8449 9597 8452
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 11333 8443 11391 8449
rect 12894 8440 12900 8452
rect 12952 8480 12958 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 12952 8452 14105 8480
rect 12952 8440 12958 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14826 8440 14832 8492
rect 14884 8480 14890 8492
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 14884 8452 15025 8480
rect 14884 8440 14890 8452
rect 15013 8449 15025 8452
rect 15059 8449 15071 8483
rect 15013 8443 15071 8449
rect 15654 8440 15660 8492
rect 15712 8480 15718 8492
rect 15749 8483 15807 8489
rect 15749 8480 15761 8483
rect 15712 8452 15761 8480
rect 15712 8440 15718 8452
rect 15749 8449 15761 8452
rect 15795 8480 15807 8483
rect 15795 8452 18368 8480
rect 15795 8449 15807 8452
rect 15749 8443 15807 8449
rect 4801 8415 4859 8421
rect 4801 8381 4813 8415
rect 4847 8381 4859 8415
rect 5074 8412 5080 8424
rect 5035 8384 5080 8412
rect 4801 8375 4859 8381
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4816 8344 4844 8375
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 5442 8412 5448 8424
rect 5355 8384 5448 8412
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 7377 8415 7435 8421
rect 7377 8381 7389 8415
rect 7423 8412 7435 8415
rect 7558 8412 7564 8424
rect 7423 8384 7564 8412
rect 7423 8381 7435 8384
rect 7377 8375 7435 8381
rect 7558 8372 7564 8384
rect 7616 8412 7622 8424
rect 9490 8412 9496 8424
rect 7616 8384 9496 8412
rect 7616 8372 7622 8384
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 11422 8412 11428 8424
rect 9600 8384 11428 8412
rect 4019 8316 4844 8344
rect 5460 8344 5488 8372
rect 7466 8344 7472 8356
rect 5460 8316 7472 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 8158 8347 8216 8353
rect 8158 8313 8170 8347
rect 8204 8344 8216 8347
rect 8662 8344 8668 8356
rect 8204 8316 8668 8344
rect 8204 8313 8216 8316
rect 8158 8307 8216 8313
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4212 8248 4257 8276
rect 4212 8236 4218 8248
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 7653 8279 7711 8285
rect 7653 8276 7665 8279
rect 7432 8248 7665 8276
rect 7432 8236 7438 8248
rect 7653 8245 7665 8248
rect 7699 8276 7711 8279
rect 8173 8276 8201 8307
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 9600 8344 9628 8384
rect 11422 8372 11428 8384
rect 11480 8372 11486 8424
rect 16500 8421 16528 8452
rect 18340 8424 18368 8452
rect 18616 8424 18644 8520
rect 20070 8508 20076 8560
rect 20128 8548 20134 8560
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 20128 8520 20729 8548
rect 20128 8508 20134 8520
rect 20717 8517 20729 8520
rect 20763 8548 20775 8551
rect 23014 8548 23020 8560
rect 20763 8520 23020 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 23014 8508 23020 8520
rect 23072 8508 23078 8560
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8480 19211 8483
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19199 8452 19717 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19705 8449 19717 8452
rect 19751 8480 19763 8483
rect 19978 8480 19984 8492
rect 19751 8452 19984 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8480 20407 8483
rect 20990 8480 20996 8492
rect 20395 8452 20996 8480
rect 20395 8449 20407 8452
rect 20349 8443 20407 8449
rect 20990 8440 20996 8452
rect 21048 8440 21054 8492
rect 21266 8440 21272 8492
rect 21324 8480 21330 8492
rect 21634 8480 21640 8492
rect 21324 8452 21369 8480
rect 21595 8452 21640 8480
rect 21324 8440 21330 8452
rect 21634 8440 21640 8452
rect 21692 8440 21698 8492
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8381 16543 8415
rect 16666 8412 16672 8424
rect 16627 8384 16672 8412
rect 16485 8375 16543 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 18322 8412 18328 8424
rect 18283 8384 18328 8412
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 18598 8412 18604 8424
rect 18559 8384 18604 8412
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 18785 8415 18843 8421
rect 18785 8381 18797 8415
rect 18831 8412 18843 8415
rect 19426 8412 19432 8424
rect 18831 8384 19432 8412
rect 18831 8381 18843 8384
rect 18785 8375 18843 8381
rect 19426 8372 19432 8384
rect 19484 8372 19490 8424
rect 8772 8316 9628 8344
rect 8772 8288 8800 8316
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 9906 8347 9964 8353
rect 9906 8344 9918 8347
rect 9824 8316 9918 8344
rect 9824 8304 9830 8316
rect 9906 8313 9918 8316
rect 9952 8344 9964 8347
rect 12158 8344 12164 8356
rect 9952 8316 12164 8344
rect 9952 8313 9964 8316
rect 9906 8307 9964 8313
rect 12158 8304 12164 8316
rect 12216 8344 12222 8356
rect 13262 8353 13268 8356
rect 12713 8347 12771 8353
rect 12713 8344 12725 8347
rect 12216 8316 12725 8344
rect 12216 8304 12222 8316
rect 12713 8313 12725 8316
rect 12759 8344 12771 8347
rect 13218 8347 13268 8353
rect 13218 8344 13230 8347
rect 12759 8316 13230 8344
rect 12759 8313 12771 8316
rect 12713 8307 12771 8313
rect 13218 8313 13230 8316
rect 13264 8313 13268 8347
rect 13218 8307 13268 8313
rect 13262 8304 13268 8307
rect 13320 8304 13326 8356
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 14734 8344 14740 8356
rect 13688 8316 14740 8344
rect 13688 8304 13694 8316
rect 14734 8304 14740 8316
rect 14792 8304 14798 8356
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8313 14887 8347
rect 14829 8307 14887 8313
rect 8754 8276 8760 8288
rect 7699 8248 8201 8276
rect 8667 8248 8760 8276
rect 7699 8245 7711 8248
rect 7653 8239 7711 8245
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 9122 8276 9128 8288
rect 9083 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 10505 8279 10563 8285
rect 10505 8276 10517 8279
rect 9640 8248 10517 8276
rect 9640 8236 9646 8248
rect 10505 8245 10517 8248
rect 10551 8245 10563 8279
rect 11790 8276 11796 8288
rect 11751 8248 11796 8276
rect 10505 8239 10563 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 13817 8279 13875 8285
rect 13817 8245 13829 8279
rect 13863 8276 13875 8279
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 13863 8248 14473 8276
rect 13863 8245 13875 8248
rect 13817 8239 13875 8245
rect 14461 8245 14473 8248
rect 14507 8276 14519 8279
rect 14844 8276 14872 8307
rect 17034 8304 17040 8356
rect 17092 8344 17098 8356
rect 19521 8347 19579 8353
rect 19521 8344 19533 8347
rect 17092 8316 19533 8344
rect 17092 8304 17098 8316
rect 19521 8313 19533 8316
rect 19567 8344 19579 8347
rect 19797 8347 19855 8353
rect 19797 8344 19809 8347
rect 19567 8316 19809 8344
rect 19567 8313 19579 8316
rect 19521 8307 19579 8313
rect 19797 8313 19809 8316
rect 19843 8344 19855 8347
rect 21361 8347 21419 8353
rect 21361 8344 21373 8347
rect 19843 8316 21373 8344
rect 19843 8313 19855 8316
rect 19797 8307 19855 8313
rect 21361 8313 21373 8316
rect 21407 8313 21419 8347
rect 21361 8307 21419 8313
rect 15470 8276 15476 8288
rect 14507 8248 15476 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 21376 8276 21404 8307
rect 22189 8279 22247 8285
rect 22189 8276 22201 8279
rect 21376 8248 22201 8276
rect 22189 8245 22201 8248
rect 22235 8245 22247 8279
rect 22189 8239 22247 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1535 8075 1593 8081
rect 1535 8072 1547 8075
rect 1452 8044 1547 8072
rect 1452 8032 1458 8044
rect 1535 8041 1547 8044
rect 1581 8041 1593 8075
rect 1535 8035 1593 8041
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4246 8072 4252 8084
rect 3559 8044 4252 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4341 8075 4399 8081
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 4522 8072 4528 8084
rect 4387 8044 4528 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 8018 8072 8024 8084
rect 7883 8044 8024 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 9398 8072 9404 8084
rect 9359 8044 9404 8072
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 12802 8072 12808 8084
rect 9548 8044 11554 8072
rect 12763 8044 12808 8072
rect 9548 8032 9554 8044
rect 2498 7964 2504 8016
rect 2556 8004 2562 8016
rect 2593 8007 2651 8013
rect 2593 8004 2605 8007
rect 2556 7976 2605 8004
rect 2556 7964 2562 7976
rect 2593 7973 2605 7976
rect 2639 7973 2651 8007
rect 2593 7967 2651 7973
rect 1464 7939 1522 7945
rect 1464 7905 1476 7939
rect 1510 7936 1522 7939
rect 1762 7936 1768 7948
rect 1510 7908 1768 7936
rect 1510 7905 1522 7908
rect 1464 7899 1522 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 4540 7936 4568 8032
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 6270 8004 6276 8016
rect 5132 7976 6276 8004
rect 5132 7964 5138 7976
rect 4617 7939 4675 7945
rect 4617 7936 4629 7939
rect 4540 7908 4629 7936
rect 4617 7905 4629 7908
rect 4663 7905 4675 7939
rect 5350 7936 5356 7948
rect 5311 7908 5356 7936
rect 4617 7899 4675 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5644 7945 5672 7976
rect 6270 7964 6276 7976
rect 6328 7964 6334 8016
rect 8202 8004 8208 8016
rect 8115 7976 8208 8004
rect 8202 7964 8208 7976
rect 8260 8004 8266 8016
rect 8754 8004 8760 8016
rect 8260 7976 8760 8004
rect 8260 7964 8266 7976
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 9861 8007 9919 8013
rect 9861 7973 9873 8007
rect 9907 8004 9919 8007
rect 10134 8004 10140 8016
rect 9907 7976 10140 8004
rect 9907 7973 9919 7976
rect 9861 7967 9919 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 11422 8004 11428 8016
rect 11383 7976 11428 8004
rect 11422 7964 11428 7976
rect 11480 7964 11486 8016
rect 11526 8004 11554 8044
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14792 8044 14841 8072
rect 14792 8032 14798 8044
rect 14829 8041 14841 8044
rect 14875 8041 14887 8075
rect 14829 8035 14887 8041
rect 16114 8032 16120 8084
rect 16172 8072 16178 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16172 8044 16957 8072
rect 16172 8032 16178 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 18138 8072 18144 8084
rect 16945 8035 17003 8041
rect 17052 8044 18144 8072
rect 12894 8004 12900 8016
rect 11526 7976 12900 8004
rect 12894 7964 12900 7976
rect 12952 8004 12958 8016
rect 17052 8004 17080 8044
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18233 8075 18291 8081
rect 18233 8041 18245 8075
rect 18279 8072 18291 8075
rect 18322 8072 18328 8084
rect 18279 8044 18328 8072
rect 18279 8041 18291 8044
rect 18233 8035 18291 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 20622 8072 20628 8084
rect 20583 8044 20628 8072
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 12952 7976 17080 8004
rect 17313 8007 17371 8013
rect 12952 7964 12958 7976
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7905 5687 7939
rect 5629 7899 5687 7905
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7936 6055 7939
rect 6178 7936 6184 7948
rect 6043 7908 6184 7936
rect 6043 7905 6055 7908
rect 5997 7899 6055 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6952 7939 7010 7945
rect 6952 7936 6964 7939
rect 6696 7908 6964 7936
rect 6696 7896 6702 7908
rect 6952 7905 6964 7908
rect 6998 7905 7010 7939
rect 6952 7899 7010 7905
rect 12250 7896 12256 7948
rect 12308 7936 12314 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12308 7908 13001 7936
rect 12308 7896 12314 7908
rect 12989 7905 13001 7908
rect 13035 7936 13047 7939
rect 13170 7936 13176 7948
rect 13035 7908 13176 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13280 7945 13308 7976
rect 17313 7973 17325 8007
rect 17359 8004 17371 8007
rect 17402 8004 17408 8016
rect 17359 7976 17408 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17402 7964 17408 7976
rect 17460 7964 17466 8016
rect 18874 8004 18880 8016
rect 18835 7976 18880 8004
rect 18874 7964 18880 7976
rect 18932 7964 18938 8016
rect 21082 8004 21088 8016
rect 21043 7976 21088 8004
rect 21082 7964 21088 7976
rect 21140 7964 21146 8016
rect 21634 8004 21640 8016
rect 21595 7976 21640 8004
rect 21634 7964 21640 7976
rect 21692 7964 21698 8016
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 15930 7936 15936 7948
rect 15887 7908 15936 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 16117 7939 16175 7945
rect 16117 7905 16129 7939
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 22532 7939 22590 7945
rect 22532 7905 22544 7939
rect 22578 7936 22590 7939
rect 23014 7936 23020 7948
rect 22578 7908 23020 7936
rect 22578 7905 22590 7908
rect 22532 7899 22590 7905
rect 2498 7868 2504 7880
rect 2459 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2590 7828 2596 7880
rect 2648 7868 2654 7880
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2648 7840 3157 7868
rect 2648 7828 2654 7840
rect 3145 7837 3157 7840
rect 3191 7868 3203 7871
rect 4430 7868 4436 7880
rect 3191 7840 4436 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5040 7840 6101 7868
rect 5040 7828 5046 7840
rect 6089 7837 6101 7840
rect 6135 7868 6147 7871
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 6135 7840 6377 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 6365 7831 6423 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 8938 7868 8944 7880
rect 8803 7840 8944 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 8938 7828 8944 7840
rect 8996 7868 9002 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 8996 7840 9781 7868
rect 8996 7828 9002 7840
rect 9769 7837 9781 7840
rect 9815 7868 9827 7871
rect 9858 7868 9864 7880
rect 9815 7840 9864 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 9858 7828 9864 7840
rect 9916 7828 9922 7880
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 10836 7840 11345 7868
rect 10836 7828 10842 7840
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7868 13783 7871
rect 13771 7840 15976 7868
rect 13771 7837 13783 7840
rect 13725 7831 13783 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1670 7800 1676 7812
rect 992 7772 1676 7800
rect 992 7760 998 7772
rect 1670 7760 1676 7772
rect 1728 7800 1734 7812
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 1728 7772 1869 7800
rect 1728 7760 1734 7772
rect 1857 7769 1869 7772
rect 1903 7769 1915 7803
rect 1857 7763 1915 7769
rect 3881 7803 3939 7809
rect 3881 7769 3893 7803
rect 3927 7800 3939 7803
rect 4706 7800 4712 7812
rect 3927 7772 4712 7800
rect 3927 7769 3939 7772
rect 3881 7763 3939 7769
rect 4706 7760 4712 7772
rect 4764 7800 4770 7812
rect 5074 7800 5080 7812
rect 4764 7772 5080 7800
rect 4764 7760 4770 7772
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 9490 7760 9496 7812
rect 9548 7800 9554 7812
rect 10686 7800 10692 7812
rect 9548 7772 10692 7800
rect 9548 7760 9554 7772
rect 10686 7760 10692 7772
rect 10744 7800 10750 7812
rect 11624 7800 11652 7831
rect 10744 7772 11652 7800
rect 10744 7760 10750 7772
rect 12986 7760 12992 7812
rect 13044 7800 13050 7812
rect 13081 7803 13139 7809
rect 13081 7800 13093 7803
rect 13044 7772 13093 7800
rect 13044 7760 13050 7772
rect 13081 7769 13093 7772
rect 13127 7769 13139 7803
rect 15948 7800 15976 7840
rect 16132 7812 16160 7899
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 17218 7868 17224 7880
rect 17179 7840 17224 7868
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17678 7868 17684 7880
rect 17639 7840 17684 7868
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 18506 7828 18512 7880
rect 18564 7868 18570 7880
rect 18785 7871 18843 7877
rect 18785 7868 18797 7871
rect 18564 7840 18797 7868
rect 18564 7828 18570 7840
rect 18785 7837 18797 7840
rect 18831 7868 18843 7871
rect 20993 7871 21051 7877
rect 18831 7840 20024 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 16114 7800 16120 7812
rect 15948 7772 16120 7800
rect 13081 7763 13139 7769
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 19337 7803 19395 7809
rect 19337 7769 19349 7803
rect 19383 7769 19395 7803
rect 19996 7800 20024 7840
rect 20993 7837 21005 7871
rect 21039 7868 21051 7871
rect 21266 7868 21272 7880
rect 21039 7840 21272 7868
rect 21039 7837 21051 7840
rect 20993 7831 21051 7837
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 22603 7803 22661 7809
rect 22603 7800 22615 7803
rect 19996 7772 22615 7800
rect 19337 7763 19395 7769
rect 22603 7769 22615 7772
rect 22649 7769 22661 7803
rect 22603 7763 22661 7769
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 7055 7735 7113 7741
rect 7055 7732 7067 7735
rect 6972 7704 7067 7732
rect 6972 7692 6978 7704
rect 7055 7701 7067 7704
rect 7101 7701 7113 7735
rect 14550 7732 14556 7744
rect 14511 7704 14556 7732
rect 7055 7695 7113 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 15804 7704 16589 7732
rect 15804 7692 15810 7704
rect 16577 7701 16589 7704
rect 16623 7732 16635 7735
rect 16666 7732 16672 7744
rect 16623 7704 16672 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 19352 7732 19380 7763
rect 19886 7732 19892 7744
rect 19352 7704 19892 7732
rect 19886 7692 19892 7704
rect 19944 7692 19950 7744
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 21910 7732 21916 7744
rect 21600 7704 21916 7732
rect 21600 7692 21606 7704
rect 21910 7692 21916 7704
rect 21968 7692 21974 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2498 7528 2504 7540
rect 2179 7500 2504 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 4580 7500 6193 7528
rect 4580 7488 4586 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 6638 7528 6644 7540
rect 6599 7500 6644 7528
rect 6181 7491 6239 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 8021 7531 8079 7537
rect 8021 7497 8033 7531
rect 8067 7528 8079 7531
rect 8202 7528 8208 7540
rect 8067 7500 8208 7528
rect 8067 7497 8079 7500
rect 8021 7491 8079 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 8938 7528 8944 7540
rect 8899 7500 8944 7528
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 11241 7531 11299 7537
rect 11241 7497 11253 7531
rect 11287 7528 11299 7531
rect 11422 7528 11428 7540
rect 11287 7500 11428 7528
rect 11287 7497 11299 7500
rect 11241 7491 11299 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7528 12863 7531
rect 12894 7528 12900 7540
rect 12851 7500 12900 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 14001 7531 14059 7537
rect 14001 7528 14013 7531
rect 13004 7500 14013 7528
rect 1670 7420 1676 7472
rect 1728 7460 1734 7472
rect 8110 7460 8116 7472
rect 1728 7432 8116 7460
rect 1728 7420 1734 7432
rect 8110 7420 8116 7432
rect 8168 7460 8174 7472
rect 8389 7463 8447 7469
rect 8389 7460 8401 7463
rect 8168 7432 8401 7460
rect 8168 7420 8174 7432
rect 8389 7429 8401 7432
rect 8435 7429 8447 7463
rect 10042 7460 10048 7472
rect 10003 7432 10048 7460
rect 8389 7423 8447 7429
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3510 7392 3516 7404
rect 3283 7364 3516 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3510 7352 3516 7364
rect 3568 7392 3574 7404
rect 4154 7392 4160 7404
rect 3568 7364 4160 7392
rect 3568 7352 3574 7364
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 13004 7401 13032 7500
rect 14001 7497 14013 7500
rect 14047 7528 14059 7531
rect 14366 7528 14372 7540
rect 14047 7500 14372 7528
rect 14047 7497 14059 7500
rect 14001 7491 14059 7497
rect 14366 7488 14372 7500
rect 14424 7528 14430 7540
rect 14826 7528 14832 7540
rect 14424 7500 14832 7528
rect 14424 7488 14430 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15838 7488 15844 7540
rect 15896 7528 15902 7540
rect 16209 7531 16267 7537
rect 16209 7528 16221 7531
rect 15896 7500 16221 7528
rect 15896 7488 15902 7500
rect 16209 7497 16221 7500
rect 16255 7497 16267 7531
rect 17402 7528 17408 7540
rect 17363 7500 17408 7528
rect 16209 7491 16267 7497
rect 15657 7463 15715 7469
rect 15657 7429 15669 7463
rect 15703 7460 15715 7463
rect 15930 7460 15936 7472
rect 15703 7432 15936 7460
rect 15703 7429 15715 7432
rect 15657 7423 15715 7429
rect 15930 7420 15936 7432
rect 15988 7420 15994 7472
rect 7193 7395 7251 7401
rect 7193 7392 7205 7395
rect 6604 7364 7205 7392
rect 6604 7352 6610 7364
rect 7193 7361 7205 7364
rect 7239 7361 7251 7395
rect 7193 7355 7251 7361
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 13446 7392 13452 7404
rect 13407 7364 13452 7392
rect 12989 7355 13047 7361
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 14550 7392 14556 7404
rect 13648 7364 14556 7392
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1578 7324 1584 7336
rect 1443 7296 1584 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 6178 7324 6184 7336
rect 4755 7296 6184 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 11400 7327 11458 7333
rect 11400 7293 11412 7327
rect 11446 7324 11458 7327
rect 11882 7324 11888 7336
rect 11446 7296 11888 7324
rect 11446 7293 11458 7296
rect 11400 7287 11458 7293
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 2314 7216 2320 7268
rect 2372 7256 2378 7268
rect 3053 7259 3111 7265
rect 3053 7256 3065 7259
rect 2372 7228 3065 7256
rect 2372 7216 2378 7228
rect 3053 7225 3065 7228
rect 3099 7256 3111 7259
rect 3558 7259 3616 7265
rect 3558 7256 3570 7259
rect 3099 7228 3570 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 3558 7225 3570 7228
rect 3604 7256 3616 7259
rect 5347 7259 5405 7265
rect 5347 7256 5359 7259
rect 3604 7228 5359 7256
rect 3604 7225 3616 7228
rect 3558 7219 3616 7225
rect 5347 7225 5359 7228
rect 5393 7256 5405 7259
rect 5626 7256 5632 7268
rect 5393 7228 5632 7256
rect 5393 7225 5405 7228
rect 5347 7219 5405 7225
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 6914 7256 6920 7268
rect 6875 7228 6920 7256
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 7006 7216 7012 7268
rect 7064 7256 7070 7268
rect 9490 7256 9496 7268
rect 7064 7228 7109 7256
rect 9451 7228 9496 7256
rect 7064 7216 7070 7228
rect 9490 7216 9496 7228
rect 9548 7216 9554 7268
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 11609 7259 11667 7265
rect 9640 7228 9685 7256
rect 9640 7216 9646 7228
rect 11609 7225 11621 7259
rect 11655 7256 11667 7259
rect 11655 7228 13032 7256
rect 11655 7225 11667 7228
rect 11609 7219 11667 7225
rect 2406 7188 2412 7200
rect 2367 7160 2412 7188
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 4246 7188 4252 7200
rect 4203 7160 4252 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 5534 7148 5540 7200
rect 5592 7188 5598 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5592 7160 5917 7188
rect 5592 7148 5598 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 8720 7160 9321 7188
rect 8720 7148 8726 7160
rect 9309 7157 9321 7160
rect 9355 7188 9367 7191
rect 9600 7188 9628 7216
rect 9355 7160 9628 7188
rect 9355 7157 9367 7160
rect 9309 7151 9367 7157
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10192 7160 10425 7188
rect 10192 7148 10198 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 10413 7151 10471 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11882 7188 11888 7200
rect 11843 7160 11888 7188
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 13004 7188 13032 7228
rect 13078 7216 13084 7268
rect 13136 7256 13142 7268
rect 13136 7228 13181 7256
rect 13136 7216 13142 7228
rect 13648 7188 13676 7364
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13964 7296 14289 7324
rect 13964 7284 13970 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 16224 7324 16252 7491
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 21591 7531 21649 7537
rect 21591 7528 21603 7531
rect 20036 7500 21603 7528
rect 20036 7488 20042 7500
rect 21591 7497 21603 7500
rect 21637 7497 21649 7531
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 21591 7491 21649 7497
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 23382 7488 23388 7540
rect 23440 7528 23446 7540
rect 23799 7531 23857 7537
rect 23799 7528 23811 7531
rect 23440 7500 23811 7528
rect 23440 7488 23446 7500
rect 23799 7497 23811 7500
rect 23845 7497 23857 7531
rect 23799 7491 23857 7497
rect 20993 7463 21051 7469
rect 20993 7429 21005 7463
rect 21039 7460 21051 7463
rect 21082 7460 21088 7472
rect 21039 7432 21088 7460
rect 21039 7429 21051 7432
rect 20993 7423 21051 7429
rect 21082 7420 21088 7432
rect 21140 7420 21146 7472
rect 18138 7392 18144 7404
rect 18051 7364 18144 7392
rect 18138 7352 18144 7364
rect 18196 7392 18202 7404
rect 22603 7395 22661 7401
rect 22603 7392 22615 7395
rect 18196 7364 22615 7392
rect 18196 7352 18202 7364
rect 22603 7361 22615 7364
rect 22649 7361 22661 7395
rect 22603 7355 22661 7361
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 16224 7296 16405 7324
rect 14277 7287 14335 7293
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 14292 7256 14320 7287
rect 14645 7259 14703 7265
rect 14645 7256 14657 7259
rect 14292 7228 14657 7256
rect 14645 7225 14657 7228
rect 14691 7225 14703 7259
rect 14645 7219 14703 7225
rect 15197 7259 15255 7265
rect 15197 7225 15209 7259
rect 15243 7256 15255 7259
rect 15654 7256 15660 7268
rect 15243 7228 15660 7256
rect 15243 7225 15255 7228
rect 15197 7219 15255 7225
rect 15654 7216 15660 7228
rect 15712 7216 15718 7268
rect 16114 7216 16120 7268
rect 16172 7256 16178 7268
rect 16868 7256 16896 7287
rect 20714 7284 20720 7336
rect 20772 7324 20778 7336
rect 21488 7327 21546 7333
rect 21488 7324 21500 7327
rect 20772 7296 21500 7324
rect 20772 7284 20778 7296
rect 21488 7293 21500 7296
rect 21534 7324 21546 7327
rect 21913 7327 21971 7333
rect 21913 7324 21925 7327
rect 21534 7296 21925 7324
rect 21534 7293 21546 7296
rect 21488 7287 21546 7293
rect 21913 7293 21925 7296
rect 21959 7293 21971 7327
rect 21913 7287 21971 7293
rect 22516 7327 22574 7333
rect 22516 7293 22528 7327
rect 22562 7324 22574 7327
rect 22830 7324 22836 7336
rect 22562 7296 22836 7324
rect 22562 7293 22574 7296
rect 22516 7287 22574 7293
rect 22830 7284 22836 7296
rect 22888 7324 22894 7336
rect 23293 7327 23351 7333
rect 23293 7324 23305 7327
rect 22888 7296 23305 7324
rect 22888 7284 22894 7296
rect 23293 7293 23305 7296
rect 23339 7293 23351 7327
rect 23728 7327 23786 7333
rect 23728 7324 23740 7327
rect 23293 7287 23351 7293
rect 23446 7296 23740 7324
rect 17126 7256 17132 7268
rect 16172 7228 16896 7256
rect 17087 7228 17132 7256
rect 16172 7216 16178 7228
rect 17126 7216 17132 7228
rect 17184 7216 17190 7268
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7225 18291 7259
rect 18233 7219 18291 7225
rect 18785 7259 18843 7265
rect 18785 7225 18797 7259
rect 18831 7256 18843 7259
rect 19150 7256 19156 7268
rect 18831 7228 19156 7256
rect 18831 7225 18843 7228
rect 18785 7219 18843 7225
rect 17770 7188 17776 7200
rect 13004 7160 13676 7188
rect 17731 7160 17776 7188
rect 17770 7148 17776 7160
rect 17828 7188 17834 7200
rect 18248 7188 18276 7219
rect 19150 7216 19156 7228
rect 19208 7216 19214 7268
rect 19978 7256 19984 7268
rect 19939 7228 19984 7256
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 20070 7216 20076 7268
rect 20128 7256 20134 7268
rect 20625 7259 20683 7265
rect 20128 7228 20173 7256
rect 20128 7216 20134 7228
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 21726 7256 21732 7268
rect 20671 7228 21732 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 21726 7216 21732 7228
rect 21784 7256 21790 7268
rect 23446 7256 23474 7296
rect 23728 7293 23740 7296
rect 23774 7324 23786 7327
rect 24121 7327 24179 7333
rect 24121 7324 24133 7327
rect 23774 7296 24133 7324
rect 23774 7293 23786 7296
rect 23728 7287 23786 7293
rect 24121 7293 24133 7296
rect 24167 7293 24179 7327
rect 24121 7287 24179 7293
rect 21784 7228 23474 7256
rect 21784 7216 21790 7228
rect 18874 7188 18880 7200
rect 17828 7160 18880 7188
rect 17828 7148 17834 7160
rect 18874 7148 18880 7160
rect 18932 7188 18938 7200
rect 19061 7191 19119 7197
rect 19061 7188 19073 7191
rect 18932 7160 19073 7188
rect 18932 7148 18938 7160
rect 19061 7157 19073 7160
rect 19107 7157 19119 7191
rect 19061 7151 19119 7157
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 19705 7191 19763 7197
rect 19705 7188 19717 7191
rect 19576 7160 19717 7188
rect 19576 7148 19582 7160
rect 19705 7157 19717 7160
rect 19751 7157 19763 7191
rect 21266 7188 21272 7200
rect 21227 7160 21272 7188
rect 19705 7151 19763 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1762 6944 1768 6996
rect 1820 6984 1826 6996
rect 1857 6987 1915 6993
rect 1857 6984 1869 6987
rect 1820 6956 1869 6984
rect 1820 6944 1826 6956
rect 1857 6953 1869 6956
rect 1903 6953 1915 6987
rect 3510 6984 3516 6996
rect 3471 6956 3516 6984
rect 1857 6947 1915 6953
rect 3510 6944 3516 6956
rect 3568 6944 3574 6996
rect 3786 6984 3792 6996
rect 3747 6956 3792 6984
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5350 6984 5356 6996
rect 5215 6956 5356 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5537 6987 5595 6993
rect 5537 6953 5549 6987
rect 5583 6984 5595 6987
rect 5626 6984 5632 6996
rect 5583 6956 5632 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 5626 6944 5632 6956
rect 5684 6984 5690 6996
rect 5684 6956 6868 6984
rect 5684 6944 5690 6956
rect 2406 6916 2412 6928
rect 2367 6888 2412 6916
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 4246 6916 4252 6928
rect 3068 6888 4252 6916
rect 1578 6857 1584 6860
rect 1432 6851 1490 6857
rect 1432 6817 1444 6851
rect 1478 6817 1490 6851
rect 1432 6811 1490 6817
rect 1535 6851 1584 6857
rect 1535 6817 1547 6851
rect 1581 6817 1584 6851
rect 1535 6811 1584 6817
rect 1447 6780 1475 6811
rect 1578 6808 1584 6811
rect 1636 6848 1642 6860
rect 2225 6851 2283 6857
rect 2225 6848 2237 6851
rect 1636 6820 2237 6848
rect 1636 6808 1642 6820
rect 2225 6817 2237 6820
rect 2271 6817 2283 6851
rect 2225 6811 2283 6817
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3068 6857 3096 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 5994 6916 6000 6928
rect 5955 6888 6000 6916
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 6546 6916 6552 6928
rect 6507 6888 6552 6916
rect 6546 6876 6552 6888
rect 6604 6876 6610 6928
rect 6840 6916 6868 6956
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 6972 6956 7665 6984
rect 6972 6944 6978 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 7653 6947 7711 6953
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6984 11207 6987
rect 11238 6984 11244 6996
rect 11195 6956 11244 6984
rect 11195 6953 11207 6956
rect 11149 6947 11207 6953
rect 11238 6944 11244 6956
rect 11296 6984 11302 6996
rect 12986 6984 12992 6996
rect 11296 6956 11738 6984
rect 12947 6956 12992 6984
rect 11296 6944 11302 6956
rect 7374 6916 7380 6928
rect 6840 6888 7380 6916
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 10134 6916 10140 6928
rect 8803 6888 10140 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 11422 6916 11428 6928
rect 10336 6888 11428 6916
rect 10336 6860 10364 6888
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 3053 6851 3111 6857
rect 3053 6848 3065 6851
rect 3016 6820 3065 6848
rect 3016 6808 3022 6820
rect 3053 6817 3065 6820
rect 3099 6817 3111 6851
rect 8662 6848 8668 6860
rect 8623 6820 8668 6848
rect 3053 6811 3111 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9122 6808 9128 6860
rect 9180 6848 9186 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9180 6820 9689 6848
rect 9180 6808 9186 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 10318 6848 10324 6860
rect 10231 6820 10324 6848
rect 9677 6811 9735 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 11710 6857 11738 6956
rect 12986 6944 12992 6956
rect 13044 6944 13050 6996
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 13136 6956 13369 6984
rect 13136 6944 13142 6956
rect 13357 6953 13369 6956
rect 13403 6953 13415 6987
rect 13357 6947 13415 6953
rect 15703 6987 15761 6993
rect 15703 6953 15715 6987
rect 15749 6984 15761 6987
rect 17218 6984 17224 6996
rect 15749 6956 17224 6984
rect 15749 6953 15761 6956
rect 15703 6947 15761 6953
rect 17218 6944 17224 6956
rect 17276 6944 17282 6996
rect 18138 6984 18144 6996
rect 18099 6956 18144 6984
rect 18138 6944 18144 6956
rect 18196 6944 18202 6996
rect 18506 6984 18512 6996
rect 18467 6956 18512 6984
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 19518 6944 19524 6996
rect 19576 6984 19582 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 19576 6956 19901 6984
rect 19576 6944 19582 6956
rect 19889 6953 19901 6956
rect 19935 6984 19947 6987
rect 20070 6984 20076 6996
rect 19935 6956 20076 6984
rect 19935 6953 19947 6956
rect 19889 6947 19947 6953
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 13817 6919 13875 6925
rect 13817 6885 13829 6919
rect 13863 6916 13875 6919
rect 13906 6916 13912 6928
rect 13863 6888 13912 6916
rect 13863 6885 13875 6888
rect 13817 6879 13875 6885
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14366 6916 14372 6928
rect 14327 6888 14372 6916
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 16114 6916 16120 6928
rect 16075 6888 16120 6916
rect 16114 6876 16120 6888
rect 16172 6916 16178 6928
rect 16393 6919 16451 6925
rect 16393 6916 16405 6919
rect 16172 6888 16405 6916
rect 16172 6876 16178 6888
rect 16393 6885 16405 6888
rect 16439 6885 16451 6919
rect 16393 6879 16451 6885
rect 16666 6876 16672 6928
rect 16724 6916 16730 6928
rect 16898 6919 16956 6925
rect 16898 6916 16910 6919
rect 16724 6888 16910 6916
rect 16724 6876 16730 6888
rect 16898 6885 16910 6888
rect 16944 6885 16956 6919
rect 19242 6916 19248 6928
rect 19203 6888 19248 6916
rect 16898 6879 16956 6885
rect 19242 6876 19248 6888
rect 19300 6876 19306 6928
rect 21082 6916 21088 6928
rect 21043 6888 21088 6916
rect 21082 6876 21088 6888
rect 21140 6876 21146 6928
rect 21637 6919 21695 6925
rect 21637 6885 21649 6919
rect 21683 6916 21695 6919
rect 21726 6916 21732 6928
rect 21683 6888 21732 6916
rect 21683 6885 21695 6888
rect 21637 6879 21695 6885
rect 21726 6876 21732 6888
rect 21784 6876 21790 6928
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 11701 6851 11759 6857
rect 11701 6817 11713 6851
rect 11747 6817 11759 6851
rect 15562 6848 15568 6860
rect 15523 6820 15568 6848
rect 11701 6811 11759 6817
rect 2590 6780 2596 6792
rect 1447 6752 2596 6780
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4430 6780 4436 6792
rect 4391 6752 4436 6780
rect 4157 6743 4215 6749
rect 4172 6712 4200 6743
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 6638 6780 6644 6792
rect 5951 6752 6644 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 9582 6780 9588 6792
rect 7984 6752 9588 6780
rect 7984 6740 7990 6752
rect 9582 6740 9588 6752
rect 9640 6780 9646 6792
rect 11256 6780 11284 6811
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 16577 6851 16635 6857
rect 16577 6848 16589 6851
rect 16356 6820 16589 6848
rect 16356 6808 16362 6820
rect 16577 6817 16589 6820
rect 16623 6817 16635 6851
rect 16577 6811 16635 6817
rect 18598 6808 18604 6860
rect 18656 6848 18662 6860
rect 18656 6820 19104 6848
rect 18656 6808 18662 6820
rect 11606 6780 11612 6792
rect 9640 6752 11612 6780
rect 9640 6740 9646 6752
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 13725 6783 13783 6789
rect 13725 6749 13737 6783
rect 13771 6749 13783 6783
rect 13725 6743 13783 6749
rect 18969 6783 19027 6789
rect 18969 6749 18981 6783
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 4338 6712 4344 6724
rect 4172 6684 4344 6712
rect 4338 6672 4344 6684
rect 4396 6712 4402 6724
rect 6546 6712 6552 6724
rect 4396 6684 6552 6712
rect 4396 6672 4402 6684
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 13740 6712 13768 6743
rect 13688 6684 13768 6712
rect 13688 6672 13694 6684
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 5592 6616 6837 6644
rect 5592 6604 5598 6616
rect 6825 6613 6837 6616
rect 6871 6644 6883 6647
rect 7006 6644 7012 6656
rect 6871 6616 7012 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 16758 6604 16764 6656
rect 16816 6644 16822 6656
rect 17497 6647 17555 6653
rect 17497 6644 17509 6647
rect 16816 6616 17509 6644
rect 16816 6604 16822 6616
rect 17497 6613 17509 6616
rect 17543 6644 17555 6647
rect 17770 6644 17776 6656
rect 17543 6616 17776 6644
rect 17543 6613 17555 6616
rect 17497 6607 17555 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18782 6644 18788 6656
rect 18743 6616 18788 6644
rect 18782 6604 18788 6616
rect 18840 6644 18846 6656
rect 18984 6644 19012 6743
rect 19076 6712 19104 6820
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 20714 6780 20720 6792
rect 19208 6752 20720 6780
rect 19208 6740 19214 6752
rect 20714 6740 20720 6752
rect 20772 6780 20778 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20772 6752 21005 6780
rect 20772 6740 20778 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 21450 6712 21456 6724
rect 19076 6684 21456 6712
rect 21450 6672 21456 6684
rect 21508 6672 21514 6724
rect 18840 6616 19012 6644
rect 18840 6604 18846 6616
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1535 6443 1593 6449
rect 1535 6409 1547 6443
rect 1581 6440 1593 6443
rect 1670 6440 1676 6452
rect 1581 6412 1676 6440
rect 1581 6409 1593 6412
rect 1535 6403 1593 6409
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 1949 6443 2007 6449
rect 1949 6409 1961 6443
rect 1995 6440 2007 6443
rect 2222 6440 2228 6452
rect 1995 6412 2228 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 1464 6239 1522 6245
rect 1464 6205 1476 6239
rect 1510 6236 1522 6239
rect 1964 6236 1992 6403
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2590 6440 2596 6452
rect 2363 6412 2596 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 3559 6443 3617 6449
rect 3559 6440 3571 6443
rect 3476 6412 3571 6440
rect 3476 6400 3482 6412
rect 3559 6409 3571 6412
rect 3605 6409 3617 6443
rect 4246 6440 4252 6452
rect 4207 6412 4252 6440
rect 3559 6403 3617 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4706 6440 4712 6452
rect 4667 6412 4712 6440
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 7101 6443 7159 6449
rect 7101 6440 7113 6443
rect 6236 6412 7113 6440
rect 6236 6400 6242 6412
rect 7101 6409 7113 6412
rect 7147 6440 7159 6443
rect 7282 6440 7288 6452
rect 7147 6412 7288 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8662 6440 8668 6452
rect 8435 6412 8668 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 10318 6440 10324 6452
rect 10279 6412 10324 6440
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11664 6412 11805 6440
rect 11664 6400 11670 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 11793 6403 11851 6409
rect 7374 6372 7380 6384
rect 7287 6344 7380 6372
rect 7374 6332 7380 6344
rect 7432 6372 7438 6384
rect 7834 6372 7840 6384
rect 7432 6344 7840 6372
rect 7432 6332 7438 6344
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 10505 6375 10563 6381
rect 10505 6372 10517 6375
rect 9088 6344 10517 6372
rect 9088 6332 9094 6344
rect 10505 6341 10517 6344
rect 10551 6372 10563 6375
rect 10597 6375 10655 6381
rect 10597 6372 10609 6375
rect 10551 6344 10609 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 10597 6341 10609 6344
rect 10643 6341 10655 6375
rect 11808 6372 11836 6403
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13357 6443 13415 6449
rect 13357 6440 13369 6443
rect 13136 6412 13369 6440
rect 13136 6400 13142 6412
rect 13357 6409 13369 6412
rect 13403 6409 13415 6443
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13357 6403 13415 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 16114 6440 16120 6452
rect 15580 6412 16120 6440
rect 15580 6372 15608 6412
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 16298 6400 16304 6452
rect 16356 6440 16362 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16356 6412 17141 6440
rect 16356 6400 16362 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 17129 6403 17187 6409
rect 18966 6400 18972 6452
rect 19024 6440 19030 6452
rect 22830 6440 22836 6452
rect 19024 6412 22836 6440
rect 19024 6400 19030 6412
rect 22830 6400 22836 6412
rect 22888 6400 22894 6452
rect 11808 6344 15608 6372
rect 10597 6335 10655 6341
rect 15654 6332 15660 6384
rect 15712 6372 15718 6384
rect 16393 6375 16451 6381
rect 16393 6372 16405 6375
rect 15712 6344 16405 6372
rect 15712 6332 15718 6344
rect 16393 6341 16405 6344
rect 16439 6341 16451 6375
rect 16393 6335 16451 6341
rect 19061 6375 19119 6381
rect 19061 6341 19073 6375
rect 19107 6372 19119 6375
rect 19242 6372 19248 6384
rect 19107 6344 19248 6372
rect 19107 6341 19119 6344
rect 19061 6335 19119 6341
rect 19242 6332 19248 6344
rect 19300 6372 19306 6384
rect 19429 6375 19487 6381
rect 19429 6372 19441 6375
rect 19300 6344 19441 6372
rect 19300 6332 19306 6344
rect 19429 6341 19441 6344
rect 19475 6372 19487 6375
rect 19521 6375 19579 6381
rect 19521 6372 19533 6375
rect 19475 6344 19533 6372
rect 19475 6341 19487 6344
rect 19429 6335 19487 6341
rect 19521 6341 19533 6344
rect 19567 6341 19579 6375
rect 19521 6335 19579 6341
rect 20625 6375 20683 6381
rect 20625 6341 20637 6375
rect 20671 6372 20683 6375
rect 21082 6372 21088 6384
rect 20671 6344 21088 6372
rect 20671 6341 20683 6344
rect 20625 6335 20683 6341
rect 21082 6332 21088 6344
rect 21140 6372 21146 6384
rect 22465 6375 22523 6381
rect 22465 6372 22477 6375
rect 21140 6344 22477 6372
rect 21140 6332 21146 6344
rect 22465 6341 22477 6344
rect 22511 6341 22523 6375
rect 22465 6335 22523 6341
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2498 6304 2504 6316
rect 2455 6276 2504 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 5994 6304 6000 6316
rect 5951 6276 6000 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 5994 6264 6000 6276
rect 6052 6304 6058 6316
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 6052 6276 6193 6304
rect 6052 6264 6058 6276
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 6638 6304 6644 6316
rect 6551 6276 6644 6304
rect 6181 6267 6239 6273
rect 6638 6264 6644 6276
rect 6696 6304 6702 6316
rect 8938 6304 8944 6316
rect 6696 6276 8944 6304
rect 6696 6264 6702 6276
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9784 6276 11284 6304
rect 1510 6208 1992 6236
rect 3488 6239 3546 6245
rect 1510 6205 1522 6208
rect 1464 6199 1522 6205
rect 3488 6205 3500 6239
rect 3534 6236 3546 6239
rect 3970 6236 3976 6248
rect 3534 6208 3976 6236
rect 3534 6205 3546 6208
rect 3488 6199 3546 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6236 5135 6239
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5123 6208 5273 6236
rect 5123 6205 5135 6208
rect 5077 6199 5135 6205
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 5534 6236 5540 6248
rect 5307 6208 5540 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 7282 6236 7288 6248
rect 7243 6208 7288 6236
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6205 7619 6239
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 7561 6199 7619 6205
rect 9048 6208 9229 6236
rect 3970 6100 3976 6112
rect 3931 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7576 6100 7604 6199
rect 9048 6112 9076 6208
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 9784 6245 9812 6276
rect 11256 6248 11284 6276
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12434 6304 12440 6316
rect 12032 6276 12440 6304
rect 12032 6264 12038 6276
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 14366 6304 14372 6316
rect 14323 6276 14372 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14642 6304 14648 6316
rect 14603 6276 14648 6304
rect 14642 6264 14648 6276
rect 14700 6264 14706 6316
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6304 15899 6307
rect 16206 6304 16212 6316
rect 15887 6276 16212 6304
rect 15887 6273 15899 6276
rect 15841 6267 15899 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 18782 6304 18788 6316
rect 18743 6276 18788 6304
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 19306 6276 20913 6304
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9364 6208 9781 6236
rect 9364 6196 9370 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 10505 6239 10563 6245
rect 10505 6205 10517 6239
rect 10551 6236 10563 6239
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10551 6208 10793 6236
rect 10551 6205 10563 6208
rect 10505 6199 10563 6205
rect 10781 6205 10793 6208
rect 10827 6236 10839 6239
rect 10870 6236 10876 6248
rect 10827 6208 10876 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11238 6236 11244 6248
rect 11199 6208 11244 6236
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 12158 6196 12164 6248
rect 12216 6236 12222 6248
rect 18141 6239 18199 6245
rect 12216 6208 12802 6236
rect 12216 6196 12222 6208
rect 9953 6171 10011 6177
rect 9953 6137 9965 6171
rect 9999 6168 10011 6171
rect 11146 6168 11152 6180
rect 9999 6140 11152 6168
rect 9999 6137 10011 6140
rect 9953 6131 10011 6137
rect 11146 6128 11152 6140
rect 11204 6128 11210 6180
rect 11517 6171 11575 6177
rect 11517 6137 11529 6171
rect 11563 6168 11575 6171
rect 12618 6168 12624 6180
rect 11563 6140 12624 6168
rect 11563 6137 11575 6140
rect 11517 6131 11575 6137
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12774 6177 12802 6208
rect 18141 6205 18153 6239
rect 18187 6236 18199 6239
rect 18414 6236 18420 6248
rect 18187 6208 18420 6236
rect 18187 6205 18199 6208
rect 18141 6199 18199 6205
rect 12759 6171 12817 6177
rect 12759 6137 12771 6171
rect 12805 6137 12817 6171
rect 12759 6131 12817 6137
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14369 6171 14427 6177
rect 14369 6168 14381 6171
rect 14056 6140 14381 6168
rect 14056 6128 14062 6140
rect 14369 6137 14381 6140
rect 14415 6168 14427 6171
rect 15197 6171 15255 6177
rect 15197 6168 15209 6171
rect 14415 6140 15209 6168
rect 14415 6137 14427 6140
rect 14369 6131 14427 6137
rect 15197 6137 15209 6140
rect 15243 6168 15255 6171
rect 15933 6171 15991 6177
rect 15933 6168 15945 6171
rect 15243 6140 15945 6168
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 15933 6137 15945 6140
rect 15979 6137 15991 6171
rect 15933 6131 15991 6137
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 17773 6171 17831 6177
rect 17773 6168 17785 6171
rect 16172 6140 17785 6168
rect 16172 6128 16178 6140
rect 17773 6137 17785 6140
rect 17819 6168 17831 6171
rect 18156 6168 18184 6199
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18598 6236 18604 6248
rect 18559 6208 18604 6236
rect 18598 6196 18604 6208
rect 18656 6236 18662 6248
rect 19306 6236 19334 6276
rect 20901 6273 20913 6276
rect 20947 6304 20959 6307
rect 20947 6276 21956 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 18656 6208 19334 6236
rect 19705 6239 19763 6245
rect 18656 6196 18662 6208
rect 19705 6205 19717 6239
rect 19751 6236 19763 6239
rect 20162 6236 20168 6248
rect 19751 6208 20168 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 20162 6196 20168 6208
rect 20220 6236 20226 6248
rect 20220 6208 21404 6236
rect 20220 6196 20226 6208
rect 19426 6168 19432 6180
rect 17819 6140 18184 6168
rect 19339 6140 19432 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 19426 6128 19432 6140
rect 19484 6168 19490 6180
rect 20026 6171 20084 6177
rect 20026 6168 20038 6171
rect 19484 6140 20038 6168
rect 19484 6128 19490 6140
rect 20026 6137 20038 6140
rect 20072 6137 20084 6171
rect 20026 6131 20084 6137
rect 7742 6100 7748 6112
rect 7340 6072 7604 6100
rect 7703 6072 7748 6100
rect 7340 6060 7346 6072
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 9030 6100 9036 6112
rect 8991 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 13630 6100 13636 6112
rect 13591 6072 13636 6100
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 16761 6103 16819 6109
rect 16761 6100 16773 6103
rect 16724 6072 16773 6100
rect 16724 6060 16730 6072
rect 16761 6069 16773 6072
rect 16807 6100 16819 6103
rect 19061 6103 19119 6109
rect 19061 6100 19073 6103
rect 16807 6072 19073 6100
rect 16807 6069 16819 6072
rect 16761 6063 16819 6069
rect 19061 6069 19073 6072
rect 19107 6100 19119 6103
rect 19153 6103 19211 6109
rect 19153 6100 19165 6103
rect 19107 6072 19165 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 19153 6069 19165 6072
rect 19199 6069 19211 6103
rect 21376 6100 21404 6208
rect 21450 6196 21456 6248
rect 21508 6236 21514 6248
rect 21928 6245 21956 6276
rect 21913 6239 21971 6245
rect 21508 6208 21553 6236
rect 21508 6196 21514 6208
rect 21913 6205 21925 6239
rect 21959 6205 21971 6239
rect 21913 6199 21971 6205
rect 21545 6103 21603 6109
rect 21545 6100 21557 6103
rect 21376 6072 21557 6100
rect 19153 6063 19211 6069
rect 21545 6069 21557 6072
rect 21591 6069 21603 6103
rect 21545 6063 21603 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2547 5899 2605 5905
rect 2547 5865 2559 5899
rect 2593 5896 2605 5899
rect 3326 5896 3332 5908
rect 2593 5868 3332 5896
rect 2593 5865 2605 5868
rect 2547 5859 2605 5865
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 4338 5896 4344 5908
rect 4299 5868 4344 5896
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5353 5899 5411 5905
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 5442 5896 5448 5908
rect 5399 5868 5448 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 9306 5896 9312 5908
rect 9267 5868 9312 5896
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10091 5899 10149 5905
rect 10091 5865 10103 5899
rect 10137 5896 10149 5899
rect 10778 5896 10784 5908
rect 10137 5868 10784 5896
rect 10137 5865 10149 5868
rect 10091 5859 10149 5865
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11238 5896 11244 5908
rect 10919 5868 11244 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 12434 5896 12440 5908
rect 12395 5868 12440 5896
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 16022 5856 16028 5908
rect 16080 5896 16086 5908
rect 18141 5899 18199 5905
rect 18141 5896 18153 5899
rect 16080 5868 18153 5896
rect 16080 5856 16086 5868
rect 18141 5865 18153 5868
rect 18187 5896 18199 5899
rect 18598 5896 18604 5908
rect 18187 5868 18604 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18598 5856 18604 5868
rect 18656 5896 18662 5908
rect 19889 5899 19947 5905
rect 18656 5868 19288 5896
rect 18656 5856 18662 5868
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8570 5828 8576 5840
rect 7524 5800 8576 5828
rect 7524 5788 7530 5800
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 11511 5831 11569 5837
rect 11511 5797 11523 5831
rect 11557 5828 11569 5831
rect 12158 5828 12164 5840
rect 11557 5800 12164 5828
rect 11557 5797 11569 5800
rect 11511 5791 11569 5797
rect 12158 5788 12164 5800
rect 12216 5828 12222 5840
rect 13218 5831 13276 5837
rect 13218 5828 13230 5831
rect 12216 5800 13230 5828
rect 12216 5788 12222 5800
rect 13218 5797 13230 5800
rect 13264 5797 13276 5831
rect 15470 5828 15476 5840
rect 15431 5800 15476 5828
rect 13218 5791 13276 5797
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 17310 5828 17316 5840
rect 17271 5800 17316 5828
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 17865 5831 17923 5837
rect 17865 5797 17877 5831
rect 17911 5828 17923 5831
rect 19150 5828 19156 5840
rect 17911 5800 19156 5828
rect 17911 5797 17923 5800
rect 17865 5791 17923 5797
rect 19150 5788 19156 5800
rect 19208 5788 19214 5840
rect 19260 5772 19288 5868
rect 19889 5865 19901 5899
rect 19935 5896 19947 5899
rect 20162 5896 20168 5908
rect 19935 5868 20168 5896
rect 19935 5865 19947 5868
rect 19889 5859 19947 5865
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 21082 5828 21088 5840
rect 21043 5800 21088 5828
rect 21082 5788 21088 5800
rect 21140 5788 21146 5840
rect 21637 5831 21695 5837
rect 21637 5797 21649 5831
rect 21683 5828 21695 5831
rect 21726 5828 21732 5840
rect 21683 5800 21732 5828
rect 21683 5797 21695 5800
rect 21637 5791 21695 5797
rect 21726 5788 21732 5800
rect 21784 5788 21790 5840
rect 1464 5763 1522 5769
rect 1464 5729 1476 5763
rect 1510 5760 1522 5763
rect 2222 5760 2228 5772
rect 1510 5732 2228 5760
rect 1510 5729 1522 5732
rect 1464 5723 1522 5729
rect 2222 5720 2228 5732
rect 2280 5720 2286 5772
rect 2476 5763 2534 5769
rect 2476 5729 2488 5763
rect 2522 5760 2534 5763
rect 2866 5760 2872 5772
rect 2522 5732 2872 5760
rect 2522 5729 2534 5732
rect 2476 5723 2534 5729
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 4982 5720 4988 5772
rect 5040 5760 5046 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5040 5732 5549 5760
rect 5040 5720 5046 5732
rect 5537 5729 5549 5732
rect 5583 5760 5595 5763
rect 6178 5760 6184 5772
rect 5583 5732 6184 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 7834 5760 7840 5772
rect 7795 5732 7840 5760
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 10020 5763 10078 5769
rect 10020 5729 10032 5763
rect 10066 5760 10078 5763
rect 10134 5760 10140 5772
rect 10066 5732 10140 5760
rect 10066 5729 10078 5732
rect 10020 5723 10078 5729
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 11146 5760 11152 5772
rect 11107 5732 11152 5760
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12676 5732 12909 5760
rect 12676 5720 12682 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 18785 5763 18843 5769
rect 18785 5760 18797 5763
rect 12897 5723 12955 5729
rect 18248 5732 18797 5760
rect 18248 5704 18276 5732
rect 18785 5729 18797 5732
rect 18831 5760 18843 5763
rect 19058 5760 19064 5772
rect 18831 5732 19064 5760
rect 18831 5729 18843 5732
rect 18785 5723 18843 5729
rect 19058 5720 19064 5732
rect 19116 5720 19122 5772
rect 19242 5760 19248 5772
rect 19155 5732 19248 5760
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 15378 5692 15384 5704
rect 15339 5664 15384 5692
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 17218 5692 17224 5704
rect 17179 5664 17224 5692
rect 17218 5652 17224 5664
rect 17276 5652 17282 5704
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 19518 5692 19524 5704
rect 19479 5664 19524 5692
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 20993 5695 21051 5701
rect 20993 5661 21005 5695
rect 21039 5692 21051 5695
rect 21450 5692 21456 5704
rect 21039 5664 21456 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 1535 5627 1593 5633
rect 1535 5593 1547 5627
rect 1581 5624 1593 5627
rect 7374 5624 7380 5636
rect 1581 5596 7380 5624
rect 1581 5593 1593 5596
rect 1535 5587 1593 5593
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 12069 5627 12127 5633
rect 12069 5624 12081 5627
rect 11020 5596 12081 5624
rect 11020 5584 11026 5596
rect 12069 5593 12081 5596
rect 12115 5624 12127 5627
rect 13906 5624 13912 5636
rect 12115 5596 13912 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 13906 5584 13912 5596
rect 13964 5624 13970 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 13964 5596 14105 5624
rect 13964 5584 13970 5596
rect 14093 5593 14105 5596
rect 14139 5593 14151 5627
rect 14093 5587 14151 5593
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 8110 5556 8116 5568
rect 8071 5528 8116 5556
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14458 5556 14464 5568
rect 13872 5528 13917 5556
rect 14419 5528 14464 5556
rect 13872 5516 13878 5528
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 16206 5516 16212 5568
rect 16264 5556 16270 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 16264 5528 16313 5556
rect 16264 5516 16270 5528
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 20714 5556 20720 5568
rect 20675 5528 20720 5556
rect 16301 5519 16359 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1535 5355 1593 5361
rect 1535 5321 1547 5355
rect 1581 5352 1593 5355
rect 1854 5352 1860 5364
rect 1581 5324 1860 5352
rect 1581 5321 1593 5324
rect 1535 5315 1593 5321
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2685 5355 2743 5361
rect 2685 5321 2697 5355
rect 2731 5352 2743 5355
rect 2866 5352 2872 5364
rect 2731 5324 2872 5352
rect 2731 5321 2743 5324
rect 2685 5315 2743 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 8076 5324 9137 5352
rect 8076 5312 8082 5324
rect 9125 5321 9137 5324
rect 9171 5352 9183 5355
rect 9214 5352 9220 5364
rect 9171 5324 9220 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12158 5352 12164 5364
rect 11931 5324 12164 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 12713 5355 12771 5361
rect 12713 5352 12725 5355
rect 12676 5324 12725 5352
rect 12676 5312 12682 5324
rect 12713 5321 12725 5324
rect 12759 5321 12771 5355
rect 12713 5315 12771 5321
rect 13035 5355 13093 5361
rect 13035 5321 13047 5355
rect 13081 5352 13093 5355
rect 14458 5352 14464 5364
rect 13081 5324 14464 5352
rect 13081 5321 13093 5324
rect 13035 5315 13093 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15657 5355 15715 5361
rect 15657 5352 15669 5355
rect 15436 5324 15669 5352
rect 15436 5312 15442 5324
rect 15657 5321 15669 5324
rect 15703 5321 15715 5355
rect 19058 5352 19064 5364
rect 19019 5324 19064 5352
rect 15657 5315 15715 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19484 5324 19533 5352
rect 19484 5312 19490 5324
rect 19521 5321 19533 5324
rect 19567 5321 19579 5355
rect 19521 5315 19579 5321
rect 20625 5355 20683 5361
rect 20625 5321 20637 5355
rect 20671 5352 20683 5355
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20671 5324 21005 5352
rect 20671 5321 20683 5324
rect 20625 5315 20683 5321
rect 20993 5321 21005 5324
rect 21039 5352 21051 5355
rect 21082 5352 21088 5364
rect 21039 5324 21088 5352
rect 21039 5321 21051 5324
rect 20993 5315 21051 5321
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 7193 5287 7251 5293
rect 7193 5253 7205 5287
rect 7239 5284 7251 5287
rect 7561 5287 7619 5293
rect 7561 5284 7573 5287
rect 7239 5256 7573 5284
rect 7239 5253 7251 5256
rect 7193 5247 7251 5253
rect 7561 5253 7573 5256
rect 7607 5284 7619 5287
rect 7834 5284 7840 5296
rect 7607 5256 7840 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 7834 5244 7840 5256
rect 7892 5284 7898 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 7892 5256 8125 5284
rect 7892 5244 7898 5256
rect 8113 5253 8125 5256
rect 8159 5253 8171 5287
rect 11790 5284 11796 5296
rect 8113 5247 8171 5253
rect 9692 5256 11796 5284
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 7929 5219 7987 5225
rect 7929 5216 7941 5219
rect 7340 5188 7941 5216
rect 7340 5176 7346 5188
rect 7929 5185 7941 5188
rect 7975 5216 7987 5219
rect 8757 5219 8815 5225
rect 7975 5188 8340 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 8312 5160 8340 5188
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9692 5216 9720 5256
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 12176 5284 12204 5312
rect 13725 5287 13783 5293
rect 13725 5284 13737 5287
rect 12176 5256 13737 5284
rect 13725 5253 13737 5256
rect 13771 5253 13783 5287
rect 13725 5247 13783 5253
rect 8803 5188 9720 5216
rect 10045 5219 10103 5225
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10134 5216 10140 5228
rect 10091 5188 10140 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10134 5176 10140 5188
rect 10192 5216 10198 5228
rect 12526 5216 12532 5228
rect 10192 5188 12532 5216
rect 10192 5176 10198 5188
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 1464 5151 1522 5157
rect 1464 5117 1476 5151
rect 1510 5148 1522 5151
rect 1854 5148 1860 5160
rect 1510 5120 1860 5148
rect 1510 5117 1522 5120
rect 1464 5111 1522 5117
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 8018 5148 8024 5160
rect 7979 5120 8024 5148
rect 8018 5108 8024 5120
rect 8076 5108 8082 5160
rect 8294 5148 8300 5160
rect 8255 5120 8300 5148
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 12964 5151 13022 5157
rect 12964 5117 12976 5151
rect 13010 5148 13022 5151
rect 13354 5148 13360 5160
rect 13010 5120 13360 5148
rect 13010 5117 13022 5120
rect 12964 5111 13022 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 10870 5080 10876 5092
rect 1728 5052 10876 5080
rect 1728 5040 1734 5052
rect 10870 5040 10876 5052
rect 10928 5040 10934 5092
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 11517 5083 11575 5089
rect 11020 5052 11065 5080
rect 11020 5040 11026 5052
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 12802 5080 12808 5092
rect 11563 5052 12808 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 12802 5040 12808 5052
rect 12860 5040 12866 5092
rect 10689 5015 10747 5021
rect 10689 4981 10701 5015
rect 10735 5012 10747 5015
rect 10980 5012 11008 5040
rect 10735 4984 11008 5012
rect 13740 5012 13768 5247
rect 21450 5244 21456 5296
rect 21508 5284 21514 5296
rect 22465 5287 22523 5293
rect 22465 5284 22477 5287
rect 21508 5256 22477 5284
rect 21508 5244 21514 5256
rect 22465 5253 22477 5256
rect 22511 5253 22523 5287
rect 22465 5247 22523 5253
rect 13998 5216 14004 5228
rect 13911 5188 14004 5216
rect 13998 5176 14004 5188
rect 14056 5216 14062 5228
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14056 5188 14933 5216
rect 14056 5176 14062 5188
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5216 15439 5219
rect 15470 5216 15476 5228
rect 15427 5188 15476 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 14700 5120 14745 5148
rect 14700 5108 14706 5120
rect 14093 5083 14151 5089
rect 14093 5049 14105 5083
rect 14139 5080 14151 5083
rect 14182 5080 14188 5092
rect 14139 5052 14188 5080
rect 14139 5049 14151 5052
rect 14093 5043 14151 5049
rect 14182 5040 14188 5052
rect 14240 5080 14246 5092
rect 15396 5080 15424 5179
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 19705 5219 19763 5225
rect 19705 5216 19717 5219
rect 19576 5188 19717 5216
rect 19576 5176 19582 5188
rect 19705 5185 19717 5188
rect 19751 5185 19763 5219
rect 19705 5179 19763 5185
rect 20714 5176 20720 5228
rect 20772 5216 20778 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 20772 5188 21833 5216
rect 20772 5176 20778 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 16209 5151 16267 5157
rect 16209 5117 16221 5151
rect 16255 5148 16267 5151
rect 16298 5148 16304 5160
rect 16255 5120 16304 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 16530 5083 16588 5089
rect 16530 5080 16542 5083
rect 14240 5052 15424 5080
rect 16040 5052 16542 5080
rect 14240 5040 14246 5052
rect 16040 5021 16068 5052
rect 16530 5049 16542 5052
rect 16576 5080 16588 5083
rect 16666 5080 16672 5092
rect 16576 5052 16672 5080
rect 16576 5049 16588 5052
rect 16530 5043 16588 5049
rect 16666 5040 16672 5052
rect 16724 5040 16730 5092
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18138 5080 18144 5092
rect 17911 5052 18144 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 18233 5083 18291 5089
rect 18233 5049 18245 5083
rect 18279 5049 18291 5083
rect 18782 5080 18788 5092
rect 18743 5052 18788 5080
rect 18233 5043 18291 5049
rect 16025 5015 16083 5021
rect 16025 5012 16037 5015
rect 13740 4984 16037 5012
rect 10735 4981 10747 4984
rect 10689 4975 10747 4981
rect 16025 4981 16037 4984
rect 16071 4981 16083 5015
rect 16025 4975 16083 4981
rect 17129 5015 17187 5021
rect 17129 4981 17141 5015
rect 17175 5012 17187 5015
rect 17310 5012 17316 5024
rect 17175 4984 17316 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17310 4972 17316 4984
rect 17368 5012 17374 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 17368 4984 17417 5012
rect 17368 4972 17374 4984
rect 17405 4981 17417 4984
rect 17451 5012 17463 5015
rect 18248 5012 18276 5043
rect 18782 5040 18788 5052
rect 18840 5040 18846 5092
rect 19426 5040 19432 5092
rect 19484 5080 19490 5092
rect 20026 5083 20084 5089
rect 20026 5080 20038 5083
rect 19484 5052 20038 5080
rect 19484 5040 19490 5052
rect 20026 5049 20038 5052
rect 20072 5049 20084 5083
rect 21542 5080 21548 5092
rect 21503 5052 21548 5080
rect 20026 5043 20084 5049
rect 21542 5040 21548 5052
rect 21600 5040 21606 5092
rect 21637 5083 21695 5089
rect 21637 5049 21649 5083
rect 21683 5049 21695 5083
rect 21637 5043 21695 5049
rect 17451 4984 18276 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21361 5015 21419 5021
rect 21361 5012 21373 5015
rect 20956 4984 21373 5012
rect 20956 4972 20962 4984
rect 21361 4981 21373 4984
rect 21407 5012 21419 5015
rect 21652 5012 21680 5043
rect 21407 4984 21680 5012
rect 21407 4981 21419 4984
rect 21361 4975 21419 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1535 4811 1593 4817
rect 1535 4777 1547 4811
rect 1581 4808 1593 4811
rect 1670 4808 1676 4820
rect 1581 4780 1676 4808
rect 1581 4777 1593 4780
rect 1535 4771 1593 4777
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10137 4811 10195 4817
rect 10137 4808 10149 4811
rect 10008 4780 10149 4808
rect 10008 4768 10014 4780
rect 10137 4777 10149 4780
rect 10183 4808 10195 4811
rect 10686 4808 10692 4820
rect 10183 4780 10692 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 10870 4808 10876 4820
rect 10831 4780 10876 4808
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11146 4808 11152 4820
rect 11107 4780 11152 4808
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 13078 4808 13084 4820
rect 12299 4780 13084 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 13078 4768 13084 4780
rect 13136 4808 13142 4820
rect 14182 4808 14188 4820
rect 13136 4780 13308 4808
rect 14143 4780 14188 4808
rect 13136 4768 13142 4780
rect 11695 4743 11753 4749
rect 11695 4709 11707 4743
rect 11741 4740 11753 4743
rect 12158 4740 12164 4752
rect 11741 4712 12164 4740
rect 11741 4709 11753 4712
rect 11695 4703 11753 4709
rect 12158 4700 12164 4712
rect 12216 4700 12222 4752
rect 13280 4749 13308 4780
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 15565 4811 15623 4817
rect 15565 4808 15577 4811
rect 15436 4780 15577 4808
rect 15436 4768 15442 4780
rect 15565 4777 15577 4780
rect 15611 4777 15623 4811
rect 15565 4771 15623 4777
rect 15841 4811 15899 4817
rect 15841 4777 15853 4811
rect 15887 4808 15899 4811
rect 16022 4808 16028 4820
rect 15887 4780 16028 4808
rect 15887 4777 15899 4780
rect 15841 4771 15899 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 17276 4780 17785 4808
rect 17276 4768 17282 4780
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 19242 4808 19248 4820
rect 19203 4780 19248 4808
rect 17773 4771 17831 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 20165 4811 20223 4817
rect 20165 4808 20177 4811
rect 19576 4780 20177 4808
rect 19576 4768 19582 4780
rect 20165 4777 20177 4780
rect 20211 4777 20223 4811
rect 20165 4771 20223 4777
rect 13265 4743 13323 4749
rect 13265 4709 13277 4743
rect 13311 4709 13323 4743
rect 13265 4703 13323 4709
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 16758 4740 16764 4752
rect 16623 4712 16764 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 16758 4700 16764 4712
rect 16816 4700 16822 4752
rect 17862 4700 17868 4752
rect 17920 4740 17926 4752
rect 18319 4743 18377 4749
rect 18319 4740 18331 4743
rect 17920 4712 18331 4740
rect 17920 4700 17926 4712
rect 18319 4709 18331 4712
rect 18365 4740 18377 4743
rect 19426 4740 19432 4752
rect 18365 4712 19432 4740
rect 18365 4709 18377 4712
rect 18319 4703 18377 4709
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 20070 4740 20076 4752
rect 19755 4712 20076 4740
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9214 4672 9220 4684
rect 8904 4644 9220 4672
rect 8904 4632 8910 4644
rect 9214 4632 9220 4644
rect 9272 4672 9278 4684
rect 9674 4672 9680 4684
rect 9272 4644 9680 4672
rect 9272 4632 9278 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 9950 4672 9956 4684
rect 9911 4644 9956 4672
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 15378 4672 15384 4684
rect 15243 4644 15384 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 17218 4632 17224 4684
rect 17276 4672 17282 4684
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17276 4644 17969 4672
rect 17276 4632 17282 4644
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 19058 4632 19064 4684
rect 19116 4672 19122 4684
rect 19755 4681 19783 4712
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 19740 4675 19798 4681
rect 19740 4672 19752 4675
rect 19116 4644 19752 4672
rect 19116 4632 19122 4644
rect 19740 4641 19752 4644
rect 19786 4641 19798 4675
rect 19740 4635 19798 4641
rect 19843 4675 19901 4681
rect 19843 4641 19855 4675
rect 19889 4672 19901 4675
rect 21453 4675 21511 4681
rect 21453 4672 21465 4675
rect 19889 4644 21465 4672
rect 19889 4641 19901 4644
rect 19843 4635 19901 4641
rect 21453 4641 21465 4644
rect 21499 4672 21511 4675
rect 21542 4672 21548 4684
rect 21499 4644 21548 4672
rect 21499 4641 21511 4644
rect 21453 4635 21511 4641
rect 21542 4632 21548 4644
rect 21600 4632 21606 4684
rect 11330 4604 11336 4616
rect 11291 4576 11336 4604
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13446 4604 13452 4616
rect 13407 4576 13452 4604
rect 13173 4567 13231 4573
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 9766 4536 9772 4548
rect 7892 4508 9772 4536
rect 7892 4496 7898 4508
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 7926 4468 7932 4480
rect 7887 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 13188 4468 13216 4567
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16408 4576 16497 4604
rect 13464 4536 13492 4564
rect 16408 4548 16436 4576
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 17494 4604 17500 4616
rect 17175 4576 17500 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 13722 4536 13728 4548
rect 13464 4508 13728 4536
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 16390 4496 16396 4548
rect 16448 4496 16454 4548
rect 14642 4468 14648 4480
rect 12860 4440 14648 4468
rect 12860 4428 12866 4440
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 16298 4468 16304 4480
rect 16259 4440 16304 4468
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 17405 4471 17463 4477
rect 17405 4468 17417 4471
rect 17368 4440 17417 4468
rect 17368 4428 17374 4440
rect 17405 4437 17417 4440
rect 17451 4437 17463 4471
rect 18874 4468 18880 4480
rect 18835 4440 18880 4468
rect 17405 4431 17463 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 20990 4428 20996 4480
rect 21048 4468 21054 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 21048 4440 21097 4468
rect 21048 4428 21054 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 106 4224 112 4276
rect 164 4264 170 4276
rect 1394 4264 1400 4276
rect 164 4236 1400 4264
rect 164 4224 170 4236
rect 1394 4224 1400 4236
rect 1452 4264 1458 4276
rect 1581 4267 1639 4273
rect 1581 4264 1593 4267
rect 1452 4236 1593 4264
rect 1452 4224 1458 4236
rect 1581 4233 1593 4236
rect 1627 4233 1639 4267
rect 1581 4227 1639 4233
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 7248 4236 7573 4264
rect 7248 4224 7254 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 9950 4264 9956 4276
rect 7561 4227 7619 4233
rect 9324 4236 9956 4264
rect 7576 4060 7604 4227
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8478 4128 8484 4140
rect 7984 4100 8064 4128
rect 8439 4100 8484 4128
rect 7984 4088 7990 4100
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7576 4032 7757 4060
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7285 3927 7343 3933
rect 7285 3893 7297 3927
rect 7331 3924 7343 3927
rect 7558 3924 7564 3936
rect 7331 3896 7564 3924
rect 7331 3893 7343 3896
rect 7285 3887 7343 3893
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7760 3924 7788 4023
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 8036 4069 8064 4100
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9324 4069 9352 4236
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 12158 4264 12164 4276
rect 11931 4236 12164 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12802 4264 12808 4276
rect 12763 4236 12808 4264
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 13078 4264 13084 4276
rect 13039 4236 13084 4264
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 15378 4264 15384 4276
rect 15339 4236 15384 4264
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 16758 4264 16764 4276
rect 16719 4236 16764 4264
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 17126 4224 17132 4276
rect 17184 4264 17190 4276
rect 17405 4267 17463 4273
rect 17405 4264 17417 4267
rect 17184 4236 17417 4264
rect 17184 4224 17190 4236
rect 17405 4233 17417 4236
rect 17451 4233 17463 4267
rect 17862 4264 17868 4276
rect 17823 4236 17868 4264
rect 17405 4227 17463 4233
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 18874 4224 18880 4276
rect 18932 4264 18938 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18932 4236 19073 4264
rect 18932 4224 18938 4236
rect 19061 4233 19073 4236
rect 19107 4264 19119 4267
rect 19426 4264 19432 4276
rect 19107 4236 19432 4264
rect 19107 4233 19119 4236
rect 19061 4227 19119 4233
rect 19426 4224 19432 4236
rect 19484 4264 19490 4276
rect 20898 4264 20904 4276
rect 19484 4236 20904 4264
rect 19484 4224 19490 4236
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 9766 4196 9772 4208
rect 9727 4168 9772 4196
rect 9766 4156 9772 4168
rect 9824 4156 9830 4208
rect 14369 4199 14427 4205
rect 14369 4196 14381 4199
rect 13556 4168 14381 4196
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9732 4100 10057 4128
rect 9732 4088 9738 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 13449 4131 13507 4137
rect 13449 4097 13461 4131
rect 13495 4128 13507 4131
rect 13556 4128 13584 4168
rect 14369 4165 14381 4168
rect 14415 4196 14427 4199
rect 15654 4196 15660 4208
rect 14415 4168 15660 4196
rect 14415 4165 14427 4168
rect 14369 4159 14427 4165
rect 15654 4156 15660 4168
rect 15712 4156 15718 4208
rect 19978 4196 19984 4208
rect 19536 4168 19984 4196
rect 13722 4128 13728 4140
rect 13495 4100 13584 4128
rect 13683 4100 13728 4128
rect 13495 4097 13507 4100
rect 13449 4091 13507 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19536 4137 19564 4168
rect 19978 4156 19984 4168
rect 20036 4156 20042 4208
rect 20070 4156 20076 4208
rect 20128 4196 20134 4208
rect 20165 4199 20223 4205
rect 20165 4196 20177 4199
rect 20128 4168 20177 4196
rect 20128 4156 20134 4168
rect 20165 4165 20177 4168
rect 20211 4165 20223 4199
rect 20165 4159 20223 4165
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 18840 4100 19533 4128
rect 18840 4088 18846 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19521 4091 19579 4097
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 20990 4128 20996 4140
rect 20855 4100 20996 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 8021 4063 8079 4069
rect 7892 4032 7937 4060
rect 7892 4020 7898 4032
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 8067 4032 8769 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8757 4029 8769 4032
rect 8803 4060 8815 4063
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 8803 4032 9321 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 10686 4020 10692 4072
rect 10744 4060 10750 4072
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10744 4032 10793 4060
rect 10744 4020 10750 4032
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 10781 4023 10839 4029
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 15746 4060 15752 4072
rect 15707 4032 15752 4060
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 16022 4020 16028 4072
rect 16080 4060 16086 4072
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 16080 4032 16221 4060
rect 16080 4020 16086 4032
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 18084 4063 18142 4069
rect 18084 4029 18096 4063
rect 18130 4029 18142 4063
rect 18084 4023 18142 4029
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 11388 3964 11529 3992
rect 11388 3952 11394 3964
rect 11517 3961 11529 3964
rect 11563 3992 11575 3995
rect 12161 3995 12219 4001
rect 12161 3992 12173 3995
rect 11563 3964 12173 3992
rect 11563 3961 11575 3964
rect 11517 3955 11575 3961
rect 12161 3961 12173 3964
rect 12207 3961 12219 3995
rect 12161 3955 12219 3961
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3992 13599 3995
rect 13814 3992 13820 4004
rect 13587 3964 13820 3992
rect 13587 3961 13599 3964
rect 13541 3955 13599 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 15562 3952 15568 4004
rect 15620 3992 15626 4004
rect 18099 3992 18127 4023
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 15620 3964 18521 3992
rect 15620 3952 15626 3964
rect 18509 3961 18521 3964
rect 18555 3961 18567 3995
rect 19242 3992 19248 4004
rect 19203 3964 19248 3992
rect 18509 3955 18567 3961
rect 19242 3952 19248 3964
rect 19300 3952 19306 4004
rect 19337 3995 19395 4001
rect 19337 3961 19349 3995
rect 19383 3992 19395 3995
rect 19426 3992 19432 4004
rect 19383 3964 19432 3992
rect 19383 3961 19395 3964
rect 19337 3955 19395 3961
rect 19426 3952 19432 3964
rect 19484 3952 19490 4004
rect 20898 3952 20904 4004
rect 20956 3992 20962 4004
rect 21450 3992 21456 4004
rect 20956 3964 21001 3992
rect 21411 3964 21456 3992
rect 20956 3952 20962 3964
rect 21450 3952 21456 3964
rect 21508 3952 21514 4004
rect 8018 3924 8024 3936
rect 7760 3896 8024 3924
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 17126 3924 17132 3936
rect 13504 3896 17132 3924
rect 13504 3884 13510 3896
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 18187 3927 18245 3933
rect 18187 3924 18199 3927
rect 17276 3896 18199 3924
rect 17276 3884 17282 3896
rect 18187 3893 18199 3896
rect 18233 3893 18245 3927
rect 18187 3887 18245 3893
rect 20625 3927 20683 3933
rect 20625 3893 20637 3927
rect 20671 3924 20683 3927
rect 20916 3924 20944 3952
rect 20671 3896 20944 3924
rect 20671 3893 20683 3896
rect 20625 3887 20683 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11238 3720 11244 3732
rect 10919 3692 11244 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 13630 3720 13636 3732
rect 13591 3692 13636 3720
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 15746 3720 15752 3732
rect 15707 3692 15752 3720
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 18923 3723 18981 3729
rect 18923 3689 18935 3723
rect 18969 3720 18981 3723
rect 19242 3720 19248 3732
rect 18969 3692 19248 3720
rect 18969 3689 18981 3692
rect 18923 3683 18981 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 3099 3655 3157 3661
rect 3099 3621 3111 3655
rect 3145 3652 3157 3655
rect 8662 3652 8668 3664
rect 3145 3624 8668 3652
rect 3145 3621 3157 3624
rect 3099 3615 3157 3621
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 8757 3655 8815 3661
rect 8757 3621 8769 3655
rect 8803 3652 8815 3655
rect 9122 3652 9128 3664
rect 8803 3624 9128 3652
rect 8803 3621 8815 3624
rect 8757 3615 8815 3621
rect 9122 3612 9128 3624
rect 9180 3612 9186 3664
rect 13449 3655 13507 3661
rect 13449 3621 13461 3655
rect 13495 3652 13507 3655
rect 13814 3652 13820 3664
rect 13495 3624 13820 3652
rect 13495 3621 13507 3624
rect 13449 3615 13507 3621
rect 13814 3612 13820 3624
rect 13872 3612 13878 3664
rect 15427 3655 15485 3661
rect 15427 3621 15439 3655
rect 15473 3652 15485 3655
rect 16206 3652 16212 3664
rect 15473 3624 16212 3652
rect 15473 3621 15485 3624
rect 15427 3615 15485 3621
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 16390 3652 16396 3664
rect 16351 3624 16396 3652
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 17310 3652 17316 3664
rect 17271 3624 17316 3652
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 2996 3587 3054 3593
rect 2996 3553 3008 3587
rect 3042 3553 3054 3587
rect 8018 3584 8024 3596
rect 7979 3556 8024 3584
rect 2996 3547 3054 3553
rect 3011 3516 3039 3547
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8297 3587 8355 3593
rect 8297 3553 8309 3587
rect 8343 3584 8355 3587
rect 8386 3584 8392 3596
rect 8343 3556 8392 3584
rect 8343 3553 8355 3556
rect 8297 3547 8355 3553
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 12688 3587 12746 3593
rect 12688 3553 12700 3587
rect 12734 3584 12746 3587
rect 13078 3584 13084 3596
rect 12734 3556 13084 3584
rect 12734 3553 12746 3556
rect 12688 3547 12746 3553
rect 13078 3544 13084 3556
rect 13136 3584 13142 3596
rect 13722 3584 13728 3596
rect 13136 3556 13728 3584
rect 13136 3544 13142 3556
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 15197 3587 15255 3593
rect 15197 3553 15209 3587
rect 15243 3584 15255 3587
rect 15286 3584 15292 3596
rect 15243 3556 15292 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3584 20867 3587
rect 20990 3584 20996 3596
rect 20855 3556 20996 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 3142 3516 3148 3528
rect 3011 3488 3148 3516
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 17218 3516 17224 3528
rect 17179 3488 17224 3516
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17494 3476 17500 3488
rect 17552 3516 17558 3528
rect 21450 3516 21456 3528
rect 17552 3488 21456 3516
rect 17552 3476 17558 3488
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 5500 3420 7757 3448
rect 5500 3408 5506 3420
rect 7745 3417 7757 3420
rect 7791 3448 7803 3451
rect 7834 3448 7840 3460
rect 7791 3420 7840 3448
rect 7791 3417 7803 3420
rect 7745 3411 7803 3417
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 8110 3448 8116 3460
rect 8071 3420 8116 3448
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 12759 3383 12817 3389
rect 12759 3380 12771 3383
rect 12492 3352 12771 3380
rect 12492 3340 12498 3352
rect 12759 3349 12771 3352
rect 12805 3349 12817 3383
rect 12759 3343 12817 3349
rect 18693 3383 18751 3389
rect 18693 3349 18705 3383
rect 18739 3380 18751 3383
rect 18782 3380 18788 3392
rect 18739 3352 18788 3380
rect 18739 3349 18751 3352
rect 18693 3343 18751 3349
rect 18782 3340 18788 3352
rect 18840 3380 18846 3392
rect 20622 3380 20628 3392
rect 18840 3352 20628 3380
rect 18840 3340 18846 3352
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 10100 3148 10149 3176
rect 10100 3136 10106 3148
rect 10137 3145 10149 3148
rect 10183 3145 10195 3179
rect 13078 3176 13084 3188
rect 13039 3148 13084 3176
rect 10137 3139 10195 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 13771 3179 13829 3185
rect 13771 3145 13783 3179
rect 13817 3176 13829 3179
rect 13998 3176 14004 3188
rect 13817 3148 14004 3176
rect 13817 3145 13829 3148
rect 13771 3139 13829 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 17221 3179 17279 3185
rect 17221 3145 17233 3179
rect 17267 3176 17279 3179
rect 17310 3176 17316 3188
rect 17267 3148 17316 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 20395 3179 20453 3185
rect 20395 3145 20407 3179
rect 20441 3176 20453 3179
rect 20806 3176 20812 3188
rect 20441 3148 20812 3176
rect 20441 3145 20453 3148
rect 20395 3139 20453 3145
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 20990 3176 20996 3188
rect 20951 3148 20996 3176
rect 20990 3136 20996 3148
rect 21048 3136 21054 3188
rect 22462 3136 22468 3188
rect 22520 3176 22526 3188
rect 23891 3179 23949 3185
rect 23891 3176 23903 3179
rect 22520 3148 23903 3176
rect 22520 3136 22526 3148
rect 23891 3145 23903 3148
rect 23937 3145 23949 3179
rect 23891 3139 23949 3145
rect 7285 3111 7343 3117
rect 7285 3077 7297 3111
rect 7331 3108 7343 3111
rect 8110 3108 8116 3120
rect 7331 3080 8116 3108
rect 7331 3077 7343 3080
rect 7285 3071 7343 3077
rect 8110 3068 8116 3080
rect 8168 3108 8174 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 8168 3080 8217 3108
rect 8168 3068 8174 3080
rect 8205 3077 8217 3080
rect 8251 3108 8263 3111
rect 9125 3111 9183 3117
rect 9125 3108 9137 3111
rect 8251 3080 9137 3108
rect 8251 3077 8263 3080
rect 8205 3071 8263 3077
rect 9125 3077 9137 3080
rect 9171 3077 9183 3111
rect 9125 3071 9183 3077
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 9582 3040 9588 3052
rect 8895 3012 9588 3040
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 17218 3000 17224 3052
rect 17276 3040 17282 3052
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17276 3012 17509 3040
rect 17276 3000 17282 3012
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 18138 3040 18144 3052
rect 18095 3012 18144 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2941 8171 2975
rect 8386 2972 8392 2984
rect 8347 2944 8392 2972
rect 8113 2935 8171 2941
rect 8128 2904 8156 2935
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 9744 2975 9802 2981
rect 9744 2941 9756 2975
rect 9790 2972 9802 2975
rect 10042 2972 10048 2984
rect 9790 2944 10048 2972
rect 9790 2941 9802 2944
rect 9744 2935 9802 2941
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 12253 2975 12311 2981
rect 12253 2941 12265 2975
rect 12299 2972 12311 2975
rect 12434 2972 12440 2984
rect 12299 2944 12440 2972
rect 12299 2941 12311 2944
rect 12253 2935 12311 2941
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 13668 2975 13726 2981
rect 13668 2972 13680 2975
rect 12584 2944 13680 2972
rect 12584 2932 12590 2944
rect 13668 2941 13680 2944
rect 13714 2972 13726 2975
rect 20165 2975 20223 2981
rect 13714 2944 13814 2972
rect 13714 2941 13726 2944
rect 13668 2935 13726 2941
rect 8846 2904 8852 2916
rect 8128 2876 8852 2904
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3142 2836 3148 2848
rect 3099 2808 3148 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 7558 2836 7564 2848
rect 7519 2808 7564 2836
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 9815 2839 9873 2845
rect 9815 2836 9827 2839
rect 9272 2808 9827 2836
rect 9272 2796 9278 2808
rect 9815 2805 9827 2808
rect 9861 2805 9873 2839
rect 9815 2799 9873 2805
rect 12621 2839 12679 2845
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 12894 2836 12900 2848
rect 12667 2808 12900 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 13786 2836 13814 2944
rect 20165 2941 20177 2975
rect 20211 2972 20223 2975
rect 20324 2975 20382 2981
rect 20324 2972 20336 2975
rect 20211 2944 20336 2972
rect 20211 2941 20223 2944
rect 20165 2935 20223 2941
rect 20324 2941 20336 2944
rect 20370 2972 20382 2975
rect 21358 2972 21364 2984
rect 20370 2944 21364 2972
rect 20370 2941 20382 2944
rect 20324 2935 20382 2941
rect 21358 2932 21364 2944
rect 21416 2932 21422 2984
rect 23820 2975 23878 2981
rect 23820 2941 23832 2975
rect 23866 2972 23878 2975
rect 23866 2944 24348 2972
rect 23866 2941 23878 2944
rect 23820 2935 23878 2941
rect 14182 2836 14188 2848
rect 13786 2808 14188 2836
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 18782 2836 18788 2848
rect 18743 2808 18788 2836
rect 18782 2796 18788 2808
rect 18840 2796 18846 2848
rect 24320 2845 24348 2944
rect 24305 2839 24363 2845
rect 24305 2805 24317 2839
rect 24351 2836 24363 2839
rect 25406 2836 25412 2848
rect 24351 2808 25412 2836
rect 24351 2805 24363 2808
rect 24305 2799 24363 2805
rect 25406 2796 25412 2808
rect 25464 2796 25470 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 7558 2592 7564 2644
rect 7616 2632 7622 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7616 2604 8125 2632
rect 7616 2592 7622 2604
rect 8113 2601 8125 2604
rect 8159 2632 8171 2635
rect 8386 2632 8392 2644
rect 8159 2604 8392 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 8938 2592 8944 2644
rect 8996 2632 9002 2644
rect 9999 2635 10057 2641
rect 9999 2632 10011 2635
rect 8996 2604 10011 2632
rect 8996 2592 9002 2604
rect 9999 2601 10011 2604
rect 10045 2601 10057 2635
rect 9999 2595 10057 2601
rect 19751 2635 19809 2641
rect 19751 2601 19763 2635
rect 19797 2632 19809 2635
rect 21266 2632 21272 2644
rect 19797 2604 21272 2632
rect 19797 2601 19809 2604
rect 19751 2595 19809 2601
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 21499 2635 21557 2641
rect 21499 2601 21511 2635
rect 21545 2632 21557 2635
rect 21910 2632 21916 2644
rect 21545 2604 21916 2632
rect 21545 2601 21557 2604
rect 21499 2595 21557 2601
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 22787 2635 22845 2641
rect 22787 2632 22799 2635
rect 22336 2604 22799 2632
rect 22336 2592 22342 2604
rect 22787 2601 22799 2604
rect 22833 2601 22845 2635
rect 22787 2595 22845 2601
rect 8846 2524 8852 2576
rect 8904 2564 8910 2576
rect 9033 2567 9091 2573
rect 9033 2564 9045 2567
rect 8904 2536 9045 2564
rect 8904 2524 8910 2536
rect 9033 2533 9045 2536
rect 9079 2533 9091 2567
rect 9033 2527 9091 2533
rect 22186 2524 22192 2576
rect 22244 2564 22250 2576
rect 24167 2567 24225 2573
rect 24167 2564 24179 2567
rect 22244 2536 24179 2564
rect 22244 2524 22250 2536
rect 24167 2533 24179 2536
rect 24213 2533 24225 2567
rect 24167 2527 24225 2533
rect 7837 2499 7895 2505
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7883 2468 8401 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 8389 2465 8401 2468
rect 8435 2496 8447 2499
rect 9214 2496 9220 2508
rect 8435 2468 9220 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9928 2499 9986 2505
rect 9928 2465 9940 2499
rect 9974 2496 9986 2499
rect 13541 2499 13599 2505
rect 9974 2468 10456 2496
rect 9974 2465 9986 2468
rect 9928 2459 9986 2465
rect 8573 2363 8631 2369
rect 8573 2329 8585 2363
rect 8619 2360 8631 2363
rect 9122 2360 9128 2372
rect 8619 2332 9128 2360
rect 8619 2329 8631 2332
rect 8573 2323 8631 2329
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 10428 2301 10456 2468
rect 13541 2465 13553 2499
rect 13587 2496 13599 2499
rect 14182 2496 14188 2508
rect 13587 2468 14188 2496
rect 13587 2465 13599 2468
rect 13541 2459 13599 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 19680 2499 19738 2505
rect 19680 2465 19692 2499
rect 19726 2496 19738 2499
rect 20070 2496 20076 2508
rect 19726 2468 20076 2496
rect 19726 2465 19738 2468
rect 19680 2459 19738 2465
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 21428 2499 21486 2505
rect 21428 2465 21440 2499
rect 21474 2496 21486 2499
rect 22716 2499 22774 2505
rect 21474 2468 21956 2496
rect 21474 2465 21486 2468
rect 21428 2459 21486 2465
rect 13725 2363 13783 2369
rect 13725 2329 13737 2363
rect 13771 2360 13783 2363
rect 14366 2360 14372 2372
rect 13771 2332 14372 2360
rect 13771 2329 13783 2332
rect 13725 2323 13783 2329
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 10413 2295 10471 2301
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 11422 2292 11428 2304
rect 10459 2264 11428 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 11422 2252 11428 2264
rect 11480 2252 11486 2304
rect 14182 2292 14188 2304
rect 14095 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2292 14246 2304
rect 15654 2292 15660 2304
rect 14240 2264 15660 2292
rect 14240 2252 14246 2264
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 20070 2292 20076 2304
rect 20031 2264 20076 2292
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 21928 2301 21956 2468
rect 22716 2465 22728 2499
rect 22762 2496 22774 2499
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22762 2468 23121 2496
rect 22762 2465 22774 2468
rect 22716 2459 22774 2465
rect 23109 2465 23121 2468
rect 23155 2496 23167 2499
rect 24080 2499 24138 2505
rect 23155 2468 23474 2496
rect 23155 2465 23167 2468
rect 23109 2459 23167 2465
rect 23446 2428 23474 2468
rect 24080 2465 24092 2499
rect 24126 2496 24138 2499
rect 24126 2468 24624 2496
rect 24126 2465 24138 2468
rect 24080 2459 24138 2465
rect 24210 2428 24216 2440
rect 23446 2400 24216 2428
rect 24210 2388 24216 2400
rect 24268 2388 24274 2440
rect 21913 2295 21971 2301
rect 21913 2261 21925 2295
rect 21959 2292 21971 2295
rect 22646 2292 22652 2304
rect 21959 2264 22652 2292
rect 21959 2261 21971 2264
rect 21913 2255 21971 2261
rect 22646 2252 22652 2264
rect 22704 2252 22710 2304
rect 24596 2301 24624 2468
rect 24581 2295 24639 2301
rect 24581 2261 24593 2295
rect 24627 2292 24639 2295
rect 26878 2292 26884 2304
rect 24627 2264 26884 2292
rect 24627 2261 24639 2264
rect 24581 2255 24639 2261
rect 26878 2252 26884 2264
rect 26936 2252 26942 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 6178 76 6184 128
rect 6236 116 6242 128
rect 7466 116 7472 128
rect 6236 88 7472 116
rect 6236 76 6242 88
rect 7466 76 7472 88
rect 7524 76 7530 128
<< via1 >>
rect 19248 27480 19300 27532
rect 19892 27480 19944 27532
rect 24860 27480 24912 27532
rect 25780 27480 25832 27532
rect 26240 27480 26292 27532
rect 27252 27480 27304 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 15476 24556 15528 24608
rect 19064 24556 19116 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 21364 24216 21416 24268
rect 21548 24012 21600 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 11060 23808 11112 23860
rect 12624 23851 12676 23860
rect 12624 23817 12633 23851
rect 12633 23817 12667 23851
rect 12667 23817 12676 23851
rect 12624 23808 12676 23817
rect 13728 23851 13780 23860
rect 13728 23817 13737 23851
rect 13737 23817 13771 23851
rect 13771 23817 13780 23851
rect 13728 23808 13780 23817
rect 21088 23808 21140 23860
rect 21364 23808 21416 23860
rect 22560 23851 22612 23860
rect 22560 23817 22569 23851
rect 22569 23817 22603 23851
rect 22603 23817 22612 23851
rect 22560 23808 22612 23817
rect 1124 23672 1176 23724
rect 6092 23604 6144 23656
rect 11520 23604 11572 23656
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 19064 23604 19116 23656
rect 22008 23740 22060 23792
rect 22560 23604 22612 23656
rect 21272 23536 21324 23588
rect 1768 23468 1820 23520
rect 22836 23468 22888 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 112 23264 164 23316
rect 1676 23128 1728 23180
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 12900 22763 12952 22772
rect 12900 22729 12909 22763
rect 12909 22729 12943 22763
rect 12943 22729 12952 22763
rect 12900 22720 12952 22729
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 15752 22720 15804 22772
rect 16948 22720 17000 22772
rect 18052 22380 18104 22432
rect 18604 22423 18656 22432
rect 18604 22389 18613 22423
rect 18613 22389 18647 22423
rect 18647 22389 18656 22423
rect 18604 22380 18656 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 7104 20204 7156 20256
rect 8668 20204 8720 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 13544 20000 13596 20052
rect 5172 19864 5224 19916
rect 6644 19864 6696 19916
rect 13176 19864 13228 19916
rect 8484 19771 8536 19780
rect 8484 19737 8493 19771
rect 8493 19737 8527 19771
rect 8527 19737 8536 19771
rect 8484 19728 8536 19737
rect 7196 19660 7248 19712
rect 7840 19660 7892 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 6092 19456 6144 19508
rect 7840 19499 7892 19508
rect 7840 19465 7849 19499
rect 7849 19465 7883 19499
rect 7883 19465 7892 19499
rect 7840 19456 7892 19465
rect 9588 19499 9640 19508
rect 9588 19465 9597 19499
rect 9597 19465 9631 19499
rect 9631 19465 9640 19499
rect 9588 19456 9640 19465
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 3884 19252 3936 19304
rect 7656 19320 7708 19372
rect 8576 19320 8628 19372
rect 2504 19116 2556 19168
rect 7840 19252 7892 19304
rect 9588 19252 9640 19304
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 8484 19184 8536 19236
rect 9864 19184 9916 19236
rect 25136 19252 25188 19304
rect 6460 19116 6512 19168
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 6644 19116 6696 19125
rect 6920 19159 6972 19168
rect 6920 19125 6929 19159
rect 6929 19125 6963 19159
rect 6963 19125 6972 19159
rect 6920 19116 6972 19125
rect 7012 19116 7064 19168
rect 8944 19116 8996 19168
rect 11704 19116 11756 19168
rect 12348 19116 12400 19168
rect 12716 19159 12768 19168
rect 12716 19125 12725 19159
rect 12725 19125 12759 19159
rect 12759 19125 12768 19159
rect 12716 19116 12768 19125
rect 16764 19116 16816 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1492 18912 1544 18964
rect 112 18844 164 18896
rect 7012 18912 7064 18964
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 6368 18887 6420 18896
rect 6368 18853 6377 18887
rect 6377 18853 6411 18887
rect 6411 18853 6420 18887
rect 6368 18844 6420 18853
rect 7656 18844 7708 18896
rect 7840 18887 7892 18896
rect 7840 18853 7849 18887
rect 7849 18853 7883 18887
rect 7883 18853 7892 18887
rect 7840 18844 7892 18853
rect 7932 18887 7984 18896
rect 7932 18853 7941 18887
rect 7941 18853 7975 18887
rect 7975 18853 7984 18887
rect 7932 18844 7984 18853
rect 10140 18844 10192 18896
rect 11704 18844 11756 18896
rect 12256 18887 12308 18896
rect 12256 18853 12265 18887
rect 12265 18853 12299 18887
rect 12299 18853 12308 18887
rect 12256 18844 12308 18853
rect 12440 18844 12492 18896
rect 1952 18776 2004 18828
rect 5172 18776 5224 18828
rect 13912 18776 13964 18828
rect 19340 18776 19392 18828
rect 24216 18776 24268 18828
rect 6276 18751 6328 18760
rect 6276 18717 6285 18751
rect 6285 18717 6319 18751
rect 6319 18717 6328 18751
rect 6276 18708 6328 18717
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 9864 18708 9916 18760
rect 10968 18708 11020 18760
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 12808 18683 12860 18692
rect 12808 18649 12817 18683
rect 12817 18649 12851 18683
rect 12851 18649 12860 18683
rect 12808 18640 12860 18649
rect 4804 18572 4856 18624
rect 7748 18572 7800 18624
rect 8300 18572 8352 18624
rect 12532 18572 12584 18624
rect 19892 18572 19944 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 5172 18411 5224 18420
rect 5172 18377 5181 18411
rect 5181 18377 5215 18411
rect 5215 18377 5224 18411
rect 5172 18368 5224 18377
rect 6368 18368 6420 18420
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 12716 18411 12768 18420
rect 12716 18377 12725 18411
rect 12725 18377 12759 18411
rect 12759 18377 12768 18411
rect 12716 18368 12768 18377
rect 13912 18411 13964 18420
rect 13912 18377 13921 18411
rect 13921 18377 13955 18411
rect 13955 18377 13964 18411
rect 19340 18411 19392 18420
rect 13912 18368 13964 18377
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 19340 18368 19392 18377
rect 24768 18411 24820 18420
rect 24768 18377 24777 18411
rect 24777 18377 24811 18411
rect 24811 18377 24820 18411
rect 24768 18368 24820 18377
rect 7564 18300 7616 18352
rect 7748 18300 7800 18352
rect 7196 18232 7248 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 9772 18300 9824 18352
rect 17040 18300 17092 18352
rect 9588 18232 9640 18284
rect 1492 18164 1544 18216
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 17500 18232 17552 18284
rect 19892 18275 19944 18284
rect 3332 18096 3384 18148
rect 1676 18028 1728 18080
rect 4712 18071 4764 18080
rect 4712 18037 4721 18071
rect 4721 18037 4755 18071
rect 4755 18037 4764 18071
rect 4712 18028 4764 18037
rect 16304 18164 16356 18216
rect 16580 18164 16632 18216
rect 7380 18096 7432 18148
rect 8484 18096 8536 18148
rect 6368 18028 6420 18080
rect 7932 18028 7984 18080
rect 9772 18096 9824 18148
rect 11612 18096 11664 18148
rect 18328 18139 18380 18148
rect 10140 18028 10192 18080
rect 12440 18028 12492 18080
rect 12716 18028 12768 18080
rect 18328 18105 18337 18139
rect 18337 18105 18371 18139
rect 18371 18105 18380 18139
rect 18328 18096 18380 18105
rect 19892 18241 19901 18275
rect 19901 18241 19935 18275
rect 19935 18241 19944 18275
rect 19892 18232 19944 18241
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 24216 18164 24268 18216
rect 14280 18028 14332 18080
rect 18236 18028 18288 18080
rect 21364 18096 21416 18148
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 7840 17824 7892 17876
rect 8944 17867 8996 17876
rect 8944 17833 8953 17867
rect 8953 17833 8987 17867
rect 8987 17833 8996 17867
rect 8944 17824 8996 17833
rect 11612 17867 11664 17876
rect 11612 17833 11621 17867
rect 11621 17833 11655 17867
rect 11655 17833 11664 17867
rect 11612 17824 11664 17833
rect 12256 17867 12308 17876
rect 12256 17833 12265 17867
rect 12265 17833 12299 17867
rect 12299 17833 12308 17867
rect 12256 17824 12308 17833
rect 17040 17867 17092 17876
rect 17040 17833 17049 17867
rect 17049 17833 17083 17867
rect 17083 17833 17092 17867
rect 17040 17824 17092 17833
rect 18328 17867 18380 17876
rect 18328 17833 18337 17867
rect 18337 17833 18371 17867
rect 18371 17833 18380 17867
rect 18328 17824 18380 17833
rect 19984 17824 20036 17876
rect 20168 17867 20220 17876
rect 20168 17833 20177 17867
rect 20177 17833 20211 17867
rect 20211 17833 20220 17867
rect 20168 17824 20220 17833
rect 21548 17867 21600 17876
rect 21548 17833 21557 17867
rect 21557 17833 21591 17867
rect 21591 17833 21600 17867
rect 21548 17824 21600 17833
rect 25504 17824 25556 17876
rect 6920 17756 6972 17808
rect 7380 17799 7432 17808
rect 7380 17765 7389 17799
rect 7389 17765 7423 17799
rect 7423 17765 7432 17799
rect 7380 17756 7432 17765
rect 7656 17756 7708 17808
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 12348 17756 12400 17808
rect 13544 17756 13596 17808
rect 17500 17756 17552 17808
rect 18420 17756 18472 17808
rect 19156 17756 19208 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2596 17688 2648 17740
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 22468 17688 22520 17740
rect 24216 17688 24268 17740
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 8484 17620 8536 17672
rect 10600 17620 10652 17672
rect 12808 17620 12860 17672
rect 13176 17663 13228 17672
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13176 17620 13228 17629
rect 13360 17620 13412 17672
rect 18512 17620 18564 17672
rect 1768 17552 1820 17604
rect 8208 17552 8260 17604
rect 10968 17552 11020 17604
rect 3608 17484 3660 17536
rect 5080 17527 5132 17536
rect 5080 17493 5089 17527
rect 5089 17493 5123 17527
rect 5123 17493 5132 17527
rect 5080 17484 5132 17493
rect 7656 17484 7708 17536
rect 15936 17484 15988 17536
rect 18420 17484 18472 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 4712 17280 4764 17332
rect 5080 17280 5132 17332
rect 5448 17280 5500 17332
rect 6368 17280 6420 17332
rect 6552 17323 6604 17332
rect 6552 17289 6561 17323
rect 6561 17289 6595 17323
rect 6595 17289 6604 17323
rect 6552 17280 6604 17289
rect 9496 17280 9548 17332
rect 9864 17280 9916 17332
rect 10600 17323 10652 17332
rect 10600 17289 10609 17323
rect 10609 17289 10643 17323
rect 10643 17289 10652 17323
rect 10600 17280 10652 17289
rect 11520 17280 11572 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 17500 17280 17552 17332
rect 17684 17280 17736 17332
rect 112 17144 164 17196
rect 2596 17144 2648 17196
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 7104 17212 7156 17264
rect 7748 17255 7800 17264
rect 7748 17221 7757 17255
rect 7757 17221 7791 17255
rect 7791 17221 7800 17255
rect 7748 17212 7800 17221
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 22468 17280 22520 17332
rect 24216 17280 24268 17332
rect 20536 17255 20588 17264
rect 20536 17221 20545 17255
rect 20545 17221 20579 17255
rect 20579 17221 20588 17255
rect 20536 17212 20588 17221
rect 21732 17212 21784 17264
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 20168 17144 20220 17196
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 1400 17076 1452 17128
rect 3332 17076 3384 17128
rect 12348 17076 12400 17128
rect 13176 17076 13228 17128
rect 15660 17119 15712 17128
rect 15660 17085 15669 17119
rect 15669 17085 15703 17119
rect 15703 17085 15712 17119
rect 15660 17076 15712 17085
rect 3976 17008 4028 17060
rect 4988 17008 5040 17060
rect 1492 16940 1544 16992
rect 2688 16940 2740 16992
rect 5080 16940 5132 16992
rect 6460 17008 6512 17060
rect 6552 17008 6604 17060
rect 7932 17008 7984 17060
rect 9772 17051 9824 17060
rect 9772 17017 9781 17051
rect 9781 17017 9815 17051
rect 9815 17017 9824 17051
rect 9772 17008 9824 17017
rect 10876 17008 10928 17060
rect 8852 16940 8904 16992
rect 15568 17051 15620 17060
rect 15568 17017 15577 17051
rect 15577 17017 15611 17051
rect 15611 17017 15620 17051
rect 15568 17008 15620 17017
rect 18328 17051 18380 17060
rect 18328 17017 18337 17051
rect 18337 17017 18371 17051
rect 18371 17017 18380 17051
rect 18328 17008 18380 17017
rect 20076 17051 20128 17060
rect 20076 17017 20085 17051
rect 20085 17017 20119 17051
rect 20119 17017 20128 17051
rect 21364 17051 21416 17060
rect 20076 17008 20128 17017
rect 21364 17017 21373 17051
rect 21373 17017 21407 17051
rect 21407 17017 21416 17051
rect 21364 17008 21416 17017
rect 22192 17051 22244 17060
rect 22192 17017 22201 17051
rect 22201 17017 22235 17051
rect 22235 17017 22244 17051
rect 22192 17008 22244 17017
rect 13544 16983 13596 16992
rect 13544 16949 13553 16983
rect 13553 16949 13587 16983
rect 13587 16949 13596 16983
rect 13544 16940 13596 16949
rect 19156 16983 19208 16992
rect 19156 16949 19165 16983
rect 19165 16949 19199 16983
rect 19199 16949 19208 16983
rect 19156 16940 19208 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1676 16736 1728 16788
rect 6920 16736 6972 16788
rect 10048 16779 10100 16788
rect 10048 16745 10057 16779
rect 10057 16745 10091 16779
rect 10091 16745 10100 16779
rect 10048 16736 10100 16745
rect 10140 16736 10192 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 17040 16779 17092 16788
rect 17040 16745 17049 16779
rect 17049 16745 17083 16779
rect 17083 16745 17092 16779
rect 17040 16736 17092 16745
rect 17500 16736 17552 16788
rect 19156 16736 19208 16788
rect 4804 16711 4856 16720
rect 4804 16677 4813 16711
rect 4813 16677 4847 16711
rect 4847 16677 4856 16711
rect 4804 16668 4856 16677
rect 6368 16711 6420 16720
rect 6368 16677 6377 16711
rect 6377 16677 6411 16711
rect 6411 16677 6420 16711
rect 6368 16668 6420 16677
rect 7564 16668 7616 16720
rect 7932 16711 7984 16720
rect 7932 16677 7941 16711
rect 7941 16677 7975 16711
rect 7975 16677 7984 16711
rect 7932 16668 7984 16677
rect 11612 16668 11664 16720
rect 13452 16711 13504 16720
rect 13452 16677 13461 16711
rect 13461 16677 13495 16711
rect 13495 16677 13504 16711
rect 13452 16668 13504 16677
rect 15568 16668 15620 16720
rect 19432 16711 19484 16720
rect 19432 16677 19441 16711
rect 19441 16677 19475 16711
rect 19475 16677 19484 16711
rect 19432 16668 19484 16677
rect 20536 16668 20588 16720
rect 21088 16711 21140 16720
rect 21088 16677 21097 16711
rect 21097 16677 21131 16711
rect 21131 16677 21140 16711
rect 21088 16668 21140 16677
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 13176 16600 13228 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 22008 16600 22060 16652
rect 22468 16643 22520 16652
rect 22468 16609 22477 16643
rect 22477 16609 22511 16643
rect 22511 16609 22520 16643
rect 22468 16600 22520 16609
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 6460 16532 6512 16584
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 9404 16532 9456 16584
rect 12072 16532 12124 16584
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 12348 16464 12400 16516
rect 14004 16532 14056 16584
rect 16488 16532 16540 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 18512 16532 18564 16584
rect 20720 16532 20772 16584
rect 18328 16464 18380 16516
rect 18972 16464 19024 16516
rect 20168 16464 20220 16516
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 3976 16396 4028 16448
rect 4344 16396 4396 16448
rect 7748 16396 7800 16448
rect 8484 16396 8536 16448
rect 10876 16439 10928 16448
rect 10876 16405 10885 16439
rect 10885 16405 10919 16439
rect 10919 16405 10928 16439
rect 10876 16396 10928 16405
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 5448 16192 5500 16244
rect 7932 16235 7984 16244
rect 7932 16201 7941 16235
rect 7941 16201 7975 16235
rect 7975 16201 7984 16235
rect 7932 16192 7984 16201
rect 9496 16235 9548 16244
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 9496 16192 9548 16201
rect 10048 16192 10100 16244
rect 11612 16192 11664 16244
rect 13452 16192 13504 16244
rect 15292 16192 15344 16244
rect 18512 16192 18564 16244
rect 19432 16192 19484 16244
rect 21088 16192 21140 16244
rect 22744 16192 22796 16244
rect 1676 16056 1728 16108
rect 1860 16056 1912 16108
rect 7104 16124 7156 16176
rect 10968 16167 11020 16176
rect 10968 16133 10977 16167
rect 10977 16133 11011 16167
rect 11011 16133 11020 16167
rect 10968 16124 11020 16133
rect 13360 16124 13412 16176
rect 14004 16167 14056 16176
rect 14004 16133 14013 16167
rect 14013 16133 14047 16167
rect 14047 16133 14056 16167
rect 14004 16124 14056 16133
rect 18420 16124 18472 16176
rect 4804 16056 4856 16108
rect 8116 16056 8168 16108
rect 10876 16056 10928 16108
rect 14372 16056 14424 16108
rect 16672 16056 16724 16108
rect 18880 16124 18932 16176
rect 21824 16124 21876 16176
rect 22560 16056 22612 16108
rect 4344 15988 4396 16040
rect 8484 15988 8536 16040
rect 14924 15988 14976 16040
rect 16028 16031 16080 16040
rect 16028 15997 16037 16031
rect 16037 15997 16071 16031
rect 16071 15997 16080 16031
rect 16028 15988 16080 15997
rect 16488 16031 16540 16040
rect 16488 15997 16497 16031
rect 16497 15997 16531 16031
rect 16531 15997 16540 16031
rect 16488 15988 16540 15997
rect 18972 15988 19024 16040
rect 1768 15920 1820 15972
rect 2412 15920 2464 15972
rect 4528 15920 4580 15972
rect 3332 15852 3384 15904
rect 4160 15852 4212 15904
rect 7748 15920 7800 15972
rect 10048 15920 10100 15972
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 10140 15895 10192 15904
rect 10140 15861 10149 15895
rect 10149 15861 10183 15895
rect 10183 15861 10192 15895
rect 10140 15852 10192 15861
rect 12072 15852 12124 15904
rect 13360 15852 13412 15904
rect 15660 15920 15712 15972
rect 13636 15852 13688 15904
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 15476 15852 15528 15904
rect 17040 15895 17092 15904
rect 17040 15861 17049 15895
rect 17049 15861 17083 15895
rect 17083 15861 17092 15895
rect 19432 15920 19484 15972
rect 21088 15920 21140 15972
rect 22192 15920 22244 15972
rect 22928 15920 22980 15972
rect 17040 15852 17092 15861
rect 22468 15895 22520 15904
rect 22468 15861 22477 15895
rect 22477 15861 22511 15895
rect 22511 15861 22520 15895
rect 22468 15852 22520 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 4712 15648 4764 15700
rect 4804 15648 4856 15700
rect 7012 15691 7064 15700
rect 7012 15657 7021 15691
rect 7021 15657 7055 15691
rect 7055 15657 7064 15691
rect 7012 15648 7064 15657
rect 7564 15648 7616 15700
rect 8852 15648 8904 15700
rect 9772 15648 9824 15700
rect 13544 15648 13596 15700
rect 1860 15623 1912 15632
rect 1860 15589 1869 15623
rect 1869 15589 1903 15623
rect 1903 15589 1912 15623
rect 2412 15623 2464 15632
rect 1860 15580 1912 15589
rect 2412 15589 2421 15623
rect 2421 15589 2455 15623
rect 2455 15589 2464 15623
rect 2412 15580 2464 15589
rect 3792 15580 3844 15632
rect 4160 15580 4212 15632
rect 10048 15623 10100 15632
rect 10048 15589 10051 15623
rect 10051 15589 10085 15623
rect 10085 15589 10100 15623
rect 10048 15580 10100 15589
rect 11612 15580 11664 15632
rect 14740 15648 14792 15700
rect 15844 15648 15896 15700
rect 16028 15691 16080 15700
rect 16028 15657 16037 15691
rect 16037 15657 16071 15691
rect 16071 15657 16080 15691
rect 16028 15648 16080 15657
rect 19156 15648 19208 15700
rect 19432 15691 19484 15700
rect 19432 15657 19441 15691
rect 19441 15657 19475 15691
rect 19475 15657 19484 15691
rect 19432 15648 19484 15657
rect 20076 15648 20128 15700
rect 20720 15691 20772 15700
rect 20720 15657 20729 15691
rect 20729 15657 20763 15691
rect 20763 15657 20772 15691
rect 20720 15648 20772 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 13912 15580 13964 15632
rect 16212 15580 16264 15632
rect 17040 15580 17092 15632
rect 21180 15623 21232 15632
rect 21180 15589 21189 15623
rect 21189 15589 21223 15623
rect 21223 15589 21232 15623
rect 21180 15580 21232 15589
rect 21732 15623 21784 15632
rect 21732 15589 21741 15623
rect 21741 15589 21775 15623
rect 21775 15589 21784 15623
rect 21732 15580 21784 15589
rect 22744 15623 22796 15632
rect 22744 15589 22753 15623
rect 22753 15589 22787 15623
rect 22787 15589 22796 15623
rect 22744 15580 22796 15589
rect 7932 15512 7984 15564
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 15752 15512 15804 15564
rect 16304 15512 16356 15564
rect 20168 15512 20220 15564
rect 24216 15512 24268 15564
rect 24768 15512 24820 15564
rect 27620 15512 27672 15564
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 9680 15487 9732 15496
rect 2964 15308 3016 15360
rect 4896 15308 4948 15360
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 6184 15351 6236 15360
rect 6184 15317 6193 15351
rect 6193 15317 6227 15351
rect 6227 15317 6236 15351
rect 6184 15308 6236 15317
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 17408 15444 17460 15496
rect 21088 15487 21140 15496
rect 12256 15376 12308 15428
rect 6920 15308 6972 15360
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 9404 15351 9456 15360
rect 9404 15317 9413 15351
rect 9413 15317 9447 15351
rect 9447 15317 9456 15351
rect 9404 15308 9456 15317
rect 10968 15351 11020 15360
rect 10968 15317 10977 15351
rect 10977 15317 11011 15351
rect 11011 15317 11020 15351
rect 10968 15308 11020 15317
rect 11244 15351 11296 15360
rect 11244 15317 11253 15351
rect 11253 15317 11287 15351
rect 11287 15317 11296 15351
rect 11244 15308 11296 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 14740 15308 14792 15360
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 22744 15444 22796 15496
rect 22928 15487 22980 15496
rect 22928 15453 22937 15487
rect 22937 15453 22971 15487
rect 22971 15453 22980 15487
rect 22928 15444 22980 15453
rect 19524 15308 19576 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1860 15104 1912 15156
rect 4896 15104 4948 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 10140 15104 10192 15156
rect 11612 15147 11664 15156
rect 11612 15113 11621 15147
rect 11621 15113 11655 15147
rect 11655 15113 11664 15147
rect 12164 15147 12216 15156
rect 11612 15104 11664 15113
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 13360 15147 13412 15156
rect 13360 15113 13369 15147
rect 13369 15113 13403 15147
rect 13403 15113 13412 15147
rect 13360 15104 13412 15113
rect 15752 15104 15804 15156
rect 16856 15104 16908 15156
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 18972 15147 19024 15156
rect 18972 15113 18981 15147
rect 18981 15113 19015 15147
rect 19015 15113 19024 15147
rect 18972 15104 19024 15113
rect 21180 15104 21232 15156
rect 22836 15147 22888 15156
rect 22836 15113 22845 15147
rect 22845 15113 22879 15147
rect 22879 15113 22888 15147
rect 22836 15104 22888 15113
rect 4068 15036 4120 15088
rect 3976 15011 4028 15020
rect 3976 14977 3985 15011
rect 3985 14977 4019 15011
rect 4019 14977 4028 15011
rect 3976 14968 4028 14977
rect 3424 14900 3476 14952
rect 4804 14968 4856 15020
rect 6184 14968 6236 15020
rect 6736 14968 6788 15020
rect 8760 14968 8812 15020
rect 9036 14968 9088 15020
rect 15844 15036 15896 15088
rect 14280 15011 14332 15020
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 14372 14968 14424 15020
rect 14648 14968 14700 15020
rect 19248 15036 19300 15088
rect 18052 15011 18104 15020
rect 18052 14977 18061 15011
rect 18061 14977 18095 15011
rect 18095 14977 18104 15011
rect 18052 14968 18104 14977
rect 20996 14968 21048 15020
rect 22744 14968 22796 15020
rect 3792 14875 3844 14884
rect 3792 14841 3801 14875
rect 3801 14841 3835 14875
rect 3835 14841 3844 14875
rect 3792 14832 3844 14841
rect 7012 14832 7064 14884
rect 7288 14832 7340 14884
rect 8392 14832 8444 14884
rect 9312 14832 9364 14884
rect 11244 14900 11296 14952
rect 12256 14900 12308 14952
rect 12164 14832 12216 14884
rect 12808 14832 12860 14884
rect 12992 14832 13044 14884
rect 13636 14832 13688 14884
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 10692 14807 10744 14816
rect 10692 14773 10701 14807
rect 10701 14773 10735 14807
rect 10735 14773 10744 14807
rect 10692 14764 10744 14773
rect 13912 14764 13964 14816
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 15660 14764 15712 14816
rect 16488 14900 16540 14952
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 20352 14832 20404 14884
rect 22192 14943 22244 14952
rect 22192 14909 22201 14943
rect 22201 14909 22235 14943
rect 22235 14909 22244 14943
rect 22192 14900 22244 14909
rect 27620 15036 27672 15088
rect 21088 14764 21140 14816
rect 21640 14807 21692 14816
rect 21640 14773 21649 14807
rect 21649 14773 21683 14807
rect 21683 14773 21692 14807
rect 21640 14764 21692 14773
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 24216 14764 24268 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1492 14560 1544 14612
rect 4068 14560 4120 14612
rect 6736 14603 6788 14612
rect 6736 14569 6745 14603
rect 6745 14569 6779 14603
rect 6779 14569 6788 14603
rect 6736 14560 6788 14569
rect 2320 14492 2372 14544
rect 8852 14560 8904 14612
rect 9312 14560 9364 14612
rect 9680 14560 9732 14612
rect 10692 14560 10744 14612
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 5080 14424 5132 14433
rect 5448 14467 5500 14476
rect 5448 14433 5457 14467
rect 5457 14433 5491 14467
rect 5491 14433 5500 14467
rect 5448 14424 5500 14433
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 2412 14356 2464 14408
rect 2872 14356 2924 14408
rect 7380 14424 7432 14476
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 9404 14492 9456 14544
rect 10968 14492 11020 14544
rect 13268 14560 13320 14612
rect 14280 14603 14332 14612
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 14740 14603 14792 14612
rect 14740 14569 14749 14603
rect 14749 14569 14783 14603
rect 14783 14569 14792 14603
rect 14740 14560 14792 14569
rect 16488 14560 16540 14612
rect 17408 14603 17460 14612
rect 12256 14535 12308 14544
rect 10692 14467 10744 14476
rect 10692 14433 10701 14467
rect 10701 14433 10735 14467
rect 10735 14433 10744 14467
rect 10692 14424 10744 14433
rect 10048 14356 10100 14408
rect 2136 14288 2188 14340
rect 5540 14288 5592 14340
rect 8668 14288 8720 14340
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 12256 14501 12265 14535
rect 12265 14501 12299 14535
rect 12299 14501 12308 14535
rect 12256 14492 12308 14501
rect 12808 14492 12860 14544
rect 15936 14535 15988 14544
rect 15936 14501 15945 14535
rect 15945 14501 15979 14535
rect 15979 14501 15988 14535
rect 15936 14492 15988 14501
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 21180 14560 21232 14612
rect 22652 14603 22704 14612
rect 22652 14569 22661 14603
rect 22661 14569 22695 14603
rect 22695 14569 22704 14603
rect 22652 14560 22704 14569
rect 23756 14603 23808 14612
rect 23756 14569 23765 14603
rect 23765 14569 23799 14603
rect 23799 14569 23808 14603
rect 23756 14560 23808 14569
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 17776 14467 17828 14476
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 18972 14467 19024 14476
rect 18972 14433 18981 14467
rect 18981 14433 19015 14467
rect 19015 14433 19024 14467
rect 18972 14424 19024 14433
rect 19984 14535 20036 14544
rect 19984 14501 19993 14535
rect 19993 14501 20027 14535
rect 20027 14501 20036 14535
rect 19984 14492 20036 14501
rect 21088 14492 21140 14544
rect 20812 14424 20864 14476
rect 22192 14492 22244 14544
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 16764 14356 16816 14408
rect 19524 14356 19576 14408
rect 14096 14288 14148 14340
rect 15292 14288 15344 14340
rect 16396 14331 16448 14340
rect 16396 14297 16405 14331
rect 16405 14297 16439 14331
rect 16439 14297 16448 14331
rect 16396 14288 16448 14297
rect 20168 14288 20220 14340
rect 23480 14424 23532 14476
rect 22652 14288 22704 14340
rect 4252 14220 4304 14272
rect 10140 14220 10192 14272
rect 11244 14220 11296 14272
rect 11612 14220 11664 14272
rect 21824 14220 21876 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2872 14059 2924 14068
rect 2872 14025 2881 14059
rect 2881 14025 2915 14059
rect 2915 14025 2924 14059
rect 2872 14016 2924 14025
rect 10048 14016 10100 14068
rect 15936 14016 15988 14068
rect 16764 14059 16816 14068
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 17316 14059 17368 14068
rect 17316 14025 17325 14059
rect 17325 14025 17359 14059
rect 17359 14025 17368 14059
rect 17316 14016 17368 14025
rect 17776 14059 17828 14068
rect 17776 14025 17785 14059
rect 17785 14025 17819 14059
rect 17819 14025 17828 14059
rect 17776 14016 17828 14025
rect 21088 14016 21140 14068
rect 22652 14059 22704 14068
rect 22652 14025 22661 14059
rect 22661 14025 22695 14059
rect 22695 14025 22704 14059
rect 22652 14016 22704 14025
rect 23480 14016 23532 14068
rect 112 13948 164 14000
rect 3516 13948 3568 14000
rect 5448 13948 5500 14000
rect 11428 13991 11480 14000
rect 11428 13957 11437 13991
rect 11437 13957 11471 13991
rect 11471 13957 11480 13991
rect 11428 13948 11480 13957
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 4252 13855 4304 13864
rect 4252 13821 4261 13855
rect 4261 13821 4295 13855
rect 4295 13821 4304 13855
rect 4252 13812 4304 13821
rect 4712 13855 4764 13864
rect 4712 13821 4721 13855
rect 4721 13821 4755 13855
rect 4755 13821 4764 13855
rect 4712 13812 4764 13821
rect 1584 13787 1636 13796
rect 1584 13753 1593 13787
rect 1593 13753 1627 13787
rect 1627 13753 1636 13787
rect 1584 13744 1636 13753
rect 5080 13855 5132 13864
rect 5080 13821 5089 13855
rect 5089 13821 5123 13855
rect 5123 13821 5132 13855
rect 5080 13812 5132 13821
rect 5356 13812 5408 13864
rect 7196 13812 7248 13864
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 8116 13744 8168 13796
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 4344 13676 4396 13685
rect 6920 13719 6972 13728
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 8024 13719 8076 13728
rect 8024 13685 8033 13719
rect 8033 13685 8067 13719
rect 8067 13685 8076 13719
rect 8024 13676 8076 13685
rect 8484 13719 8536 13728
rect 8484 13685 8493 13719
rect 8493 13685 8527 13719
rect 8527 13685 8536 13719
rect 8484 13676 8536 13685
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 9956 13812 10008 13864
rect 11612 13880 11664 13932
rect 11060 13855 11112 13864
rect 11060 13821 11069 13855
rect 11069 13821 11103 13855
rect 11103 13821 11112 13855
rect 11060 13812 11112 13821
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 13084 13880 13136 13932
rect 17868 13948 17920 14000
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 15384 13880 15436 13932
rect 15936 13880 15988 13932
rect 16028 13880 16080 13932
rect 16396 13923 16448 13932
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 16396 13880 16448 13889
rect 14372 13812 14424 13864
rect 22008 13948 22060 14000
rect 23572 13948 23624 14000
rect 20076 13880 20128 13932
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 9036 13744 9088 13796
rect 9864 13676 9916 13728
rect 12256 13719 12308 13728
rect 12256 13685 12265 13719
rect 12265 13685 12299 13719
rect 12299 13685 12308 13719
rect 12256 13676 12308 13685
rect 15936 13744 15988 13796
rect 22744 13812 22796 13864
rect 23572 13812 23624 13864
rect 19892 13744 19944 13796
rect 20076 13744 20128 13796
rect 20536 13719 20588 13728
rect 20536 13685 20545 13719
rect 20545 13685 20579 13719
rect 20579 13685 20588 13719
rect 20536 13676 20588 13685
rect 20812 13676 20864 13728
rect 21824 13787 21876 13796
rect 21824 13753 21833 13787
rect 21833 13753 21867 13787
rect 21867 13753 21876 13787
rect 21824 13744 21876 13753
rect 22192 13744 22244 13796
rect 22284 13676 22336 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2320 13472 2372 13524
rect 3424 13472 3476 13524
rect 7380 13472 7432 13524
rect 9036 13515 9088 13524
rect 1676 13404 1728 13456
rect 6460 13404 6512 13456
rect 7104 13447 7156 13456
rect 7104 13413 7113 13447
rect 7113 13413 7147 13447
rect 7147 13413 7156 13447
rect 7104 13404 7156 13413
rect 9036 13481 9045 13515
rect 9045 13481 9079 13515
rect 9079 13481 9088 13515
rect 9036 13472 9088 13481
rect 9312 13472 9364 13524
rect 11428 13472 11480 13524
rect 12072 13515 12124 13524
rect 12072 13481 12081 13515
rect 12081 13481 12115 13515
rect 12115 13481 12124 13515
rect 12072 13472 12124 13481
rect 12440 13472 12492 13524
rect 12808 13472 12860 13524
rect 14372 13515 14424 13524
rect 8760 13447 8812 13456
rect 4344 13379 4396 13388
rect 4344 13345 4353 13379
rect 4353 13345 4387 13379
rect 4387 13345 4396 13379
rect 4344 13336 4396 13345
rect 4528 13379 4580 13388
rect 4528 13345 4537 13379
rect 4537 13345 4571 13379
rect 4571 13345 4580 13379
rect 4528 13336 4580 13345
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 5540 13336 5592 13388
rect 8760 13413 8769 13447
rect 8769 13413 8803 13447
rect 8803 13413 8812 13447
rect 8760 13404 8812 13413
rect 14372 13481 14381 13515
rect 14381 13481 14415 13515
rect 14415 13481 14424 13515
rect 14372 13472 14424 13481
rect 19432 13515 19484 13524
rect 19432 13481 19441 13515
rect 19441 13481 19475 13515
rect 19475 13481 19484 13515
rect 19432 13472 19484 13481
rect 3700 13268 3752 13320
rect 9956 13336 10008 13388
rect 10692 13336 10744 13388
rect 10968 13336 11020 13388
rect 13820 13404 13872 13456
rect 13912 13404 13964 13456
rect 18144 13447 18196 13456
rect 18144 13413 18153 13447
rect 18153 13413 18187 13447
rect 18187 13413 18196 13447
rect 18144 13404 18196 13413
rect 21456 13447 21508 13456
rect 21456 13413 21465 13447
rect 21465 13413 21499 13447
rect 21499 13413 21508 13447
rect 21456 13404 21508 13413
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 12256 13379 12308 13388
rect 9404 13268 9456 13320
rect 11520 13268 11572 13320
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 5356 13132 5408 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 7012 13200 7064 13252
rect 6920 13132 6972 13184
rect 7196 13132 7248 13184
rect 7748 13132 7800 13184
rect 9220 13132 9272 13184
rect 11060 13200 11112 13252
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 15384 13379 15436 13388
rect 15384 13345 15393 13379
rect 15393 13345 15427 13379
rect 15427 13345 15436 13379
rect 15384 13336 15436 13345
rect 16856 13379 16908 13388
rect 16856 13345 16865 13379
rect 16865 13345 16899 13379
rect 16899 13345 16908 13379
rect 16856 13336 16908 13345
rect 18696 13336 18748 13388
rect 19524 13379 19576 13388
rect 19524 13345 19533 13379
rect 19533 13345 19567 13379
rect 19567 13345 19576 13379
rect 19524 13336 19576 13345
rect 24676 13379 24728 13388
rect 24676 13345 24694 13379
rect 24694 13345 24728 13379
rect 24676 13336 24728 13345
rect 26240 13336 26292 13388
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 16212 13200 16264 13252
rect 22468 13268 22520 13320
rect 18420 13200 18472 13252
rect 18604 13243 18656 13252
rect 18604 13209 18613 13243
rect 18613 13209 18647 13243
rect 18647 13209 18656 13243
rect 21916 13243 21968 13252
rect 18604 13200 18656 13209
rect 21916 13209 21925 13243
rect 21925 13209 21959 13243
rect 21959 13209 21968 13243
rect 21916 13200 21968 13209
rect 17132 13132 17184 13184
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 22284 13175 22336 13184
rect 22284 13141 22293 13175
rect 22293 13141 22327 13175
rect 22327 13141 22336 13175
rect 22284 13132 22336 13141
rect 22376 13132 22428 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1584 12928 1636 12980
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 5080 12928 5132 12980
rect 6184 12928 6236 12980
rect 8668 12928 8720 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 11612 12928 11664 12980
rect 13820 12928 13872 12980
rect 14740 12928 14792 12980
rect 15384 12971 15436 12980
rect 15384 12937 15393 12971
rect 15393 12937 15427 12971
rect 15427 12937 15436 12971
rect 15384 12928 15436 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 18144 12928 18196 12980
rect 21456 12928 21508 12980
rect 24676 12928 24728 12980
rect 24860 12928 24912 12980
rect 2044 12767 2096 12776
rect 2044 12733 2053 12767
rect 2053 12733 2087 12767
rect 2087 12733 2096 12767
rect 2044 12724 2096 12733
rect 2320 12724 2372 12776
rect 4528 12792 4580 12844
rect 5724 12860 5776 12912
rect 8392 12860 8444 12912
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7104 12792 7156 12844
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5356 12724 5408 12776
rect 8760 12860 8812 12912
rect 8944 12860 8996 12912
rect 12256 12903 12308 12912
rect 12256 12869 12265 12903
rect 12265 12869 12299 12903
rect 12299 12869 12308 12903
rect 12256 12860 12308 12869
rect 13636 12860 13688 12912
rect 15936 12860 15988 12912
rect 21824 12903 21876 12912
rect 21824 12869 21833 12903
rect 21833 12869 21867 12903
rect 21867 12869 21876 12903
rect 21824 12860 21876 12869
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 12992 12792 13044 12844
rect 10692 12767 10744 12776
rect 2412 12588 2464 12640
rect 2872 12588 2924 12640
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 6276 12656 6328 12708
rect 7104 12656 7156 12708
rect 4344 12588 4396 12640
rect 4528 12588 4580 12640
rect 5724 12588 5776 12640
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 8024 12588 8076 12640
rect 10692 12733 10701 12767
rect 10701 12733 10735 12767
rect 10735 12733 10744 12767
rect 10692 12724 10744 12733
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13452 12792 13504 12844
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 9220 12656 9272 12708
rect 10048 12699 10100 12708
rect 10048 12665 10057 12699
rect 10057 12665 10091 12699
rect 10091 12665 10100 12699
rect 10048 12656 10100 12665
rect 10784 12656 10836 12708
rect 16580 12792 16632 12844
rect 20352 12792 20404 12844
rect 18604 12724 18656 12776
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 15936 12656 15988 12708
rect 16212 12699 16264 12708
rect 16212 12665 16221 12699
rect 16221 12665 16255 12699
rect 16255 12665 16264 12699
rect 16212 12656 16264 12665
rect 17408 12588 17460 12640
rect 19524 12656 19576 12708
rect 19340 12588 19392 12640
rect 22376 12792 22428 12844
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 23112 12724 23164 12776
rect 25228 12699 25280 12708
rect 25228 12665 25237 12699
rect 25237 12665 25271 12699
rect 25271 12665 25280 12699
rect 25228 12656 25280 12665
rect 22652 12588 22704 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 112 12384 164 12436
rect 1676 12359 1728 12368
rect 1676 12325 1685 12359
rect 1685 12325 1719 12359
rect 1719 12325 1728 12359
rect 1676 12316 1728 12325
rect 2044 12359 2096 12368
rect 2044 12325 2053 12359
rect 2053 12325 2087 12359
rect 2087 12325 2096 12359
rect 2044 12316 2096 12325
rect 2504 12359 2556 12368
rect 2504 12325 2513 12359
rect 2513 12325 2547 12359
rect 2547 12325 2556 12359
rect 2504 12316 2556 12325
rect 3792 12384 3844 12436
rect 12440 12427 12492 12436
rect 7288 12316 7340 12368
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 12992 12384 13044 12436
rect 13176 12384 13228 12436
rect 15936 12384 15988 12436
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 18604 12427 18656 12436
rect 18604 12393 18613 12427
rect 18613 12393 18647 12427
rect 18647 12393 18656 12427
rect 18604 12384 18656 12393
rect 10140 12316 10192 12368
rect 11336 12359 11388 12368
rect 11336 12325 11345 12359
rect 11345 12325 11379 12359
rect 11379 12325 11388 12359
rect 11336 12316 11388 12325
rect 11428 12359 11480 12368
rect 11428 12325 11437 12359
rect 11437 12325 11471 12359
rect 11471 12325 11480 12359
rect 11428 12316 11480 12325
rect 3516 12248 3568 12300
rect 5724 12291 5776 12300
rect 2964 12155 3016 12164
rect 2964 12121 2973 12155
rect 2973 12121 3007 12155
rect 3007 12121 3016 12155
rect 2964 12112 3016 12121
rect 4344 12180 4396 12232
rect 5724 12257 5733 12291
rect 5733 12257 5767 12291
rect 5767 12257 5776 12291
rect 5724 12248 5776 12257
rect 6000 12248 6052 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 6920 12248 6972 12300
rect 9220 12248 9272 12300
rect 10968 12291 11020 12300
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 14464 12316 14516 12368
rect 14740 12316 14792 12368
rect 21640 12384 21692 12436
rect 22376 12384 22428 12436
rect 21364 12359 21416 12368
rect 21364 12325 21373 12359
rect 21373 12325 21407 12359
rect 21407 12325 21416 12359
rect 21364 12316 21416 12325
rect 21916 12359 21968 12368
rect 21916 12325 21925 12359
rect 21925 12325 21959 12359
rect 21959 12325 21968 12359
rect 21916 12316 21968 12325
rect 22928 12359 22980 12368
rect 22928 12325 22937 12359
rect 22937 12325 22971 12359
rect 22971 12325 22980 12359
rect 22928 12316 22980 12325
rect 24216 12316 24268 12368
rect 6092 12180 6144 12232
rect 10140 12223 10192 12232
rect 3332 12112 3384 12164
rect 1400 12044 1452 12096
rect 8208 12112 8260 12164
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 12808 12180 12860 12232
rect 17592 12248 17644 12300
rect 18972 12291 19024 12300
rect 18972 12257 18981 12291
rect 18981 12257 19015 12291
rect 19015 12257 19024 12291
rect 18972 12248 19024 12257
rect 19432 12248 19484 12300
rect 16488 12180 16540 12232
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 21088 12180 21140 12232
rect 22836 12223 22888 12232
rect 10968 12112 11020 12164
rect 12716 12112 12768 12164
rect 13820 12112 13872 12164
rect 22836 12189 22845 12223
rect 22845 12189 22879 12223
rect 22879 12189 22888 12223
rect 22836 12180 22888 12189
rect 22192 12112 22244 12164
rect 24032 12180 24084 12232
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 8852 12087 8904 12096
rect 8852 12053 8861 12087
rect 8861 12053 8895 12087
rect 8895 12053 8904 12087
rect 8852 12044 8904 12053
rect 15660 12044 15712 12096
rect 16672 12044 16724 12096
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 20076 12087 20128 12096
rect 20076 12053 20085 12087
rect 20085 12053 20119 12087
rect 20119 12053 20128 12087
rect 20076 12044 20128 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2504 11840 2556 11892
rect 4620 11840 4672 11892
rect 5540 11840 5592 11892
rect 8944 11840 8996 11892
rect 10784 11840 10836 11892
rect 11336 11840 11388 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 6276 11772 6328 11824
rect 13176 11772 13228 11824
rect 7012 11704 7064 11756
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 9680 11704 9732 11756
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 8944 11679 8996 11688
rect 2688 11611 2740 11620
rect 2688 11577 2697 11611
rect 2697 11577 2731 11611
rect 2731 11577 2740 11611
rect 2688 11568 2740 11577
rect 112 11500 164 11552
rect 5448 11500 5500 11552
rect 6092 11500 6144 11552
rect 8668 11500 8720 11552
rect 8944 11645 8953 11679
rect 8953 11645 8987 11679
rect 8987 11645 8996 11679
rect 8944 11636 8996 11645
rect 10876 11636 10928 11688
rect 15844 11772 15896 11824
rect 20536 11840 20588 11892
rect 21364 11840 21416 11892
rect 22836 11840 22888 11892
rect 23388 11883 23440 11892
rect 23388 11849 23397 11883
rect 23397 11849 23431 11883
rect 23431 11849 23440 11883
rect 23388 11840 23440 11849
rect 24032 11883 24084 11892
rect 24032 11849 24041 11883
rect 24041 11849 24075 11883
rect 24075 11849 24084 11883
rect 24032 11840 24084 11849
rect 24216 11840 24268 11892
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 18236 11772 18288 11824
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 15936 11704 15988 11756
rect 16580 11704 16632 11756
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 9680 11568 9732 11620
rect 9220 11500 9272 11552
rect 11428 11568 11480 11620
rect 13452 11568 13504 11620
rect 13544 11568 13596 11620
rect 19340 11636 19392 11688
rect 12716 11500 12768 11552
rect 14740 11500 14792 11552
rect 16028 11568 16080 11620
rect 17408 11568 17460 11620
rect 18236 11611 18288 11620
rect 18236 11577 18245 11611
rect 18245 11577 18279 11611
rect 18279 11577 18288 11611
rect 18236 11568 18288 11577
rect 22376 11772 22428 11824
rect 22192 11704 22244 11756
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 22928 11636 22980 11688
rect 24584 11679 24636 11688
rect 24584 11645 24593 11679
rect 24593 11645 24627 11679
rect 24627 11645 24636 11679
rect 24584 11636 24636 11645
rect 22836 11568 22888 11620
rect 24032 11568 24084 11620
rect 15660 11500 15712 11552
rect 18420 11500 18472 11552
rect 18972 11500 19024 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 4160 11339 4212 11348
rect 4160 11305 4169 11339
rect 4169 11305 4203 11339
rect 4203 11305 4212 11339
rect 4160 11296 4212 11305
rect 1676 11228 1728 11280
rect 2412 11228 2464 11280
rect 3884 11228 3936 11280
rect 6000 11296 6052 11348
rect 6184 11339 6236 11348
rect 6184 11305 6193 11339
rect 6193 11305 6227 11339
rect 6227 11305 6236 11339
rect 6184 11296 6236 11305
rect 9312 11296 9364 11348
rect 9680 11296 9732 11348
rect 6368 11271 6420 11280
rect 6368 11237 6377 11271
rect 6377 11237 6411 11271
rect 6411 11237 6420 11271
rect 6368 11228 6420 11237
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 4988 11203 5040 11212
rect 4988 11169 4997 11203
rect 4997 11169 5031 11203
rect 5031 11169 5040 11203
rect 4988 11160 5040 11169
rect 5540 11160 5592 11212
rect 7104 11228 7156 11280
rect 8484 11228 8536 11280
rect 8668 11271 8720 11280
rect 8668 11237 8677 11271
rect 8677 11237 8711 11271
rect 8711 11237 8720 11271
rect 8668 11228 8720 11237
rect 9864 11228 9916 11280
rect 10692 11296 10744 11348
rect 10876 11339 10928 11348
rect 10876 11305 10885 11339
rect 10885 11305 10919 11339
rect 10919 11305 10928 11339
rect 10876 11296 10928 11305
rect 10968 11296 11020 11348
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 17040 11296 17092 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 19984 11296 20036 11348
rect 21088 11339 21140 11348
rect 21088 11305 21097 11339
rect 21097 11305 21131 11339
rect 21131 11305 21140 11339
rect 21088 11296 21140 11305
rect 22284 11296 22336 11348
rect 24584 11296 24636 11348
rect 11612 11271 11664 11280
rect 11612 11237 11621 11271
rect 11621 11237 11655 11271
rect 11655 11237 11664 11271
rect 11612 11228 11664 11237
rect 15660 11271 15712 11280
rect 15660 11237 15669 11271
rect 15669 11237 15703 11271
rect 15703 11237 15712 11271
rect 15660 11228 15712 11237
rect 16212 11271 16264 11280
rect 16212 11237 16221 11271
rect 16221 11237 16255 11271
rect 16255 11237 16264 11271
rect 16212 11228 16264 11237
rect 20076 11228 20128 11280
rect 22376 11228 22428 11280
rect 8024 11203 8076 11212
rect 2780 11092 2832 11144
rect 2504 11024 2556 11076
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 1952 10999 2004 11008
rect 1952 10965 1961 10999
rect 1961 10965 1995 10999
rect 1995 10965 2004 10999
rect 1952 10956 2004 10965
rect 3332 10956 3384 11008
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 7472 10956 7524 10965
rect 7564 10956 7616 11008
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 16672 11160 16724 11212
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 19064 11203 19116 11212
rect 19064 11169 19073 11203
rect 19073 11169 19107 11203
rect 19107 11169 19116 11203
rect 19064 11160 19116 11169
rect 19432 11160 19484 11212
rect 21088 11160 21140 11212
rect 23020 11160 23072 11212
rect 23572 11160 23624 11212
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 12992 11135 13044 11144
rect 10140 11024 10192 11076
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 11980 11024 12032 11076
rect 22284 11024 22336 11076
rect 22468 11092 22520 11144
rect 9220 10956 9272 11008
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 16488 10956 16540 11008
rect 17316 10956 17368 11008
rect 19616 10956 19668 11008
rect 22192 10956 22244 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2412 10795 2464 10804
rect 2412 10761 2421 10795
rect 2421 10761 2455 10795
rect 2455 10761 2464 10795
rect 2412 10752 2464 10761
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 4160 10752 4212 10804
rect 4344 10752 4396 10804
rect 9772 10752 9824 10804
rect 10048 10752 10100 10804
rect 10692 10752 10744 10804
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 15568 10752 15620 10804
rect 21088 10752 21140 10804
rect 22008 10795 22060 10804
rect 22008 10761 22017 10795
rect 22017 10761 22051 10795
rect 22051 10761 22060 10795
rect 22008 10752 22060 10761
rect 22836 10752 22888 10804
rect 23388 10752 23440 10804
rect 2964 10684 3016 10736
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1952 10616 2004 10668
rect 5540 10684 5592 10736
rect 6276 10684 6328 10736
rect 6184 10616 6236 10668
rect 12716 10684 12768 10736
rect 15660 10684 15712 10736
rect 22376 10727 22428 10736
rect 22376 10693 22385 10727
rect 22385 10693 22419 10727
rect 22419 10693 22428 10727
rect 22376 10684 22428 10693
rect 10140 10616 10192 10668
rect 10968 10659 11020 10668
rect 10968 10625 10977 10659
rect 10977 10625 11011 10659
rect 11011 10625 11020 10659
rect 10968 10616 11020 10625
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 6828 10591 6880 10600
rect 1676 10480 1728 10532
rect 3148 10523 3200 10532
rect 1768 10412 1820 10464
rect 3148 10489 3157 10523
rect 3157 10489 3191 10523
rect 3191 10489 3200 10523
rect 3148 10480 3200 10489
rect 4988 10455 5040 10464
rect 4988 10421 4997 10455
rect 4997 10421 5031 10455
rect 5031 10421 5040 10455
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 7472 10548 7524 10600
rect 6184 10455 6236 10464
rect 4988 10412 5040 10421
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 7564 10412 7616 10464
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9312 10548 9364 10600
rect 13820 10591 13872 10600
rect 13820 10557 13829 10591
rect 13829 10557 13863 10591
rect 13863 10557 13872 10591
rect 13820 10548 13872 10557
rect 14096 10548 14148 10600
rect 15476 10616 15528 10668
rect 23020 10616 23072 10668
rect 23572 10616 23624 10668
rect 15568 10591 15620 10600
rect 15568 10557 15577 10591
rect 15577 10557 15611 10591
rect 15611 10557 15620 10591
rect 15568 10548 15620 10557
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16856 10548 16908 10600
rect 18236 10591 18288 10600
rect 9680 10523 9732 10532
rect 9680 10489 9689 10523
rect 9689 10489 9723 10523
rect 9723 10489 9732 10523
rect 9680 10480 9732 10489
rect 10692 10523 10744 10532
rect 10692 10489 10701 10523
rect 10701 10489 10735 10523
rect 10735 10489 10744 10523
rect 12532 10523 12584 10532
rect 10692 10480 10744 10489
rect 12532 10489 12541 10523
rect 12541 10489 12575 10523
rect 12575 10489 12584 10523
rect 12532 10480 12584 10489
rect 11612 10455 11664 10464
rect 11612 10421 11621 10455
rect 11621 10421 11655 10455
rect 11655 10421 11664 10455
rect 11612 10412 11664 10421
rect 12992 10480 13044 10532
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 22008 10548 22060 10600
rect 23112 10591 23164 10600
rect 23112 10557 23121 10591
rect 23121 10557 23155 10591
rect 23155 10557 23164 10591
rect 23112 10548 23164 10557
rect 24124 10548 24176 10600
rect 12716 10412 12768 10464
rect 15936 10412 15988 10464
rect 16488 10455 16540 10464
rect 16488 10421 16497 10455
rect 16497 10421 16531 10455
rect 16531 10421 16540 10455
rect 16488 10412 16540 10421
rect 16672 10412 16724 10464
rect 17868 10412 17920 10464
rect 18604 10480 18656 10532
rect 19064 10480 19116 10532
rect 19340 10480 19392 10532
rect 19616 10523 19668 10532
rect 19616 10489 19625 10523
rect 19625 10489 19659 10523
rect 19659 10489 19668 10523
rect 19616 10480 19668 10489
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 20444 10455 20496 10464
rect 20444 10421 20453 10455
rect 20453 10421 20487 10455
rect 20487 10421 20496 10455
rect 20444 10412 20496 10421
rect 21180 10523 21232 10532
rect 21180 10489 21189 10523
rect 21189 10489 21223 10523
rect 21223 10489 21232 10523
rect 21732 10523 21784 10532
rect 21180 10480 21232 10489
rect 21732 10489 21741 10523
rect 21741 10489 21775 10523
rect 21775 10489 21784 10523
rect 21732 10480 21784 10489
rect 21824 10480 21876 10532
rect 21548 10412 21600 10464
rect 24216 10455 24268 10464
rect 24216 10421 24225 10455
rect 24225 10421 24259 10455
rect 24259 10421 24268 10455
rect 24216 10412 24268 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3148 10208 3200 10260
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 4528 10208 4580 10260
rect 6000 10208 6052 10260
rect 2412 10140 2464 10192
rect 6184 10140 6236 10192
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6552 10072 6604 10124
rect 6828 10208 6880 10260
rect 8024 10208 8076 10260
rect 8484 10208 8536 10260
rect 9680 10208 9732 10260
rect 9220 10140 9272 10192
rect 10784 10183 10836 10192
rect 10784 10149 10793 10183
rect 10793 10149 10827 10183
rect 10827 10149 10836 10183
rect 10784 10140 10836 10149
rect 11520 10208 11572 10260
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 12164 10208 12216 10260
rect 14464 10208 14516 10260
rect 15660 10208 15712 10260
rect 17592 10208 17644 10260
rect 19524 10208 19576 10260
rect 22652 10208 22704 10260
rect 17132 10183 17184 10192
rect 17132 10149 17141 10183
rect 17141 10149 17175 10183
rect 17175 10149 17184 10183
rect 17132 10140 17184 10149
rect 17224 10183 17276 10192
rect 17224 10149 17233 10183
rect 17233 10149 17267 10183
rect 17267 10149 17276 10183
rect 17224 10140 17276 10149
rect 19248 10140 19300 10192
rect 19432 10140 19484 10192
rect 20904 10140 20956 10192
rect 22928 10208 22980 10260
rect 8116 10115 8168 10124
rect 2320 10004 2372 10056
rect 2688 9868 2740 9920
rect 3424 9911 3476 9920
rect 3424 9877 3433 9911
rect 3433 9877 3467 9911
rect 3467 9877 3476 9911
rect 3424 9868 3476 9877
rect 4344 10004 4396 10056
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 12164 10115 12216 10124
rect 12164 10081 12173 10115
rect 12173 10081 12207 10115
rect 12207 10081 12216 10115
rect 12164 10072 12216 10081
rect 12716 10115 12768 10124
rect 12716 10081 12725 10115
rect 12725 10081 12759 10115
rect 12759 10081 12768 10115
rect 12716 10072 12768 10081
rect 3976 9936 4028 9988
rect 4988 9936 5040 9988
rect 6368 9936 6420 9988
rect 7840 10004 7892 10056
rect 8668 10004 8720 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 13360 10072 13412 10124
rect 14096 10072 14148 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 18144 10115 18196 10124
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 21824 10072 21876 10124
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 19156 10004 19208 10056
rect 12992 9936 13044 9988
rect 13636 9936 13688 9988
rect 17684 9979 17736 9988
rect 17684 9945 17693 9979
rect 17693 9945 17727 9979
rect 17727 9945 17736 9979
rect 17684 9936 17736 9945
rect 19340 9936 19392 9988
rect 20720 10004 20772 10056
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 22928 9936 22980 9988
rect 23296 9936 23348 9988
rect 24768 10115 24820 10124
rect 24768 10081 24777 10115
rect 24777 10081 24811 10115
rect 24811 10081 24820 10115
rect 24768 10072 24820 10081
rect 4528 9868 4580 9920
rect 5172 9868 5224 9920
rect 9864 9868 9916 9920
rect 16304 9868 16356 9920
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 23204 9868 23256 9920
rect 24768 9868 24820 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1676 9707 1728 9716
rect 1676 9673 1685 9707
rect 1685 9673 1719 9707
rect 1719 9673 1728 9707
rect 1676 9664 1728 9673
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 2964 9707 3016 9716
rect 2964 9673 2973 9707
rect 2973 9673 3007 9707
rect 3007 9673 3016 9707
rect 2964 9664 3016 9673
rect 6184 9707 6236 9716
rect 6184 9673 6193 9707
rect 6193 9673 6227 9707
rect 6227 9673 6236 9707
rect 6184 9664 6236 9673
rect 8116 9664 8168 9716
rect 10784 9707 10836 9716
rect 10784 9673 10793 9707
rect 10793 9673 10827 9707
rect 10827 9673 10836 9707
rect 10784 9664 10836 9673
rect 12992 9664 13044 9716
rect 13452 9664 13504 9716
rect 13728 9664 13780 9716
rect 7748 9596 7800 9648
rect 10692 9596 10744 9648
rect 12808 9596 12860 9648
rect 15844 9664 15896 9716
rect 16028 9707 16080 9716
rect 16028 9673 16037 9707
rect 16037 9673 16071 9707
rect 16071 9673 16080 9707
rect 16028 9664 16080 9673
rect 19248 9664 19300 9716
rect 21640 9664 21692 9716
rect 22652 9707 22704 9716
rect 6368 9528 6420 9580
rect 1952 9460 2004 9512
rect 2596 9460 2648 9512
rect 2688 9460 2740 9512
rect 5172 9503 5224 9512
rect 1860 9392 1912 9444
rect 4436 9392 4488 9444
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 6736 9460 6788 9512
rect 8300 9528 8352 9580
rect 7564 9460 7616 9512
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 6092 9392 6144 9444
rect 6184 9392 6236 9444
rect 8944 9460 8996 9512
rect 11796 9528 11848 9580
rect 13636 9528 13688 9580
rect 12624 9460 12676 9512
rect 9864 9435 9916 9444
rect 9864 9401 9873 9435
rect 9873 9401 9907 9435
rect 9907 9401 9916 9435
rect 9864 9392 9916 9401
rect 4160 9324 4212 9376
rect 4528 9324 4580 9376
rect 5448 9324 5500 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 10692 9392 10744 9444
rect 13912 9435 13964 9444
rect 13912 9401 13921 9435
rect 13921 9401 13955 9435
rect 13955 9401 13964 9435
rect 13912 9392 13964 9401
rect 14832 9392 14884 9444
rect 9588 9324 9640 9333
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 13636 9324 13688 9376
rect 15660 9324 15712 9376
rect 17408 9596 17460 9648
rect 20444 9596 20496 9648
rect 21180 9596 21232 9648
rect 21824 9596 21876 9648
rect 22652 9673 22661 9707
rect 22661 9673 22695 9707
rect 22695 9673 22704 9707
rect 22652 9664 22704 9673
rect 24768 9664 24820 9716
rect 25780 9707 25832 9716
rect 25780 9673 25789 9707
rect 25789 9673 25823 9707
rect 25823 9673 25832 9707
rect 25780 9664 25832 9673
rect 17684 9528 17736 9580
rect 19340 9528 19392 9580
rect 21640 9528 21692 9580
rect 22744 9528 22796 9580
rect 16304 9460 16356 9512
rect 17040 9460 17092 9512
rect 17224 9460 17276 9512
rect 19524 9460 19576 9512
rect 18144 9435 18196 9444
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 17408 9324 17460 9376
rect 19248 9392 19300 9444
rect 20904 9435 20956 9444
rect 20904 9401 20913 9435
rect 20913 9401 20947 9435
rect 20947 9401 20956 9435
rect 20904 9392 20956 9401
rect 21272 9392 21324 9444
rect 21824 9392 21876 9444
rect 23296 9392 23348 9444
rect 25780 9460 25832 9512
rect 18788 9324 18840 9376
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 21456 9324 21508 9376
rect 23940 9324 23992 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1492 9120 1544 9172
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 2688 9027 2740 9036
rect 2136 8916 2188 8968
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 5080 9120 5132 9172
rect 6368 9163 6420 9172
rect 204 8848 256 8900
rect 5172 9052 5224 9104
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6552 9120 6604 9172
rect 7288 9120 7340 9172
rect 9128 9052 9180 9104
rect 9588 9052 9640 9104
rect 4252 8984 4304 9036
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 8024 8984 8076 9036
rect 3976 8916 4028 8968
rect 7472 8916 7524 8968
rect 9312 8984 9364 9036
rect 11796 8984 11848 9036
rect 12716 9120 12768 9172
rect 13268 9120 13320 9172
rect 13452 9120 13504 9172
rect 17132 9120 17184 9172
rect 18788 9163 18840 9172
rect 18788 9129 18797 9163
rect 18797 9129 18831 9163
rect 18831 9129 18840 9163
rect 18788 9120 18840 9129
rect 19156 9163 19208 9172
rect 19156 9129 19165 9163
rect 19165 9129 19199 9163
rect 19199 9129 19208 9163
rect 19156 9120 19208 9129
rect 20536 9120 20588 9172
rect 16028 9052 16080 9104
rect 17776 9052 17828 9104
rect 23296 9120 23348 9172
rect 21088 9095 21140 9104
rect 21088 9061 21097 9095
rect 21097 9061 21131 9095
rect 21131 9061 21140 9095
rect 21088 9052 21140 9061
rect 21272 9052 21324 9104
rect 22652 9095 22704 9104
rect 22652 9061 22661 9095
rect 22661 9061 22695 9095
rect 22695 9061 22704 9095
rect 22652 9052 22704 9061
rect 23572 9052 23624 9104
rect 13912 9027 13964 9036
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 10784 8916 10836 8968
rect 11244 8916 11296 8968
rect 13912 8993 13921 9027
rect 13921 8993 13955 9027
rect 13955 8993 13964 9027
rect 13912 8984 13964 8993
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 16856 8984 16908 9036
rect 18512 8984 18564 9036
rect 20076 8984 20128 9036
rect 25136 8984 25188 9036
rect 12808 8916 12860 8968
rect 20628 8916 20680 8968
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 21732 8916 21784 8968
rect 22928 8916 22980 8968
rect 9864 8848 9916 8900
rect 19524 8848 19576 8900
rect 21456 8848 21508 8900
rect 21548 8848 21600 8900
rect 2780 8780 2832 8832
rect 3792 8780 3844 8832
rect 6000 8780 6052 8832
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 17224 8780 17276 8832
rect 19432 8780 19484 8832
rect 20720 8780 20772 8832
rect 20996 8780 21048 8832
rect 21272 8780 21324 8832
rect 24032 8780 24084 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2688 8576 2740 8628
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 3976 8576 4028 8628
rect 112 8508 164 8560
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 5448 8576 5500 8628
rect 5540 8576 5592 8628
rect 6000 8576 6052 8628
rect 7840 8576 7892 8628
rect 8668 8576 8720 8628
rect 9772 8576 9824 8628
rect 10784 8619 10836 8628
rect 10784 8585 10793 8619
rect 10793 8585 10827 8619
rect 10827 8585 10836 8619
rect 17776 8619 17828 8628
rect 10784 8576 10836 8585
rect 5356 8508 5408 8560
rect 8116 8508 8168 8560
rect 11244 8551 11296 8560
rect 11244 8517 11253 8551
rect 11253 8517 11287 8551
rect 11287 8517 11296 8551
rect 11244 8508 11296 8517
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 3792 8372 3844 8424
rect 4528 8372 4580 8424
rect 7288 8440 7340 8492
rect 8760 8440 8812 8492
rect 9404 8440 9456 8492
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 21088 8619 21140 8628
rect 21088 8585 21097 8619
rect 21097 8585 21131 8619
rect 21131 8585 21140 8619
rect 21088 8576 21140 8585
rect 22652 8619 22704 8628
rect 22652 8585 22661 8619
rect 22661 8585 22695 8619
rect 22695 8585 22704 8619
rect 22652 8576 22704 8585
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 13268 8508 13320 8560
rect 16028 8551 16080 8560
rect 16028 8517 16037 8551
rect 16037 8517 16071 8551
rect 16071 8517 16080 8551
rect 16028 8508 16080 8517
rect 17500 8551 17552 8560
rect 17500 8517 17509 8551
rect 17509 8517 17543 8551
rect 17543 8517 17552 8551
rect 17500 8508 17552 8517
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 14832 8440 14884 8492
rect 15660 8440 15712 8492
rect 5080 8415 5132 8424
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 5448 8415 5500 8424
rect 5448 8381 5457 8415
rect 5457 8381 5491 8415
rect 5491 8381 5500 8415
rect 5448 8372 5500 8381
rect 7564 8372 7616 8424
rect 9496 8372 9548 8424
rect 7472 8304 7524 8356
rect 4160 8279 4212 8288
rect 4160 8245 4169 8279
rect 4169 8245 4203 8279
rect 4203 8245 4212 8279
rect 4160 8236 4212 8245
rect 7380 8236 7432 8288
rect 8668 8304 8720 8356
rect 11428 8372 11480 8424
rect 20076 8508 20128 8560
rect 23020 8508 23072 8560
rect 19984 8440 20036 8492
rect 20996 8440 21048 8492
rect 21272 8483 21324 8492
rect 21272 8449 21281 8483
rect 21281 8449 21315 8483
rect 21315 8449 21324 8483
rect 21640 8483 21692 8492
rect 21272 8440 21324 8449
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 18328 8415 18380 8424
rect 18328 8381 18337 8415
rect 18337 8381 18371 8415
rect 18371 8381 18380 8415
rect 18328 8372 18380 8381
rect 18604 8415 18656 8424
rect 18604 8381 18613 8415
rect 18613 8381 18647 8415
rect 18647 8381 18656 8415
rect 18604 8372 18656 8381
rect 19432 8372 19484 8424
rect 9772 8304 9824 8356
rect 12164 8347 12216 8356
rect 12164 8313 12173 8347
rect 12173 8313 12207 8347
rect 12207 8313 12216 8347
rect 12164 8304 12216 8313
rect 13268 8304 13320 8356
rect 13636 8304 13688 8356
rect 14740 8347 14792 8356
rect 14740 8313 14749 8347
rect 14749 8313 14783 8347
rect 14783 8313 14792 8347
rect 14740 8304 14792 8313
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 9588 8236 9640 8288
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 17040 8304 17092 8356
rect 15476 8236 15528 8288
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8032 1452 8084
rect 2136 8032 2188 8084
rect 4252 8032 4304 8084
rect 4528 8032 4580 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8024 8032 8076 8084
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 9496 8032 9548 8084
rect 12808 8075 12860 8084
rect 2504 7964 2556 8016
rect 1768 7896 1820 7948
rect 5080 7964 5132 8016
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 6276 7964 6328 8016
rect 8208 8007 8260 8016
rect 8208 7973 8217 8007
rect 8217 7973 8251 8007
rect 8251 7973 8260 8007
rect 8208 7964 8260 7973
rect 8760 7964 8812 8016
rect 10140 7964 10192 8016
rect 11428 8007 11480 8016
rect 11428 7973 11437 8007
rect 11437 7973 11471 8007
rect 11471 7973 11480 8007
rect 11428 7964 11480 7973
rect 12808 8041 12817 8075
rect 12817 8041 12851 8075
rect 12851 8041 12860 8075
rect 12808 8032 12860 8041
rect 14740 8032 14792 8084
rect 16120 8032 16172 8084
rect 12900 7964 12952 8016
rect 18144 8032 18196 8084
rect 18328 8032 18380 8084
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 20628 8075 20680 8084
rect 20628 8041 20637 8075
rect 20637 8041 20671 8075
rect 20671 8041 20680 8075
rect 20628 8032 20680 8041
rect 6184 7896 6236 7948
rect 6644 7896 6696 7948
rect 12256 7896 12308 7948
rect 13176 7896 13228 7948
rect 17408 7964 17460 8016
rect 18880 8007 18932 8016
rect 18880 7973 18889 8007
rect 18889 7973 18923 8007
rect 18923 7973 18932 8007
rect 18880 7964 18932 7973
rect 21088 8007 21140 8016
rect 21088 7973 21097 8007
rect 21097 7973 21131 8007
rect 21131 7973 21140 8007
rect 21088 7964 21140 7973
rect 21640 8007 21692 8016
rect 21640 7973 21649 8007
rect 21649 7973 21683 8007
rect 21683 7973 21692 8007
rect 21640 7964 21692 7973
rect 15936 7896 15988 7948
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 2596 7828 2648 7880
rect 4436 7828 4488 7880
rect 4988 7828 5040 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8944 7828 8996 7880
rect 9864 7828 9916 7880
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 10784 7828 10836 7880
rect 940 7760 992 7812
rect 1676 7760 1728 7812
rect 4712 7760 4764 7812
rect 5080 7760 5132 7812
rect 9496 7760 9548 7812
rect 10692 7760 10744 7812
rect 12992 7760 13044 7812
rect 23020 7896 23072 7948
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 18512 7828 18564 7880
rect 16120 7760 16172 7812
rect 21272 7828 21324 7880
rect 6920 7692 6972 7744
rect 14556 7735 14608 7744
rect 14556 7701 14565 7735
rect 14565 7701 14599 7735
rect 14599 7701 14608 7735
rect 14556 7692 14608 7701
rect 15752 7692 15804 7744
rect 16672 7692 16724 7744
rect 19892 7735 19944 7744
rect 19892 7701 19901 7735
rect 19901 7701 19935 7735
rect 19935 7701 19944 7735
rect 19892 7692 19944 7701
rect 21548 7692 21600 7744
rect 21916 7735 21968 7744
rect 21916 7701 21925 7735
rect 21925 7701 21959 7735
rect 21959 7701 21968 7735
rect 21916 7692 21968 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2504 7488 2556 7540
rect 4528 7488 4580 7540
rect 6644 7531 6696 7540
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 8208 7488 8260 7540
rect 8944 7531 8996 7540
rect 8944 7497 8953 7531
rect 8953 7497 8987 7531
rect 8987 7497 8996 7531
rect 8944 7488 8996 7497
rect 11428 7488 11480 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 12900 7488 12952 7540
rect 1676 7420 1728 7472
rect 8116 7420 8168 7472
rect 10048 7463 10100 7472
rect 10048 7429 10057 7463
rect 10057 7429 10091 7463
rect 10091 7429 10100 7463
rect 10048 7420 10100 7429
rect 3516 7352 3568 7404
rect 4160 7352 4212 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 6552 7352 6604 7404
rect 14372 7488 14424 7540
rect 14832 7488 14884 7540
rect 15844 7488 15896 7540
rect 17408 7531 17460 7540
rect 15936 7420 15988 7472
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 14556 7395 14608 7404
rect 1584 7284 1636 7336
rect 6184 7284 6236 7336
rect 11888 7284 11940 7336
rect 2320 7216 2372 7268
rect 5632 7216 5684 7268
rect 6920 7259 6972 7268
rect 6920 7225 6929 7259
rect 6929 7225 6963 7259
rect 6963 7225 6972 7259
rect 6920 7216 6972 7225
rect 7012 7259 7064 7268
rect 7012 7225 7021 7259
rect 7021 7225 7055 7259
rect 7055 7225 7064 7259
rect 9496 7259 9548 7268
rect 7012 7216 7064 7225
rect 9496 7225 9505 7259
rect 9505 7225 9539 7259
rect 9539 7225 9548 7259
rect 9496 7216 9548 7225
rect 9588 7259 9640 7268
rect 9588 7225 9597 7259
rect 9597 7225 9631 7259
rect 9631 7225 9640 7259
rect 9588 7216 9640 7225
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 4252 7148 4304 7200
rect 5540 7148 5592 7200
rect 8668 7148 8720 7200
rect 10140 7148 10192 7200
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 13084 7259 13136 7268
rect 13084 7225 13093 7259
rect 13093 7225 13127 7259
rect 13127 7225 13136 7259
rect 13084 7216 13136 7225
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 13912 7284 13964 7336
rect 17408 7497 17417 7531
rect 17417 7497 17451 7531
rect 17451 7497 17460 7531
rect 17408 7488 17460 7497
rect 19984 7488 20036 7540
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 23388 7488 23440 7540
rect 21088 7420 21140 7472
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 15660 7216 15712 7268
rect 16120 7216 16172 7268
rect 20720 7284 20772 7336
rect 22836 7284 22888 7336
rect 17132 7259 17184 7268
rect 17132 7225 17141 7259
rect 17141 7225 17175 7259
rect 17175 7225 17184 7259
rect 17132 7216 17184 7225
rect 17776 7191 17828 7200
rect 17776 7157 17785 7191
rect 17785 7157 17819 7191
rect 17819 7157 17828 7191
rect 19156 7216 19208 7268
rect 19984 7259 20036 7268
rect 19984 7225 19993 7259
rect 19993 7225 20027 7259
rect 20027 7225 20036 7259
rect 19984 7216 20036 7225
rect 20076 7259 20128 7268
rect 20076 7225 20085 7259
rect 20085 7225 20119 7259
rect 20119 7225 20128 7259
rect 20076 7216 20128 7225
rect 21732 7216 21784 7268
rect 17776 7148 17828 7157
rect 18880 7148 18932 7200
rect 19524 7148 19576 7200
rect 21272 7191 21324 7200
rect 21272 7157 21281 7191
rect 21281 7157 21315 7191
rect 21315 7157 21324 7191
rect 21272 7148 21324 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1768 6944 1820 6996
rect 3516 6987 3568 6996
rect 3516 6953 3525 6987
rect 3525 6953 3559 6987
rect 3559 6953 3568 6987
rect 3516 6944 3568 6953
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 5356 6944 5408 6996
rect 5632 6944 5684 6996
rect 2412 6919 2464 6928
rect 2412 6885 2421 6919
rect 2421 6885 2455 6919
rect 2455 6885 2464 6919
rect 2412 6876 2464 6885
rect 4252 6919 4304 6928
rect 1584 6808 1636 6860
rect 2964 6808 3016 6860
rect 4252 6885 4261 6919
rect 4261 6885 4295 6919
rect 4295 6885 4304 6919
rect 4252 6876 4304 6885
rect 6000 6919 6052 6928
rect 6000 6885 6009 6919
rect 6009 6885 6043 6919
rect 6043 6885 6052 6919
rect 6000 6876 6052 6885
rect 6552 6919 6604 6928
rect 6552 6885 6561 6919
rect 6561 6885 6595 6919
rect 6595 6885 6604 6919
rect 6552 6876 6604 6885
rect 6920 6944 6972 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 11244 6944 11296 6996
rect 12992 6987 13044 6996
rect 7380 6876 7432 6928
rect 10140 6876 10192 6928
rect 11428 6876 11480 6928
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 9128 6808 9180 6860
rect 10324 6851 10376 6860
rect 10324 6817 10333 6851
rect 10333 6817 10367 6851
rect 10367 6817 10376 6851
rect 10324 6808 10376 6817
rect 12992 6953 13001 6987
rect 13001 6953 13035 6987
rect 13035 6953 13044 6987
rect 12992 6944 13044 6953
rect 13084 6944 13136 6996
rect 17224 6944 17276 6996
rect 18144 6987 18196 6996
rect 18144 6953 18153 6987
rect 18153 6953 18187 6987
rect 18187 6953 18196 6987
rect 18144 6944 18196 6953
rect 18512 6987 18564 6996
rect 18512 6953 18521 6987
rect 18521 6953 18555 6987
rect 18555 6953 18564 6987
rect 18512 6944 18564 6953
rect 19524 6944 19576 6996
rect 20076 6944 20128 6996
rect 13912 6876 13964 6928
rect 14372 6919 14424 6928
rect 14372 6885 14381 6919
rect 14381 6885 14415 6919
rect 14415 6885 14424 6919
rect 14372 6876 14424 6885
rect 16120 6919 16172 6928
rect 16120 6885 16129 6919
rect 16129 6885 16163 6919
rect 16163 6885 16172 6919
rect 16120 6876 16172 6885
rect 16672 6876 16724 6928
rect 19248 6919 19300 6928
rect 19248 6885 19257 6919
rect 19257 6885 19291 6919
rect 19291 6885 19300 6919
rect 19248 6876 19300 6885
rect 21088 6919 21140 6928
rect 21088 6885 21097 6919
rect 21097 6885 21131 6919
rect 21131 6885 21140 6919
rect 21088 6876 21140 6885
rect 21732 6876 21784 6928
rect 15568 6851 15620 6860
rect 2596 6740 2648 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 6644 6740 6696 6792
rect 7932 6740 7984 6792
rect 9588 6740 9640 6792
rect 15568 6817 15577 6851
rect 15577 6817 15611 6851
rect 15611 6817 15620 6851
rect 15568 6808 15620 6817
rect 16304 6808 16356 6860
rect 18604 6808 18656 6860
rect 11612 6740 11664 6792
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 4344 6672 4396 6724
rect 6552 6672 6604 6724
rect 13636 6672 13688 6724
rect 5540 6604 5592 6656
rect 7012 6604 7064 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 16764 6604 16816 6656
rect 17776 6604 17828 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 19156 6740 19208 6792
rect 20720 6740 20772 6792
rect 21456 6672 21508 6724
rect 18788 6604 18840 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1676 6400 1728 6452
rect 2228 6400 2280 6452
rect 2596 6400 2648 6452
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 3424 6400 3476 6452
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 6184 6400 6236 6452
rect 7288 6400 7340 6452
rect 8668 6400 8720 6452
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 11612 6400 11664 6452
rect 12164 6443 12216 6452
rect 7380 6375 7432 6384
rect 7380 6341 7389 6375
rect 7389 6341 7423 6375
rect 7423 6341 7432 6375
rect 7380 6332 7432 6341
rect 7840 6332 7892 6384
rect 9036 6332 9088 6384
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 13084 6400 13136 6452
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 16120 6400 16172 6452
rect 16304 6400 16356 6452
rect 18972 6400 19024 6452
rect 22836 6400 22888 6452
rect 15660 6332 15712 6384
rect 19248 6332 19300 6384
rect 21088 6332 21140 6384
rect 2504 6264 2556 6316
rect 6000 6264 6052 6316
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 8944 6264 8996 6316
rect 3976 6196 4028 6248
rect 5540 6196 5592 6248
rect 7288 6239 7340 6248
rect 7288 6205 7297 6239
rect 7297 6205 7331 6239
rect 7331 6205 7340 6239
rect 7288 6196 7340 6205
rect 3976 6103 4028 6112
rect 3976 6069 3985 6103
rect 3985 6069 4019 6103
rect 4019 6069 4028 6103
rect 3976 6060 4028 6069
rect 7288 6060 7340 6112
rect 9312 6196 9364 6248
rect 11980 6264 12032 6316
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 14372 6264 14424 6316
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 16212 6264 16264 6316
rect 18788 6307 18840 6316
rect 18788 6273 18797 6307
rect 18797 6273 18831 6307
rect 18831 6273 18840 6307
rect 18788 6264 18840 6273
rect 10876 6196 10928 6248
rect 11244 6239 11296 6248
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 12164 6196 12216 6248
rect 11152 6128 11204 6180
rect 12624 6128 12676 6180
rect 14004 6128 14056 6180
rect 16120 6128 16172 6180
rect 18420 6196 18472 6248
rect 18604 6239 18656 6248
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 20168 6196 20220 6248
rect 19432 6171 19484 6180
rect 19432 6137 19441 6171
rect 19441 6137 19475 6171
rect 19475 6137 19484 6171
rect 19432 6128 19484 6137
rect 7748 6103 7800 6112
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 13636 6103 13688 6112
rect 13636 6069 13645 6103
rect 13645 6069 13679 6103
rect 13679 6069 13688 6103
rect 13636 6060 13688 6069
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16672 6060 16724 6112
rect 21456 6239 21508 6248
rect 21456 6205 21465 6239
rect 21465 6205 21499 6239
rect 21499 6205 21508 6239
rect 21456 6196 21508 6205
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 3332 5856 3384 5908
rect 4344 5899 4396 5908
rect 4344 5865 4353 5899
rect 4353 5865 4387 5899
rect 4387 5865 4396 5899
rect 4344 5856 4396 5865
rect 5448 5856 5500 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 10784 5856 10836 5908
rect 11244 5856 11296 5908
rect 12440 5899 12492 5908
rect 12440 5865 12449 5899
rect 12449 5865 12483 5899
rect 12483 5865 12492 5899
rect 12440 5856 12492 5865
rect 16028 5856 16080 5908
rect 18604 5856 18656 5908
rect 7472 5788 7524 5840
rect 8576 5788 8628 5840
rect 12164 5788 12216 5840
rect 15476 5831 15528 5840
rect 15476 5797 15485 5831
rect 15485 5797 15519 5831
rect 15519 5797 15528 5831
rect 15476 5788 15528 5797
rect 17316 5831 17368 5840
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 19156 5788 19208 5840
rect 20168 5856 20220 5908
rect 21088 5831 21140 5840
rect 21088 5797 21097 5831
rect 21097 5797 21131 5831
rect 21131 5797 21140 5831
rect 21088 5788 21140 5797
rect 21732 5788 21784 5840
rect 2228 5720 2280 5772
rect 2872 5720 2924 5772
rect 4988 5720 5040 5772
rect 6184 5720 6236 5772
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 10140 5720 10192 5772
rect 11152 5763 11204 5772
rect 11152 5729 11161 5763
rect 11161 5729 11195 5763
rect 11195 5729 11204 5763
rect 11152 5720 11204 5729
rect 12624 5720 12676 5772
rect 19064 5720 19116 5772
rect 19248 5763 19300 5772
rect 19248 5729 19257 5763
rect 19257 5729 19291 5763
rect 19291 5729 19300 5763
rect 19248 5720 19300 5729
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 18236 5652 18288 5704
rect 19524 5695 19576 5704
rect 19524 5661 19533 5695
rect 19533 5661 19567 5695
rect 19567 5661 19576 5695
rect 19524 5652 19576 5661
rect 21456 5652 21508 5704
rect 7380 5584 7432 5636
rect 10968 5584 11020 5636
rect 13912 5584 13964 5636
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 8116 5559 8168 5568
rect 8116 5525 8125 5559
rect 8125 5525 8159 5559
rect 8159 5525 8168 5559
rect 8116 5516 8168 5525
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 14464 5559 14516 5568
rect 13820 5516 13872 5525
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 16212 5516 16264 5568
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 20720 5516 20772 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1860 5312 1912 5364
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 2872 5312 2924 5364
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 8024 5312 8076 5364
rect 9220 5312 9272 5364
rect 12164 5312 12216 5364
rect 12624 5312 12676 5364
rect 14464 5312 14516 5364
rect 15384 5312 15436 5364
rect 19064 5355 19116 5364
rect 19064 5321 19073 5355
rect 19073 5321 19107 5355
rect 19107 5321 19116 5355
rect 19064 5312 19116 5321
rect 19432 5312 19484 5364
rect 21088 5312 21140 5364
rect 7840 5244 7892 5296
rect 7288 5176 7340 5228
rect 11796 5244 11848 5296
rect 10140 5176 10192 5228
rect 12532 5176 12584 5228
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 8024 5151 8076 5160
rect 8024 5117 8033 5151
rect 8033 5117 8067 5151
rect 8067 5117 8076 5151
rect 8024 5108 8076 5117
rect 8300 5151 8352 5160
rect 8300 5117 8309 5151
rect 8309 5117 8343 5151
rect 8343 5117 8352 5151
rect 8300 5108 8352 5117
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 1676 5040 1728 5092
rect 10876 5083 10928 5092
rect 10876 5049 10885 5083
rect 10885 5049 10919 5083
rect 10919 5049 10928 5083
rect 10876 5040 10928 5049
rect 10968 5083 11020 5092
rect 10968 5049 10977 5083
rect 10977 5049 11011 5083
rect 11011 5049 11020 5083
rect 10968 5040 11020 5049
rect 12808 5040 12860 5092
rect 21456 5244 21508 5296
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 14188 5040 14240 5092
rect 15476 5176 15528 5228
rect 19524 5176 19576 5228
rect 20720 5176 20772 5228
rect 16304 5108 16356 5160
rect 16672 5040 16724 5092
rect 18144 5083 18196 5092
rect 18144 5049 18153 5083
rect 18153 5049 18187 5083
rect 18187 5049 18196 5083
rect 18144 5040 18196 5049
rect 18788 5083 18840 5092
rect 17316 4972 17368 5024
rect 18788 5049 18797 5083
rect 18797 5049 18831 5083
rect 18831 5049 18840 5083
rect 18788 5040 18840 5049
rect 19432 5040 19484 5092
rect 21548 5083 21600 5092
rect 21548 5049 21557 5083
rect 21557 5049 21591 5083
rect 21591 5049 21600 5083
rect 21548 5040 21600 5049
rect 20904 4972 20956 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1676 4768 1728 4820
rect 9956 4768 10008 4820
rect 10692 4768 10744 4820
rect 10876 4811 10928 4820
rect 10876 4777 10885 4811
rect 10885 4777 10919 4811
rect 10919 4777 10928 4811
rect 10876 4768 10928 4777
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 13084 4768 13136 4820
rect 14188 4811 14240 4820
rect 12164 4700 12216 4752
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 15384 4768 15436 4820
rect 16028 4768 16080 4820
rect 17224 4768 17276 4820
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 19524 4768 19576 4820
rect 16764 4700 16816 4752
rect 17868 4700 17920 4752
rect 19432 4700 19484 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 8852 4632 8904 4684
rect 9220 4632 9272 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 9956 4675 10008 4684
rect 9956 4641 9965 4675
rect 9965 4641 9999 4675
rect 9999 4641 10008 4675
rect 9956 4632 10008 4641
rect 15384 4632 15436 4684
rect 17224 4632 17276 4684
rect 19064 4632 19116 4684
rect 20076 4700 20128 4752
rect 21548 4632 21600 4684
rect 11336 4607 11388 4616
rect 11336 4573 11345 4607
rect 11345 4573 11379 4607
rect 11379 4573 11388 4607
rect 11336 4564 11388 4573
rect 13452 4607 13504 4616
rect 7840 4496 7892 4548
rect 9772 4539 9824 4548
rect 9772 4505 9781 4539
rect 9781 4505 9815 4539
rect 9815 4505 9824 4539
rect 9772 4496 9824 4505
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 12808 4428 12860 4480
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 17500 4564 17552 4616
rect 13728 4496 13780 4548
rect 16396 4496 16448 4548
rect 14648 4428 14700 4480
rect 16304 4471 16356 4480
rect 16304 4437 16313 4471
rect 16313 4437 16347 4471
rect 16347 4437 16356 4471
rect 16304 4428 16356 4437
rect 17316 4428 17368 4480
rect 18880 4471 18932 4480
rect 18880 4437 18889 4471
rect 18889 4437 18923 4471
rect 18923 4437 18932 4471
rect 18880 4428 18932 4437
rect 20996 4428 21048 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 112 4224 164 4276
rect 1400 4224 1452 4276
rect 7196 4224 7248 4276
rect 7932 4088 7984 4140
rect 8484 4131 8536 4140
rect 7564 3884 7616 3936
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 9956 4224 10008 4276
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 12164 4224 12216 4276
rect 12808 4267 12860 4276
rect 12808 4233 12817 4267
rect 12817 4233 12851 4267
rect 12851 4233 12860 4267
rect 12808 4224 12860 4233
rect 13084 4267 13136 4276
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 15384 4267 15436 4276
rect 15384 4233 15393 4267
rect 15393 4233 15427 4267
rect 15427 4233 15436 4267
rect 15384 4224 15436 4233
rect 16764 4267 16816 4276
rect 16764 4233 16773 4267
rect 16773 4233 16807 4267
rect 16807 4233 16816 4267
rect 16764 4224 16816 4233
rect 17132 4224 17184 4276
rect 17868 4267 17920 4276
rect 17868 4233 17877 4267
rect 17877 4233 17911 4267
rect 17911 4233 17920 4267
rect 17868 4224 17920 4233
rect 18880 4224 18932 4276
rect 19432 4224 19484 4276
rect 20904 4224 20956 4276
rect 9772 4199 9824 4208
rect 9772 4165 9781 4199
rect 9781 4165 9815 4199
rect 9815 4165 9824 4199
rect 9772 4156 9824 4165
rect 9680 4088 9732 4140
rect 15660 4156 15712 4208
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 18788 4088 18840 4140
rect 19984 4156 20036 4208
rect 20076 4156 20128 4208
rect 20996 4088 21048 4140
rect 7840 4020 7892 4029
rect 10692 4020 10744 4072
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 15752 4063 15804 4072
rect 15752 4029 15761 4063
rect 15761 4029 15795 4063
rect 15795 4029 15804 4063
rect 15752 4020 15804 4029
rect 16028 4020 16080 4072
rect 11336 3952 11388 4004
rect 13820 3952 13872 4004
rect 15568 3952 15620 4004
rect 19248 3995 19300 4004
rect 19248 3961 19257 3995
rect 19257 3961 19291 3995
rect 19291 3961 19300 3995
rect 19248 3952 19300 3961
rect 19432 3952 19484 4004
rect 20904 3995 20956 4004
rect 20904 3961 20913 3995
rect 20913 3961 20947 3995
rect 20947 3961 20956 3995
rect 21456 3995 21508 4004
rect 20904 3952 20956 3961
rect 21456 3961 21465 3995
rect 21465 3961 21499 3995
rect 21499 3961 21508 3995
rect 21456 3952 21508 3961
rect 8024 3884 8076 3936
rect 13452 3884 13504 3936
rect 17132 3884 17184 3936
rect 17224 3884 17276 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 11244 3680 11296 3732
rect 13636 3723 13688 3732
rect 13636 3689 13645 3723
rect 13645 3689 13679 3723
rect 13679 3689 13688 3723
rect 13636 3680 13688 3689
rect 15752 3723 15804 3732
rect 15752 3689 15761 3723
rect 15761 3689 15795 3723
rect 15795 3689 15804 3723
rect 15752 3680 15804 3689
rect 19248 3723 19300 3732
rect 19248 3689 19257 3723
rect 19257 3689 19291 3723
rect 19291 3689 19300 3723
rect 19248 3680 19300 3689
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 8668 3612 8720 3664
rect 9128 3612 9180 3664
rect 13820 3612 13872 3664
rect 16212 3612 16264 3664
rect 16396 3655 16448 3664
rect 16396 3621 16405 3655
rect 16405 3621 16439 3655
rect 16439 3621 16448 3655
rect 16396 3612 16448 3621
rect 17316 3655 17368 3664
rect 17316 3621 17325 3655
rect 17325 3621 17359 3655
rect 17359 3621 17368 3655
rect 17316 3612 17368 3621
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 8392 3544 8444 3596
rect 13084 3544 13136 3596
rect 13728 3544 13780 3596
rect 15292 3544 15344 3596
rect 20996 3544 21048 3596
rect 3148 3476 3200 3528
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 21456 3476 21508 3528
rect 5448 3408 5500 3460
rect 7840 3408 7892 3460
rect 8116 3451 8168 3460
rect 8116 3417 8125 3451
rect 8125 3417 8159 3451
rect 8159 3417 8168 3451
rect 8116 3408 8168 3417
rect 12440 3340 12492 3392
rect 18788 3340 18840 3392
rect 20628 3340 20680 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 10048 3136 10100 3188
rect 13084 3179 13136 3188
rect 13084 3145 13093 3179
rect 13093 3145 13127 3179
rect 13127 3145 13136 3179
rect 13084 3136 13136 3145
rect 14004 3136 14056 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 17316 3136 17368 3188
rect 20812 3136 20864 3188
rect 20996 3179 21048 3188
rect 20996 3145 21005 3179
rect 21005 3145 21039 3179
rect 21039 3145 21048 3179
rect 20996 3136 21048 3145
rect 22468 3136 22520 3188
rect 8116 3068 8168 3120
rect 9588 3000 9640 3052
rect 17224 3000 17276 3052
rect 18144 3000 18196 3052
rect 8392 2975 8444 2984
rect 8392 2941 8401 2975
rect 8401 2941 8435 2975
rect 8435 2941 8444 2975
rect 8392 2932 8444 2941
rect 10048 2932 10100 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12532 2932 12584 2984
rect 8852 2864 8904 2916
rect 3148 2796 3200 2848
rect 7564 2839 7616 2848
rect 7564 2805 7573 2839
rect 7573 2805 7607 2839
rect 7607 2805 7616 2839
rect 7564 2796 7616 2805
rect 9220 2796 9272 2848
rect 12900 2796 12952 2848
rect 21364 2932 21416 2984
rect 14188 2839 14240 2848
rect 14188 2805 14197 2839
rect 14197 2805 14231 2839
rect 14231 2805 14240 2839
rect 14188 2796 14240 2805
rect 18788 2839 18840 2848
rect 18788 2805 18797 2839
rect 18797 2805 18831 2839
rect 18831 2805 18840 2839
rect 18788 2796 18840 2805
rect 25412 2796 25464 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 7564 2592 7616 2644
rect 8392 2592 8444 2644
rect 8944 2592 8996 2644
rect 21272 2592 21324 2644
rect 21916 2592 21968 2644
rect 22284 2592 22336 2644
rect 8852 2524 8904 2576
rect 22192 2524 22244 2576
rect 9220 2456 9272 2508
rect 9128 2320 9180 2372
rect 14188 2456 14240 2508
rect 20076 2456 20128 2508
rect 14372 2320 14424 2372
rect 11428 2252 11480 2304
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 15660 2252 15712 2304
rect 20076 2295 20128 2304
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 24216 2388 24268 2440
rect 22652 2252 22704 2304
rect 26884 2252 26936 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 6184 76 6236 128
rect 7472 76 7524 128
<< metal2 >>
rect 308 27526 704 27554
rect 110 24712 166 24721
rect 110 24647 166 24656
rect 124 23322 152 24647
rect 308 23474 336 27526
rect 676 27520 704 27526
rect 754 27520 810 28000
rect 1964 27526 2176 27554
rect 676 27492 796 27520
rect 1122 25528 1178 25537
rect 1122 25463 1178 25472
rect 1136 23730 1164 25463
rect 1124 23724 1176 23730
rect 1124 23666 1176 23672
rect 216 23446 336 23474
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 112 23316 164 23322
rect 112 23258 164 23264
rect 110 19680 166 19689
rect 110 19615 166 19624
rect 124 18902 152 19615
rect 112 18896 164 18902
rect 112 18838 164 18844
rect 112 17196 164 17202
rect 112 17138 164 17144
rect 124 17105 152 17138
rect 110 17096 166 17105
rect 110 17031 166 17040
rect 112 14000 164 14006
rect 112 13942 164 13948
rect 124 13297 152 13942
rect 110 13288 166 13297
rect 110 13223 166 13232
rect 112 12436 164 12442
rect 112 12378 164 12384
rect 124 12073 152 12378
rect 110 12064 166 12073
rect 110 11999 166 12008
rect 112 11552 164 11558
rect 112 11494 164 11500
rect 124 10713 152 11494
rect 110 10704 166 10713
rect 110 10639 166 10648
rect 216 8906 244 23446
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1688 22642 1716 23122
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1688 22545 1716 22578
rect 1674 22536 1730 22545
rect 1674 22471 1730 22480
rect 1490 21720 1546 21729
rect 1490 21655 1546 21664
rect 1504 18970 1532 21655
rect 1582 20360 1638 20369
rect 1582 20295 1638 20304
rect 1596 19514 1624 20295
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1504 18222 1532 18906
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 1676 18080 1728 18086
rect 1582 18048 1638 18057
rect 1676 18022 1728 18028
rect 1582 17983 1638 17992
rect 1596 17882 1624 17983
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1412 17134 1440 17682
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 14618 1532 16934
rect 1688 16794 1716 18022
rect 1780 17610 1808 23462
rect 1964 18834 1992 27526
rect 2148 27520 2176 27526
rect 2226 27520 2282 28000
rect 3698 27554 3754 28000
rect 3698 27526 3924 27554
rect 3698 27520 3754 27526
rect 2148 27492 2268 27520
rect 2226 26752 2282 26761
rect 2226 26687 2282 26696
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1964 18426 1992 18770
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1688 16114 1716 16730
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1780 15978 1808 16390
rect 1872 16114 1900 16594
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1872 15638 1900 16050
rect 1860 15632 1912 15638
rect 1860 15574 1912 15580
rect 1872 15162 1900 15574
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1504 13938 1532 14554
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1596 12986 1624 13738
rect 1688 13462 1716 14758
rect 2136 14340 2188 14346
rect 2136 14282 2188 14288
rect 2148 13938 2176 14282
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1688 12374 1716 13398
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12374 2084 12718
rect 1676 12368 1728 12374
rect 1676 12310 1728 12316
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11694 1440 12038
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 204 8900 256 8906
rect 204 8842 256 8848
rect 112 8560 164 8566
rect 112 8502 164 8508
rect 124 8265 152 8502
rect 110 8256 166 8265
rect 110 8191 166 8200
rect 1412 8090 1440 11630
rect 1688 11286 1716 12310
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 9178 1532 10610
rect 1688 10538 1716 10950
rect 1964 10674 1992 10950
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1676 10532 1728 10538
rect 1676 10474 1728 10480
rect 1688 9722 1716 10474
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 110 4448 166 4457
rect 110 4383 166 4392
rect 124 4282 152 4383
rect 112 4276 164 4282
rect 112 4218 164 4224
rect 662 82 718 480
rect 952 82 980 7754
rect 1596 7546 1624 8871
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 7818 1716 8366
rect 1780 7954 1808 10406
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1596 6866 1624 7278
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1688 6458 1716 7414
rect 1780 7002 1808 7890
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1872 5370 1900 9386
rect 1964 9178 1992 9454
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8498 2176 8910
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2148 8090 2176 8434
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2240 6458 2268 26687
rect 3896 19514 3924 27526
rect 5170 27520 5226 28000
rect 6642 27520 6698 28000
rect 7760 27526 8064 27554
rect 5184 19922 5212 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6092 23656 6144 23662
rect 6092 23598 6144 23604
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6104 19514 6132 23598
rect 6550 23488 6606 23497
rect 6656 23474 6684 27520
rect 6606 23446 6684 23474
rect 6550 23423 6606 23432
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 3896 19310 3924 19450
rect 3884 19304 3936 19310
rect 6656 19281 6684 19858
rect 3884 19246 3936 19252
rect 6642 19272 6698 19281
rect 6642 19207 6698 19216
rect 6656 19174 6684 19207
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2424 15638 2452 15914
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 2332 13530 2360 14486
rect 2424 14414 2452 15574
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2516 13814 2544 19110
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2608 17202 2636 17682
rect 3344 17338 3372 18090
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 3344 17134 3372 17274
rect 3620 17202 3648 17478
rect 4724 17338 4752 18022
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2700 15706 2728 16934
rect 3988 16454 4016 17002
rect 4816 16946 4844 18566
rect 5184 18426 5212 18770
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17338 5120 17478
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4894 17232 4950 17241
rect 4894 17167 4950 17176
rect 4724 16918 4844 16946
rect 4724 16590 4752 16918
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2884 14074 2912 14350
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2976 13870 3004 15302
rect 2424 13786 2544 13814
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2332 12782 2360 13466
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2424 12646 2452 13786
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2516 11898 2544 12310
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2424 10810 2452 11222
rect 2516 11082 2544 11834
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2424 10198 2452 10746
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2332 9178 2360 9998
rect 2424 9722 2452 10134
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2608 9518 2636 10202
rect 2700 9926 2728 11562
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2792 10810 2820 11086
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2700 9042 2728 9454
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2700 8634 2728 8978
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8634 2820 8774
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2504 8016 2556 8022
rect 2424 7976 2504 8004
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2226 6352 2282 6361
rect 2226 6287 2282 6296
rect 2240 5778 2268 6287
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2240 5370 2268 5714
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 1858 5264 1914 5273
rect 1858 5199 1914 5208
rect 1872 5166 1900 5199
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1688 4826 1716 5034
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 4282 1440 4626
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 662 54 980 82
rect 2042 82 2098 480
rect 2332 82 2360 7210
rect 2424 7206 2452 7976
rect 2504 7958 2556 7964
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2516 7546 2544 7822
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 6934 2452 7142
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2516 6322 2544 7482
rect 2608 6798 2636 7822
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6458 2636 6734
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2884 5778 2912 12582
rect 3344 12288 3372 15846
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 13530 3464 14894
rect 3804 14890 3832 15574
rect 3988 15026 4016 16390
rect 4356 16046 4384 16390
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15638 4200 15846
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 15094 4108 15438
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 4080 14618 4108 15030
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4264 14278 4292 14418
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3528 12986 3556 13942
rect 4264 13870 4292 14214
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4264 13376 4292 13806
rect 4356 13734 4384 15982
rect 4528 15972 4580 15978
rect 4448 15932 4528 15960
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4344 13388 4396 13394
rect 4264 13348 4344 13376
rect 4344 13330 4396 13336
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3712 12646 3740 13262
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3804 12442 3832 13126
rect 4356 12646 4384 13330
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3516 12300 3568 12306
rect 3344 12260 3516 12288
rect 3516 12242 3568 12248
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 2976 11762 3004 12106
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 10742 3004 11698
rect 3344 11014 3372 12106
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2976 9722 3004 10678
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 3160 10266 3188 10474
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2976 6458 3004 6802
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3344 5914 3372 10950
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 6458 3464 9862
rect 3528 9178 3556 12242
rect 4356 12238 4384 12582
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3896 10266 3924 11222
rect 4172 10810 4200 11290
rect 4356 11218 4384 12174
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4356 10810 4384 11154
rect 4160 10804 4212 10810
rect 4344 10804 4396 10810
rect 4160 10746 4212 10752
rect 4264 10764 4344 10792
rect 4264 10690 4292 10764
rect 4344 10746 4396 10752
rect 4080 10662 4292 10690
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 4080 10130 4108 10662
rect 4068 10124 4120 10130
rect 4120 10084 4200 10112
rect 4068 10066 4120 10072
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3988 8974 4016 9930
rect 4172 9382 4200 10084
rect 4344 10056 4396 10062
rect 4264 10016 4344 10044
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4264 9042 4292 10016
rect 4344 9998 4396 10004
rect 4448 9450 4476 15932
rect 4528 15914 4580 15920
rect 4724 15706 4752 16526
rect 4816 16114 4844 16662
rect 4908 16425 4936 17167
rect 4988 17060 5040 17066
rect 4988 17002 5040 17008
rect 5000 16590 5028 17002
rect 5092 16998 5120 17274
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 4988 16584 5040 16590
rect 5184 16561 5212 18362
rect 6288 17882 6316 18702
rect 6380 18426 6408 18838
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6366 18184 6422 18193
rect 6366 18119 6422 18128
rect 6380 18086 6408 18119
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 17338 5488 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 4988 16526 5040 16532
rect 5170 16552 5226 16561
rect 5170 16487 5226 16496
rect 4894 16416 4950 16425
rect 4894 16351 4950 16360
rect 5460 16250 5488 17274
rect 6380 16726 6408 17274
rect 6472 17066 6500 19110
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 17338 6592 18362
rect 6932 17814 6960 19110
rect 7024 18970 7052 19110
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6564 17066 6592 17274
rect 6460 17060 6512 17066
rect 6460 17002 6512 17008
rect 6552 17060 6604 17066
rect 6552 17002 6604 17008
rect 6368 16720 6420 16726
rect 6368 16662 6420 16668
rect 6472 16590 6500 17002
rect 6932 16794 6960 17750
rect 7116 17270 7144 20198
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 18970 7236 19654
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7208 18290 7236 18906
rect 7668 18902 7696 19314
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7760 18630 7788 27526
rect 8036 27418 8064 27526
rect 8114 27520 8170 28000
rect 9586 27520 9642 28000
rect 11058 27520 11114 28000
rect 12530 27554 12586 28000
rect 12530 27526 12664 27554
rect 12530 27520 12586 27526
rect 8128 27418 8156 27520
rect 8036 27390 8156 27418
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7852 19514 7880 19654
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7852 19310 7880 19450
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 8496 19242 8524 19722
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7564 18352 7616 18358
rect 7564 18294 7616 18300
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7392 17814 7420 18090
rect 7380 17808 7432 17814
rect 7380 17750 7432 17756
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7576 16726 7604 18294
rect 7656 17808 7708 17814
rect 7656 17750 7708 17756
rect 7668 17542 7696 17750
rect 7760 17678 7788 18294
rect 7852 17882 7880 18838
rect 7944 18086 7972 18838
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4816 15706 4844 16050
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 4816 15026 4844 15642
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 4908 15162 4936 15302
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 5552 14958 5580 15302
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6196 15026 6224 15302
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 4724 13870 4752 14418
rect 5092 13870 5120 14418
rect 5460 14006 5488 14418
rect 5552 14346 5580 14894
rect 6748 14618 6776 14962
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 4712 13864 4764 13870
rect 5080 13864 5132 13870
rect 4712 13806 4764 13812
rect 5000 13824 5080 13852
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4540 12850 4568 13330
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4540 12646 4568 12786
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4632 11898 4660 12718
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 5000 11218 5028 13824
rect 5080 13806 5132 13812
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5092 12986 5120 13330
rect 5368 13190 5396 13806
rect 5460 13376 5488 13942
rect 6564 13938 6592 14418
rect 6642 14376 6698 14385
rect 6642 14311 6698 14320
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6564 13841 6592 13874
rect 6550 13832 6606 13841
rect 6550 13767 6606 13776
rect 6460 13456 6512 13462
rect 6380 13416 6460 13444
rect 5540 13388 5592 13394
rect 5460 13348 5540 13376
rect 5540 13330 5592 13336
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5368 12782 5396 13126
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 11540 5396 12718
rect 5552 11898 5580 13330
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12646 5764 12854
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5736 12306 5764 12582
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5448 11552 5500 11558
rect 5368 11512 5448 11540
rect 5448 11494 5500 11500
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4988 11212 5040 11218
rect 4988 11154 5040 11160
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4540 9926 4568 10202
rect 4816 10130 4844 11154
rect 5000 10713 5028 11154
rect 4986 10704 5042 10713
rect 5042 10662 5120 10690
rect 4986 10639 5042 10648
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 5000 9994 5028 10406
rect 5092 10130 5120 10662
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4540 9042 4568 9318
rect 5092 9178 5120 10066
rect 5184 9926 5212 10542
rect 5460 10130 5488 11494
rect 5552 11218 5580 11834
rect 6012 11354 6040 12242
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6104 11558 6132 12174
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6196 11354 6224 12922
rect 6288 12714 6316 13126
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6380 12646 6408 13416
rect 6460 13398 6512 13404
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6288 11830 6316 12242
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10742 5580 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 6012 10266 6040 11290
rect 6196 10674 6224 11290
rect 6288 10742 6316 11766
rect 6380 11286 6408 12582
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 6184 10668 6236 10674
rect 6104 10628 6184 10656
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9518 5212 9862
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5184 9110 5212 9454
rect 5460 9382 5488 10066
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6104 9450 6132 10628
rect 6184 10610 6236 10616
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10198 6224 10406
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6196 9722 6224 10134
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8430 3832 8774
rect 3988 8634 4016 8910
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3528 7002 3556 7346
rect 3804 7002 3832 8366
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4172 7410 4200 8230
rect 4264 8090 4292 8978
rect 4540 8430 4568 8978
rect 5460 8634 5488 9318
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5552 8634 5580 8978
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8634 6040 8774
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4540 8090 4568 8366
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 4264 6934 4292 7142
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4264 6458 4292 6870
rect 4448 6798 4476 7822
rect 4540 7546 4568 8026
rect 5092 8022 5120 8366
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 3976 6248 4028 6254
rect 3974 6216 3976 6225
rect 4028 6216 4030 6225
rect 3974 6151 4030 6160
rect 3988 6118 4016 6151
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 4356 5914 4384 6666
rect 4724 6458 4752 7754
rect 5000 7410 5028 7822
rect 5092 7818 5120 7958
rect 5368 7954 5396 8502
rect 5460 8430 5488 8570
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5368 7002 5396 7890
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 5460 5914 5488 8366
rect 6196 7954 6224 9386
rect 6288 8022 6316 10678
rect 6656 10577 6684 14311
rect 6932 13734 6960 15302
rect 7024 14890 7052 15642
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 7116 13462 7144 16118
rect 7576 15706 7604 16662
rect 7668 16436 7696 17478
rect 7760 17270 7788 17614
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 7748 17264 7800 17270
rect 7748 17206 7800 17212
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7944 16726 7972 17002
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7748 16448 7800 16454
rect 7668 16408 7748 16436
rect 7748 16390 7800 16396
rect 7760 15978 7788 16390
rect 7944 16250 7972 16662
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7760 15162 7788 15914
rect 7944 15570 7972 16186
rect 8128 16114 8156 16526
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12850 6960 13126
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6932 12753 6960 12786
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6932 12209 6960 12242
rect 6918 12200 6974 12209
rect 6918 12135 6974 12144
rect 7024 12102 7052 13194
rect 7116 12850 7144 13398
rect 7208 13190 7236 13806
rect 7300 13705 7328 14826
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7392 13870 7420 14418
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7286 13696 7342 13705
rect 7286 13631 7342 13640
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7024 11762 7052 12038
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7116 11286 7144 12650
rect 7300 12374 7328 13631
rect 7392 13530 7420 13806
rect 8036 13734 8064 14418
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8024 13728 8076 13734
rect 7944 13688 8024 13716
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7300 11762 7328 12310
rect 7288 11756 7340 11762
rect 7340 11716 7420 11744
rect 7288 11698 7340 11704
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 6828 10600 6880 10606
rect 6642 10568 6698 10577
rect 6828 10542 6880 10548
rect 6642 10503 6698 10512
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10130 6592 10406
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9586 6408 9930
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6380 9178 6408 9522
rect 6564 9178 6592 10066
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6656 7954 6684 10503
rect 6840 10266 6868 10542
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6196 7342 6224 7890
rect 6656 7546 6684 7890
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6662 5580 7142
rect 5644 7002 5672 7210
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6254 5580 6598
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6322 6040 6870
rect 6196 6458 6224 7278
rect 6564 6934 6592 7346
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6564 6730 6592 6870
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 6196 5778 6224 6394
rect 6656 6322 6684 6734
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 2884 5370 2912 5714
rect 5000 5370 5028 5714
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 2884 5137 2912 5306
rect 2870 5128 2926 5137
rect 2870 5063 2926 5072
rect 5000 4154 5028 5306
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 4908 4126 5028 4154
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 3160 2854 3188 3470
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2042 54 2360 82
rect 3160 82 3188 2790
rect 4908 1193 4936 4126
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 3369 5488 3402
rect 5446 3360 5502 3369
rect 5446 3295 5502 3304
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5078 1864 5134 1873
rect 5078 1799 5134 1808
rect 4894 1184 4950 1193
rect 4894 1119 4950 1128
rect 3422 82 3478 480
rect 3160 54 3478 82
rect 662 0 718 54
rect 2042 0 2098 54
rect 3422 0 3478 54
rect 4802 82 4858 480
rect 5092 82 5120 1799
rect 4802 54 5120 82
rect 6182 128 6238 480
rect 6182 76 6184 128
rect 6236 76 6238 128
rect 6748 105 6776 9454
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9178 7328 9318
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7300 8498 7328 9114
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7392 8294 7420 11716
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7484 10606 7512 10950
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 10033 7512 10542
rect 7576 10470 7604 10950
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7470 10024 7526 10033
rect 7470 9959 7526 9968
rect 7576 9518 7604 10406
rect 7760 9654 7788 13126
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 9042 7604 9454
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7484 8362 7512 8910
rect 7576 8430 7604 8978
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7274 6960 7686
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 7012 7268 7064 7274
rect 7012 7210 7064 7216
rect 6932 7002 6960 7210
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7024 6662 7052 7210
rect 7392 6934 7420 8230
rect 7484 8090 7512 8298
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7300 6254 7328 6394
rect 7392 6390 7420 6598
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7288 6248 7340 6254
rect 7208 6208 7288 6236
rect 7208 4282 7236 6208
rect 7288 6190 7340 6196
rect 7760 6118 7788 9590
rect 7852 9518 7880 9998
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 9042 7880 9454
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7852 8634 7880 8978
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7944 6798 7972 13688
rect 8024 13670 8076 13676
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 11694 8064 12582
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 11218 8064 11630
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8036 9518 8064 10202
rect 8128 10130 8156 13738
rect 8220 12170 8248 17546
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8128 9722 8156 10066
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 9042 8064 9454
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8036 8090 8064 8978
rect 8128 8566 8156 9658
rect 8312 9586 8340 18566
rect 8496 18154 8524 18702
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8496 17678 8524 18090
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 16046 8524 16390
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 14890 8432 15846
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8496 13734 8524 15982
rect 8588 15570 8616 19314
rect 8680 16153 8708 20198
rect 9600 19514 9628 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 11072 23866 11100 27520
rect 12636 23866 12664 27526
rect 13740 27526 13952 27554
rect 13740 23866 13768 27526
rect 13924 27418 13952 27526
rect 14002 27520 14058 28000
rect 15474 27520 15530 28000
rect 16946 27520 17002 28000
rect 18418 27554 18474 28000
rect 18418 27526 18736 27554
rect 18418 27520 18474 27526
rect 14016 27418 14044 27520
rect 13924 27390 14044 27418
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15488 24614 15516 27520
rect 15476 24608 15528 24614
rect 15476 24550 15528 24556
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 12898 23760 12954 23769
rect 12898 23695 12954 23704
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9600 19310 9628 19450
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8956 18290 8984 19110
rect 9600 18290 9628 19246
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9876 18766 9904 19178
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9784 18358 9812 18702
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 8956 17882 8984 18226
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 8944 17876 8996 17882
rect 8944 17818 8996 17824
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8666 16144 8722 16153
rect 8666 16079 8722 16088
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 15162 8616 15506
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8680 15042 8708 16079
rect 8864 15706 8892 16934
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 9416 15366 9444 16526
rect 9508 16250 9536 17274
rect 9784 17066 9812 18090
rect 10152 18086 10180 18838
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9876 17338 9904 17750
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9784 15706 9812 17002
rect 10152 16794 10180 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10612 17338 10640 17614
rect 10980 17610 11008 18702
rect 10968 17604 11020 17610
rect 10968 17546 11020 17552
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10060 16250 10088 16730
rect 10888 16454 10916 17002
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10060 15978 10088 16186
rect 10888 16114 10916 16390
rect 10980 16182 11008 17546
rect 11532 17338 11560 23598
rect 12912 22778 12940 23695
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 13556 20058 13584 23598
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 16960 22778 16988 27520
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18902 11744 19110
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11612 18148 11664 18154
rect 11612 18090 11664 18096
rect 11624 17882 11652 18090
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11808 17377 11836 19246
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12268 17882 12296 18838
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12360 17814 12388 19110
rect 12440 18896 12492 18902
rect 12440 18838 12492 18844
rect 12452 18086 12480 18838
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 11794 17368 11850 17377
rect 11520 17332 11572 17338
rect 11794 17303 11850 17312
rect 11520 17274 11572 17280
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11624 16250 11652 16662
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 10060 15638 10088 15914
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 15632 10100 15638
rect 10048 15574 10100 15580
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 8588 15014 8708 15042
rect 9048 15026 9076 15302
rect 8760 15020 8812 15026
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 8404 11694 8432 12854
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8496 11286 8524 12038
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8496 10266 8524 11222
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7478 8156 7822
rect 8220 7546 8248 7958
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7300 5574 7328 6054
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5234 7328 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7392 5137 7420 5578
rect 7378 5128 7434 5137
rect 7378 5063 7434 5072
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 7484 134 7512 5782
rect 7852 5778 7880 6326
rect 8588 5846 8616 15014
rect 8760 14962 8812 14968
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8668 14340 8720 14346
rect 8668 14282 8720 14288
rect 8680 12986 8708 14282
rect 8772 13462 8800 14962
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9324 14618 9352 14826
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 8864 13870 8892 14554
rect 9416 14550 9444 15302
rect 9692 14618 9720 15438
rect 10152 15162 10180 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 11624 15638 11652 16186
rect 12084 15910 12112 16526
rect 12360 16522 12388 17070
rect 12452 16658 12480 18022
rect 12544 17202 12572 18566
rect 12728 18426 12756 19110
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12728 18086 12756 18362
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12820 17678 12848 18634
rect 13188 18290 13216 19858
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13924 18426 13952 18770
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13188 17678 13216 18226
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 12820 17202 12848 17614
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16794 12848 17138
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13188 16658 13216 17070
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13372 16590 13400 17614
rect 13556 16998 13584 17750
rect 13924 17241 13952 18362
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 13910 17232 13966 17241
rect 13910 17167 13966 17176
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 13372 16182 13400 16526
rect 13464 16250 13492 16662
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 14758
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10980 14550 11008 15302
rect 11256 14958 11284 15302
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 9404 14544 9456 14550
rect 10968 14544 11020 14550
rect 9404 14486 9456 14492
rect 10046 14512 10102 14521
rect 10968 14486 11020 14492
rect 10046 14447 10102 14456
rect 10692 14476 10744 14482
rect 10060 14414 10088 14447
rect 10692 14418 10744 14424
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10060 14074 10088 14350
rect 10140 14272 10192 14278
rect 10140 14214 10192 14220
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8772 12084 8800 12854
rect 8864 12850 8892 13806
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9048 13530 9076 13738
rect 9876 13734 9904 13806
rect 9864 13728 9916 13734
rect 9678 13696 9734 13705
rect 9864 13670 9916 13676
rect 9678 13631 9734 13640
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8852 12096 8904 12102
rect 8772 12056 8852 12084
rect 8852 12038 8904 12044
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 11286 8708 11494
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8864 10713 8892 12038
rect 8956 11898 8984 12854
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8956 11694 8984 11834
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 8850 10704 8906 10713
rect 8850 10639 8906 10648
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8680 10062 8708 10542
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8956 9518 8984 11630
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8680 8362 8708 8570
rect 8772 8498 8800 8910
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 8022 8800 8230
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7546 8984 7822
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8680 6866 8708 7142
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8680 6458 8708 6802
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 9048 6390 9076 13466
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12714 9260 13126
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12306 9260 12650
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 9232 11558 9260 12242
rect 9324 12209 9352 13466
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12986 9444 13262
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9310 12200 9366 12209
rect 9310 12135 9366 12144
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11014 9260 11494
rect 9324 11354 9352 12135
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10606 9260 10950
rect 9324 10606 9352 11290
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9232 10198 9260 10542
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9140 8294 9168 9046
rect 9324 9042 9352 10542
rect 9416 9081 9444 12922
rect 9692 11762 9720 13631
rect 9968 13394 9996 13806
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9692 11626 9720 11698
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11354 9720 11562
rect 9680 11348 9732 11354
rect 9732 11308 9812 11336
rect 9680 11290 9732 11296
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10538 9720 11086
rect 9784 10810 9812 11308
rect 9864 11280 9916 11286
rect 9968 11268 9996 13330
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 9916 11240 9996 11268
rect 9864 11222 9916 11228
rect 10060 10810 10088 12650
rect 10152 12374 10180 14214
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13394 10732 14418
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13870 11284 14214
rect 11440 14006 11468 15438
rect 11624 15162 11652 15574
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11520 14476 11572 14482
rect 11572 14436 11652 14464
rect 11520 14418 11572 14424
rect 11624 14278 11652 14436
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11624 13938 11652 14214
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11244 13864 11296 13870
rect 11296 13812 11468 13814
rect 11244 13806 11468 13812
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10152 11082 10180 12174
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10704 11354 10732 12718
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10796 11898 10824 12650
rect 10980 12306 11008 13330
rect 11072 13258 11100 13806
rect 11256 13786 11468 13806
rect 11440 13530 11468 13786
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11624 13394 11652 13874
rect 12084 13530 12112 15846
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12176 14890 12204 15098
rect 12268 14958 12296 15370
rect 13372 15366 13400 15846
rect 13556 15706 13584 16934
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14016 16182 14044 16526
rect 14004 16176 14056 16182
rect 14004 16118 14056 16124
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 15162 13400 15302
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12268 14550 12296 14894
rect 13648 14890 13676 15846
rect 13912 15632 13964 15638
rect 13912 15574 13964 15580
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 12820 14550 12848 14826
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12268 13394 12296 13670
rect 12452 13530 12480 13806
rect 12820 13530 12848 14486
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11354 10916 11630
rect 10980 11354 11008 12106
rect 11348 11898 11376 12310
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11440 11626 11468 12310
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 10692 11348 10744 11354
rect 10876 11348 10928 11354
rect 10744 11308 10824 11336
rect 10692 11290 10744 11296
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10152 10674 10180 11018
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10704 10538 10732 10746
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 9692 10266 9720 10474
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 10796 10198 10824 11308
rect 10876 11290 10928 11296
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11532 11150 11560 13262
rect 11624 12986 11652 13330
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 12268 12918 12296 13330
rect 12256 12912 12308 12918
rect 12256 12854 12308 12860
rect 12452 12782 12480 13466
rect 13004 12850 13032 14826
rect 13924 14822 13952 15574
rect 14292 15026 14320 18022
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14646 17368 14702 17377
rect 14956 17360 15252 17380
rect 15396 17338 15424 17682
rect 14646 17303 14702 17312
rect 15384 17332 15436 17338
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 15910 14412 16050
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15502 14412 15846
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14384 15026 14412 15438
rect 14660 15026 14688 17303
rect 15384 17274 15436 17280
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16594
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14922 16144 14978 16153
rect 14922 16079 14978 16088
rect 14936 16046 14964 16079
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14752 15366 14780 15642
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 13938 13124 14350
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13280 13870 13308 14554
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12850 13492 13262
rect 13648 12918 13676 13806
rect 13924 13462 13952 14758
rect 14108 14346 14136 14758
rect 14292 14618 14320 14962
rect 14752 14618 14780 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 15304 13814 15332 14282
rect 15396 13938 15424 17274
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15580 16726 15608 17002
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15488 15910 15516 16594
rect 15672 15978 15700 17070
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 14384 13530 14412 13806
rect 15304 13786 15424 13814
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13912 13456 13964 13462
rect 13912 13398 13964 13404
rect 13832 12986 13860 13398
rect 15396 13394 15424 13786
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15396 12986 15424 13330
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 13636 12912 13688 12918
rect 13636 12854 13688 12860
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 13004 12442 13032 12786
rect 13648 12782 13676 12854
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12728 11558 12756 12106
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9450 9904 9862
rect 10704 9654 10732 9998
rect 10796 9722 10824 10134
rect 10980 10062 11008 10610
rect 11532 10266 11560 11086
rect 11624 10470 11652 11222
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11992 10266 12020 11018
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10538 12572 10950
rect 12728 10742 12756 11494
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12820 10674 12848 12174
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12176 10130 12204 10202
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 9588 9376 9640 9382
rect 9876 9353 9904 9386
rect 9588 9318 9640 9324
rect 9862 9344 9918 9353
rect 9600 9110 9628 9318
rect 9862 9279 9918 9288
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9588 9104 9640 9110
rect 9402 9072 9458 9081
rect 9312 9036 9364 9042
rect 9232 8996 9312 9024
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 6866 9168 8230
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6384 9088 6390
rect 9088 6344 9168 6372
rect 9036 6326 9088 6332
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5302 7880 5714
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7852 4554 7880 5238
rect 8036 5166 8064 5306
rect 8024 5160 8076 5166
rect 8024 5102 8076 5108
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7852 4078 7880 4490
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4146 7972 4422
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 2854 7604 3878
rect 7852 3466 7880 4014
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3602 8064 3878
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 8036 3194 8064 3538
rect 8128 3466 8156 5510
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8312 4690 8340 5102
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8312 3584 8340 4626
rect 8482 4176 8538 4185
rect 8482 4111 8484 4120
rect 8536 4111 8538 4120
rect 8484 4082 8536 4088
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8392 3596 8444 3602
rect 8312 3556 8392 3584
rect 8392 3538 8444 3544
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8128 3126 8156 3402
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8404 2990 8432 3538
rect 8680 3505 8708 3606
rect 8666 3496 8722 3505
rect 8666 3431 8722 3440
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7576 2650 7604 2790
rect 8404 2650 8432 2926
rect 8864 2922 8892 4626
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 7576 2417 7604 2586
rect 8864 2582 8892 2858
rect 8956 2650 8984 6258
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 4185 9076 6054
rect 9034 4176 9090 4185
rect 9034 4111 9090 4120
rect 9140 3670 9168 6344
rect 9232 5370 9260 8996
rect 9588 9046 9640 9052
rect 9954 9072 10010 9081
rect 9402 9007 9458 9016
rect 9954 9007 10010 9016
rect 9312 8978 9364 8984
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9416 8090 9444 8434
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 8090 9536 8366
rect 9784 8362 9812 8570
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 7274 9536 7754
rect 9600 7274 9628 8230
rect 9876 7886 9904 8842
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9508 7002 9536 7210
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4690 9260 5306
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 9600 3058 9628 6734
rect 9968 4826 9996 9007
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 7478 10088 7822
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9692 4146 9720 4626
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9784 4214 9812 4490
rect 9968 4282 9996 4626
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 10060 3194 10088 7414
rect 10152 7206 10180 7958
rect 10704 7818 10732 9386
rect 11808 9042 11836 9522
rect 12176 9382 12204 10066
rect 12544 9761 12572 10474
rect 12716 10464 12768 10470
rect 12636 10424 12716 10452
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12636 9518 12664 10424
rect 12716 10406 12768 10412
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12728 9178 12756 10066
rect 12820 9654 12848 10610
rect 13004 10538 13032 11086
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10796 8634 10824 8910
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 11256 8566 11284 8910
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10796 7206 10824 7822
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10152 6934 10180 7142
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6458 10364 6802
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10796 5914 10824 7142
rect 11256 7002 11284 8502
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11440 8022 11468 8366
rect 11808 8294 11836 8978
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11428 8016 11480 8022
rect 11428 7958 11480 7964
rect 11440 7546 11468 7958
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11256 6254 11284 6938
rect 11440 6934 11468 7482
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11624 6458 11652 6734
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5817 10916 6190
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 10874 5808 10930 5817
rect 10140 5772 10192 5778
rect 11164 5778 11192 6122
rect 11256 5914 11284 6190
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 10874 5743 10930 5752
rect 11152 5772 11204 5778
rect 10140 5714 10192 5720
rect 11152 5714 11204 5720
rect 10152 5234 10180 5714
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10980 5098 11008 5578
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10888 4826 10916 5034
rect 11164 4826 11192 5714
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10138 4720 10194 4729
rect 10138 4655 10194 4664
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 10060 2990 10088 3130
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 9232 2514 9260 2790
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 7562 2408 7618 2417
rect 7562 2343 7618 2352
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 7562 2000 7618 2009
rect 7562 1935 7618 1944
rect 7472 128 7524 134
rect 4802 0 4858 54
rect 6182 0 6238 76
rect 6734 96 6790 105
rect 7472 70 7524 76
rect 7576 82 7604 1935
rect 7654 82 7710 480
rect 7576 54 7710 82
rect 6734 31 6790 40
rect 7654 0 7710 54
rect 9034 82 9090 480
rect 9140 82 9168 2314
rect 9034 54 9168 82
rect 10152 82 10180 4655
rect 10704 4282 10732 4762
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10704 4078 10732 4218
rect 11256 4078 11284 5850
rect 11808 5302 11836 8230
rect 11888 7336 11940 7342
rect 11886 7304 11888 7313
rect 11940 7304 11942 7313
rect 11886 7239 11942 7248
rect 11900 7206 11928 7239
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6322 12020 6734
rect 12176 6458 12204 8298
rect 12820 8090 12848 8910
rect 12912 8498 12940 9998
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13004 9722 13032 9930
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 12268 7546 12296 7890
rect 12912 7546 12940 7958
rect 12992 7812 13044 7818
rect 13096 7800 13124 12718
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13188 11830 13216 12378
rect 14752 12374 14780 12922
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14740 12368 14792 12374
rect 14740 12310 14792 12316
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13542 11792 13598 11801
rect 13188 7954 13216 11766
rect 13542 11727 13598 11736
rect 13556 11626 13584 11727
rect 13832 11694 13860 12106
rect 14476 11762 14504 12310
rect 14752 11898 14780 12310
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13464 11218 13492 11562
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13464 10810 13492 11154
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13268 9172 13320 9178
rect 13372 9160 13400 10066
rect 13556 10010 13584 11562
rect 13818 10704 13874 10713
rect 13818 10639 13874 10648
rect 13832 10606 13860 10639
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14108 10130 14136 10542
rect 14476 10266 14504 11698
rect 14752 11558 14780 11834
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14936 11354 14964 11630
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15488 10674 15516 15846
rect 15764 15570 15792 22714
rect 18050 22536 18106 22545
rect 18050 22471 18106 22480
rect 18064 22438 18092 22471
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 16578 19272 16634 19281
rect 16578 19207 16634 19216
rect 16592 18222 16620 19207
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15764 15162 15792 15506
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15856 15094 15884 15642
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 13841 15700 14758
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15672 12102 15700 13767
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15856 11830 15884 15030
rect 15948 14550 15976 17478
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 16040 15706 16068 15982
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 14822 16252 15574
rect 16316 15570 16344 18158
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16500 16046 16528 16526
rect 16684 16114 16712 16526
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16500 14958 16528 15982
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16500 14618 16528 14894
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 15936 14544 15988 14550
rect 15936 14486 15988 14492
rect 15948 14074 15976 14486
rect 16776 14414 16804 19110
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 17052 17882 17080 18294
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17040 17876 17092 17882
rect 17040 17818 17092 17824
rect 17512 17814 17540 18226
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 17512 17338 17540 17750
rect 17696 17338 17724 18702
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17512 16794 17540 17274
rect 18248 17048 18276 18022
rect 18340 17882 18368 18090
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 18432 17542 18460 17750
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18328 17060 18380 17066
rect 18248 17020 18328 17048
rect 18328 17002 18380 17008
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17052 15910 17080 16730
rect 18340 16522 18368 17002
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 18432 16182 18460 17478
rect 18524 17202 18552 17614
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18524 16590 18552 17138
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18524 16250 18552 16526
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18420 16176 18472 16182
rect 18420 16118 18472 16124
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15638 17080 15846
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17420 15162 17448 15438
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16408 13938 16436 14282
rect 16776 14074 16804 14350
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 15948 13802 15976 13874
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15948 12714 15976 12854
rect 16040 12753 16068 13874
rect 16868 13394 16896 15098
rect 17420 14618 17448 15098
rect 18064 15026 18092 15302
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17328 14074 17356 14418
rect 17788 14074 17816 14418
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16212 13252 16264 13258
rect 16212 13194 16264 13200
rect 16026 12744 16082 12753
rect 15936 12708 15988 12714
rect 16224 12714 16252 13194
rect 16868 12986 16896 13330
rect 17132 13184 17184 13190
rect 17132 13126 17184 13132
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16026 12679 16082 12688
rect 16212 12708 16264 12714
rect 15936 12650 15988 12656
rect 16212 12650 16264 12656
rect 15948 12442 15976 12650
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15672 11286 15700 11494
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15580 10810 15608 11086
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15672 10742 15700 11222
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14096 10124 14148 10130
rect 15580 10112 15608 10542
rect 15672 10266 15700 10678
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15856 10130 15884 11766
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 10606 15976 11698
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15948 10470 15976 10542
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15660 10124 15712 10130
rect 15580 10084 15660 10112
rect 14096 10066 14148 10072
rect 15660 10066 15712 10072
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 14108 10033 14136 10066
rect 13464 9982 13584 10010
rect 13726 10024 13782 10033
rect 13636 9988 13688 9994
rect 13464 9722 13492 9982
rect 13726 9959 13782 9968
rect 14094 10024 14150 10033
rect 14094 9959 14150 9968
rect 13636 9930 13688 9936
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13648 9586 13676 9930
rect 13740 9722 13768 9959
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13452 9172 13504 9178
rect 13372 9132 13452 9160
rect 13268 9114 13320 9120
rect 13452 9114 13504 9120
rect 13280 8566 13308 9114
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13280 8362 13308 8502
rect 13648 8362 13676 9318
rect 13924 9042 13952 9386
rect 13912 9036 13964 9042
rect 13964 8996 14044 9024
rect 13912 8978 13964 8984
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13044 7772 13124 7800
rect 12992 7754 13044 7760
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 13004 7002 13032 7754
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 13096 7002 13124 7210
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 6458 13124 6938
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12176 6254 12204 6394
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12176 5846 12204 6190
rect 12452 5914 12480 6258
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12176 5370 12204 5782
rect 12636 5778 12664 6122
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12636 5370 12664 5714
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 12176 4758 12204 5306
rect 13358 5264 13414 5273
rect 12532 5228 12584 5234
rect 13358 5199 13414 5208
rect 12532 5170 12584 5176
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 11256 3738 11284 4014
rect 11348 4010 11376 4558
rect 12176 4282 12204 4694
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 2990 12480 3334
rect 12544 2990 12572 5170
rect 13372 5166 13400 5199
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12820 4486 12848 5034
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4282 12848 4422
rect 13096 4282 13124 4762
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13372 4154 13400 5102
rect 13464 4622 13492 7346
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13924 6934 13952 7278
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13648 6118 13676 6666
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13372 4126 13492 4154
rect 13464 3942 13492 4126
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13648 3738 13676 6054
rect 13924 5642 13952 6870
rect 14016 6458 14044 8996
rect 14844 8498 14872 9386
rect 15672 9382 15700 10066
rect 15856 9722 15884 10066
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15672 8498 15700 9318
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 14740 8356 14792 8362
rect 14740 8298 14792 8304
rect 14752 8090 14780 8298
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14384 6934 14412 7482
rect 14568 7410 14596 7686
rect 14844 7546 14872 8434
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14016 6186 14044 6394
rect 14372 6316 14424 6322
rect 14648 6316 14700 6322
rect 14424 6276 14504 6304
rect 14372 6258 14424 6264
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 14476 5574 14504 6276
rect 14648 6258 14700 6264
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13740 4146 13768 4490
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13740 3602 13768 4082
rect 13832 4010 13860 5510
rect 14476 5370 14504 5510
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3670 13860 3946
rect 13820 3664 13872 3670
rect 13820 3606 13872 3612
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13096 3194 13124 3538
rect 14016 3194 14044 5170
rect 14660 5166 14688 6258
rect 15488 5846 15516 8230
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15580 6118 15608 6802
rect 15672 6390 15700 7210
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15396 5370 15424 5646
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14200 4826 14228 5034
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14660 4486 14688 5102
rect 15396 4826 15424 5306
rect 15488 5234 15516 5782
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15382 4720 15438 4729
rect 15382 4655 15384 4664
rect 15436 4655 15438 4664
rect 15384 4626 15436 4632
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15396 4282 15424 4626
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15580 4010 15608 6054
rect 15672 5710 15700 6326
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 4214 15700 5646
rect 15660 4208 15712 4214
rect 15764 4185 15792 7686
rect 15856 7546 15884 9658
rect 15948 7954 15976 10406
rect 16040 9722 16068 11562
rect 16224 11286 16252 12650
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11898 16528 12174
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16592 11762 16620 12786
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16684 11218 16712 12038
rect 17052 11354 17080 12174
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10470 16528 10950
rect 16684 10470 16712 11154
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 16040 8566 16068 9046
rect 16132 9042 16160 9998
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9518 16344 9862
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16132 8090 16160 8978
rect 16316 8294 16344 9454
rect 16684 8430 16712 10406
rect 16868 9042 16896 10542
rect 17144 10198 17172 13126
rect 17328 11014 17356 14010
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12442 17448 12582
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17420 11626 17448 12378
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17604 11218 17632 12242
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17604 10266 17632 11154
rect 17880 10470 17908 13942
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 18156 12986 18184 13398
rect 18616 13258 18644 22374
rect 18708 13394 18736 27526
rect 19248 27532 19300 27538
rect 19890 27532 19946 28000
rect 21362 27554 21418 28000
rect 19890 27520 19892 27532
rect 19248 27474 19300 27480
rect 19944 27520 19946 27532
rect 21100 27526 21418 27554
rect 19892 27474 19944 27480
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19076 23662 19104 24550
rect 19064 23656 19116 23662
rect 19064 23598 19116 23604
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 16182 18920 16390
rect 18880 16176 18932 16182
rect 18880 16118 18932 16124
rect 18984 16046 19012 16458
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18984 15162 19012 15982
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 19076 14521 19104 23598
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19168 16998 19196 17750
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 19168 16794 19196 16934
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19168 15706 19196 16730
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19260 15094 19288 27474
rect 19904 27443 19932 27474
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 21100 23866 21128 27526
rect 21362 27520 21418 27526
rect 22834 27520 22890 28000
rect 23860 27526 24256 27554
rect 22558 26752 22614 26761
rect 22558 26687 22614 26696
rect 21362 25528 21418 25537
rect 21362 25463 21418 25472
rect 21376 24274 21404 25463
rect 21364 24268 21416 24274
rect 21364 24210 21416 24216
rect 21376 23866 21404 24210
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21272 23588 21324 23594
rect 21272 23530 21324 23536
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19352 18426 19380 18770
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19904 18290 19932 18566
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19904 18068 19932 18226
rect 19904 18040 20024 18068
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17882 20024 18040
rect 20180 17882 20208 18226
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20180 17202 20208 17818
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19444 16250 19472 16662
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19444 15706 19472 15914
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20088 15706 20116 17002
rect 20180 16522 20208 17138
rect 20548 16726 20576 17206
rect 20536 16720 20588 16726
rect 20536 16662 20588 16668
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20732 15706 20760 16526
rect 21100 16250 21128 16662
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20168 15564 20220 15570
rect 20168 15506 20220 15512
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19062 14512 19118 14521
rect 18972 14476 19024 14482
rect 19062 14447 19118 14456
rect 18972 14418 19024 14424
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18604 13252 18656 13258
rect 18604 13194 18656 13200
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11830 18276 12038
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18156 11354 18184 11698
rect 18248 11626 18276 11766
rect 18432 11762 18460 13194
rect 18984 13172 19012 14418
rect 19536 14414 19564 15302
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14550 20024 14894
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 20180 14346 20208 15506
rect 21100 15502 21128 15914
rect 21180 15632 21232 15638
rect 21180 15574 21232 15580
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21192 15162 21220 15574
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13530 19472 13806
rect 20088 13802 20116 13874
rect 19892 13796 19944 13802
rect 20076 13796 20128 13802
rect 19944 13756 20024 13784
rect 19892 13738 19944 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19064 13184 19116 13190
rect 18984 13144 19064 13172
rect 19064 13126 19116 13132
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18616 12442 18644 12718
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18984 11558 19012 12242
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 17052 8838 17080 9454
rect 17144 9178 17172 10134
rect 17236 9518 17264 10134
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17684 9988 17736 9994
rect 17684 9930 17736 9936
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17420 9382 17448 9590
rect 17696 9586 17724 9930
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15948 7478 15976 7890
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 16132 7274 16160 7754
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16132 6934 16160 7210
rect 16120 6928 16172 6934
rect 16040 6888 16120 6916
rect 16040 5914 16068 6888
rect 16120 6870 16172 6876
rect 16316 6866 16344 7822
rect 16684 7750 16712 8366
rect 17052 8362 17080 8774
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17236 7886 17264 8774
rect 17420 8022 17448 9318
rect 17498 9072 17554 9081
rect 17498 9007 17554 9016
rect 17512 8566 17540 9007
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 6458 16344 6802
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16132 6186 16160 6394
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16040 4826 16068 5850
rect 16224 5574 16252 6258
rect 16684 6118 16712 6870
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15660 4150 15712 4156
rect 15750 4176 15806 4185
rect 15750 4111 15806 4120
rect 15764 4078 15792 4111
rect 16040 4078 16068 4762
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15568 4004 15620 4010
rect 15568 3946 15620 3952
rect 15382 3632 15438 3641
rect 15292 3596 15344 3602
rect 15344 3576 15382 3584
rect 15344 3567 15438 3576
rect 15344 3556 15424 3567
rect 15292 3538 15344 3544
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15396 3194 15424 3556
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 10414 82 10470 480
rect 10152 54 10470 82
rect 11440 82 11468 2246
rect 11794 82 11850 480
rect 11440 54 11850 82
rect 12912 82 12940 2790
rect 14200 2514 14228 2790
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 14200 2310 14228 2450
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 13174 82 13230 480
rect 12912 54 13230 82
rect 14384 82 14412 2314
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15580 1873 15608 3946
rect 15764 3738 15792 4014
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 16224 3670 16252 5510
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16316 4486 16344 5102
rect 16684 5098 16712 6054
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16776 4758 16804 6598
rect 16764 4752 16816 4758
rect 16764 4694 16816 4700
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16316 4146 16344 4422
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16408 3670 16436 4490
rect 16776 4282 16804 4694
rect 17144 4672 17172 7210
rect 17236 7002 17264 7822
rect 17420 7546 17448 7958
rect 17696 7886 17724 9522
rect 18156 9450 18184 10066
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17788 8634 17816 9046
rect 18248 8809 18276 10542
rect 18234 8800 18290 8809
rect 18156 8758 18234 8786
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 18156 8090 18184 8758
rect 18234 8735 18290 8744
rect 18326 8528 18382 8537
rect 18326 8463 18382 8472
rect 18340 8430 18368 8463
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18340 8090 18368 8366
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17788 6662 17816 7142
rect 18156 7002 18184 7346
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 18432 6254 18460 11494
rect 19076 11218 19104 13126
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 11694 19380 12582
rect 19444 12306 19472 13466
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19536 12714 19564 13330
rect 19706 13288 19762 13297
rect 19706 13223 19762 13232
rect 19720 13190 19748 13223
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11762 19472 12242
rect 19996 11762 20024 13756
rect 20076 13738 20128 13744
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 20088 12102 20116 12718
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19340 11688 19392 11694
rect 19260 11648 19340 11676
rect 19064 11212 19116 11218
rect 19064 11154 19116 11160
rect 19076 10538 19104 11154
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18524 8090 18552 8978
rect 18616 8430 18644 10474
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18800 9178 18828 9318
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18524 7002 18552 7822
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18616 6866 18644 8366
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18892 7206 18920 7958
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6322 18828 6598
rect 18984 6458 19012 10406
rect 19260 10198 19288 11648
rect 19340 11630 19392 11636
rect 19444 11218 19472 11698
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19996 11354 20024 11698
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 20088 11286 20116 12038
rect 20076 11280 20128 11286
rect 20076 11222 20128 11228
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19340 10532 19392 10538
rect 19340 10474 19392 10480
rect 19248 10192 19300 10198
rect 19248 10134 19300 10140
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19062 9616 19118 9625
rect 19062 9551 19118 9560
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 5914 18644 6190
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 18234 5808 18290 5817
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17236 5137 17264 5646
rect 17222 5128 17278 5137
rect 17222 5063 17278 5072
rect 17236 4826 17264 5063
rect 17328 5030 17356 5782
rect 19076 5778 19104 9551
rect 19168 9178 19196 9998
rect 19260 9722 19288 10134
rect 19352 9994 19380 10474
rect 19444 10198 19472 11154
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10538 19656 10950
rect 19616 10532 19668 10538
rect 19536 10492 19616 10520
rect 19536 10266 19564 10492
rect 19616 10474 19668 10480
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19260 9450 19288 9658
rect 19352 9586 19380 9930
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19156 9172 19208 9178
rect 19156 9114 19208 9120
rect 19536 8906 19564 9454
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19444 8430 19472 8774
rect 20088 8566 20116 8978
rect 20076 8560 20128 8566
rect 20076 8502 20128 8508
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19156 7268 19208 7274
rect 19904 7256 19932 7686
rect 19996 7546 20024 8434
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19984 7268 20036 7274
rect 19904 7228 19984 7256
rect 19156 7210 19208 7216
rect 19984 7210 20036 7216
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 19168 6798 19196 7210
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19536 7002 19564 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19168 5846 19196 6734
rect 19260 6390 19288 6870
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 18234 5743 18290 5752
rect 19064 5772 19116 5778
rect 18248 5710 18276 5743
rect 19064 5714 19116 5720
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 19076 5370 19104 5714
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17224 4684 17276 4690
rect 17144 4644 17224 4672
rect 17144 4282 17172 4644
rect 17224 4626 17276 4632
rect 17328 4486 17356 4966
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 17500 4616 17552 4622
rect 17500 4558 17552 4564
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16408 3505 16436 3606
rect 16394 3496 16450 3505
rect 16394 3431 16450 3440
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15566 1864 15622 1873
rect 15566 1799 15622 1808
rect 14646 82 14702 480
rect 14384 54 14702 82
rect 15672 82 15700 2246
rect 16026 82 16082 480
rect 15672 54 16082 82
rect 17144 82 17172 3878
rect 17236 3534 17264 3878
rect 17328 3670 17356 4422
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17236 3058 17264 3470
rect 17328 3194 17356 3606
rect 17512 3534 17540 4558
rect 17880 4282 17908 4694
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 18156 3058 18184 5034
rect 18800 4146 18828 5034
rect 19260 4826 19288 5714
rect 19444 5370 19472 6122
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19444 5098 19472 5306
rect 19536 5234 19564 5646
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19444 4758 19472 5034
rect 19536 4826 19564 5170
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18892 4282 18920 4422
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18800 2854 18828 3334
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18800 2009 18828 2790
rect 18786 2000 18842 2009
rect 18786 1935 18842 1944
rect 17406 82 17462 480
rect 17144 54 17462 82
rect 9034 0 9090 54
rect 10414 0 10470 54
rect 11794 0 11850 54
rect 13174 0 13230 54
rect 14646 0 14702 54
rect 16026 0 16082 54
rect 17406 0 17462 54
rect 18786 82 18842 480
rect 19076 82 19104 4626
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19444 4010 19472 4218
rect 19996 4214 20024 7210
rect 20088 7002 20116 7210
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 20180 6338 20208 14282
rect 20364 12850 20392 14826
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 13734 20852 14418
rect 20536 13728 20588 13734
rect 20536 13670 20588 13676
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20548 11898 20576 13670
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20456 9654 20484 10406
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 9178 20576 9318
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20640 8090 20668 8910
rect 20732 8838 20760 9998
rect 20824 9625 20852 13670
rect 20904 10192 20956 10198
rect 20904 10134 20956 10140
rect 20810 9616 20866 9625
rect 20810 9551 20866 9560
rect 20916 9450 20944 10134
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 21008 8956 21036 14962
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 14550 21128 14758
rect 21192 14618 21220 15098
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21100 14074 21128 14486
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21100 11354 21128 12174
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21088 11212 21140 11218
rect 21088 11154 21140 11160
rect 21100 10810 21128 11154
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21100 10577 21128 10746
rect 21086 10568 21142 10577
rect 21086 10503 21142 10512
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 21192 9654 21220 10474
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21284 9450 21312 23530
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 17066 21404 18090
rect 21560 17882 21588 24006
rect 22572 23866 22600 26687
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22008 23792 22060 23798
rect 22008 23734 22060 23740
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21560 17202 21588 17818
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21364 17060 21416 17066
rect 21364 17002 21416 17008
rect 21744 15638 21772 17206
rect 22020 16658 22048 23734
rect 22572 23662 22600 23802
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22848 23526 22876 27520
rect 22836 23520 22888 23526
rect 23860 23474 23888 27526
rect 24228 27520 24256 27526
rect 24306 27520 24362 28000
rect 24860 27532 24912 27538
rect 24228 27492 24348 27520
rect 25778 27532 25834 28000
rect 25778 27520 25780 27532
rect 24860 27474 24912 27480
rect 25832 27520 25834 27532
rect 26240 27532 26292 27538
rect 25780 27474 25832 27480
rect 27250 27532 27306 28000
rect 27250 27520 27252 27532
rect 26240 27474 26292 27480
rect 27304 27520 27306 27532
rect 27252 27474 27304 27480
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24766 24032 24822 24041
rect 24289 23964 24585 23984
rect 24766 23967 24822 23976
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 22836 23462 22888 23468
rect 23768 23446 23888 23474
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 17338 22508 17682
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21824 16176 21876 16182
rect 21824 16118 21876 16124
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21836 14822 21864 16118
rect 22204 15978 22232 17002
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22480 15910 22508 16594
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22480 15473 22508 15846
rect 22466 15464 22522 15473
rect 22466 15399 22522 15408
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21468 12986 21496 13398
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21652 12442 21680 14758
rect 22204 14550 22232 14894
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 13802 21864 14214
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21836 12918 21864 13738
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21824 12912 21876 12918
rect 21824 12854 21876 12860
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21364 12368 21416 12374
rect 21364 12310 21416 12316
rect 21376 11898 21404 12310
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 21284 9110 21312 9386
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 20824 8928 21036 8956
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20720 7336 20772 7342
rect 20088 6310 20208 6338
rect 20640 7296 20720 7324
rect 20088 4758 20116 6310
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20180 5914 20208 6190
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20088 4214 20116 4694
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 20076 4208 20128 4214
rect 20076 4150 20128 4156
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19260 3738 19288 3946
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 20640 3398 20668 7296
rect 20720 7278 20772 7284
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20732 5574 20760 6734
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20732 5234 20760 5510
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20824 3194 20852 8928
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 21008 8498 21036 8774
rect 21100 8634 21128 9046
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21284 8838 21312 8910
rect 21468 8906 21496 9318
rect 21560 8906 21588 10406
rect 21652 9722 21680 12378
rect 21928 12374 21956 13194
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 22020 10810 22048 13942
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22204 12170 22232 13738
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22296 13190 22324 13670
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22204 11014 22232 11698
rect 22296 11354 22324 13126
rect 22388 12850 22416 13126
rect 22480 12850 22508 13262
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22388 12442 22416 12786
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22376 11824 22428 11830
rect 22376 11766 22428 11772
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22388 11286 22416 11766
rect 22480 11762 22508 12786
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22376 11280 22428 11286
rect 22376 11222 22428 11228
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 21100 8022 21128 8570
rect 21652 8498 21680 9522
rect 21744 8974 21772 10474
rect 21836 10130 21864 10474
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 21824 9648 21876 9654
rect 21824 9590 21876 9596
rect 21836 9450 21864 9590
rect 21824 9444 21876 9450
rect 21824 9386 21876 9392
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21272 8492 21324 8498
rect 21640 8492 21692 8498
rect 21324 8452 21588 8480
rect 21272 8434 21324 8440
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21100 7478 21128 7958
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 21284 7206 21312 7822
rect 21560 7750 21588 8452
rect 21640 8434 21692 8440
rect 21652 8022 21680 8434
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21088 6928 21140 6934
rect 21088 6870 21140 6876
rect 21100 6390 21128 6870
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 21100 5370 21128 5782
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4282 20944 4966
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 20916 4010 20944 4218
rect 21008 4146 21036 4422
rect 20996 4140 21048 4146
rect 21048 4100 21128 4128
rect 20996 4082 21048 4088
rect 20904 4004 20956 4010
rect 20904 3946 20956 3952
rect 20994 3904 21050 3913
rect 20994 3839 21050 3848
rect 21008 3602 21036 3839
rect 21100 3738 21128 4100
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 21008 3194 21036 3538
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 21284 2650 21312 7142
rect 21744 6934 21772 7210
rect 21732 6928 21784 6934
rect 21732 6870 21784 6876
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21468 6254 21496 6666
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21744 5846 21772 6870
rect 21732 5840 21784 5846
rect 21732 5782 21784 5788
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21468 5302 21496 5646
rect 21456 5296 21508 5302
rect 21456 5238 21508 5244
rect 21468 4010 21496 5238
rect 21548 5092 21600 5098
rect 21548 5034 21600 5040
rect 21560 4690 21588 5034
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 21468 3534 21496 3946
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20088 2310 20116 2450
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 18786 54 19104 82
rect 20088 82 20116 2246
rect 20166 82 20222 480
rect 20088 54 20222 82
rect 21376 82 21404 2926
rect 21928 2650 21956 7686
rect 22020 6225 22048 10542
rect 22006 6216 22062 6225
rect 22006 6151 22062 6160
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 22204 2582 22232 10950
rect 22296 9926 22324 11018
rect 22388 10742 22416 11222
rect 22480 11150 22508 11698
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22376 10736 22428 10742
rect 22376 10678 22428 10684
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22296 2650 22324 9862
rect 22572 4154 22600 16050
rect 22756 15638 22784 16186
rect 22928 15972 22980 15978
rect 22928 15914 22980 15920
rect 22744 15632 22796 15638
rect 22796 15592 22876 15620
rect 22744 15574 22796 15580
rect 22744 15496 22796 15502
rect 22650 15464 22706 15473
rect 22744 15438 22796 15444
rect 22650 15399 22706 15408
rect 22664 14618 22692 15399
rect 22756 15026 22784 15438
rect 22848 15162 22876 15592
rect 22940 15502 22968 15914
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 23768 14618 23796 23446
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 24228 18222 24256 18770
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 18426 24808 23967
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24228 17338 24256 17682
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24766 16552 24822 16561
rect 24766 16487 24822 16496
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24780 15706 24808 16487
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24216 15564 24268 15570
rect 24216 15506 24268 15512
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24228 14822 24256 15506
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 24122 14512 24178 14521
rect 23480 14476 23532 14482
rect 24122 14447 24178 14456
rect 23480 14418 23532 14424
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22664 14074 22692 14282
rect 23492 14074 23520 14418
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23572 14000 23624 14006
rect 23478 13968 23534 13977
rect 23572 13942 23624 13948
rect 23478 13903 23534 13912
rect 22744 13864 22796 13870
rect 22664 13824 22744 13852
rect 22664 12646 22692 13824
rect 22744 13806 22796 13812
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22664 10690 22692 12582
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22848 11898 22876 12174
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22940 11694 22968 12310
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22836 11620 22888 11626
rect 22836 11562 22888 11568
rect 22848 10810 22876 11562
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22664 10662 22876 10690
rect 23032 10674 23060 11154
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22664 9722 22692 10202
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22756 9586 22784 9998
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22664 8634 22692 9046
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22848 7342 22876 10662
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22940 9994 22968 10202
rect 23032 10062 23060 10610
rect 23124 10606 23152 12718
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23400 10810 23428 11834
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23492 10690 23520 13903
rect 23584 13870 23612 13942
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24044 11898 24072 12174
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 24044 11626 24072 11834
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23400 10662 23520 10690
rect 23584 10674 23612 11154
rect 23572 10668 23624 10674
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23216 9625 23244 9862
rect 23202 9616 23258 9625
rect 23202 9551 23258 9560
rect 23308 9450 23336 9930
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 23308 9178 23336 9386
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23018 9072 23074 9081
rect 23018 9007 23074 9016
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22940 8634 22968 8910
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23032 8566 23060 9007
rect 23020 8560 23072 8566
rect 23308 8537 23336 9114
rect 23020 8502 23072 8508
rect 23294 8528 23350 8537
rect 23032 7954 23060 8502
rect 23294 8463 23350 8472
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23032 7546 23060 7890
rect 23400 7546 23428 10662
rect 23572 10610 23624 10616
rect 23584 9110 23612 10610
rect 24136 10606 24164 14447
rect 24228 13977 24256 14758
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24214 13968 24270 13977
rect 24214 13903 24270 13912
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12986 24716 13330
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24216 12368 24268 12374
rect 24216 12310 24268 12316
rect 24228 11898 24256 12310
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 15506
rect 24872 12986 24900 27474
rect 25792 27443 25820 27474
rect 25502 22944 25558 22953
rect 25502 22879 25558 22888
rect 25134 20360 25190 20369
rect 25134 20295 25190 20304
rect 25148 19514 25176 20295
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25148 19310 25176 19450
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25134 19136 25190 19145
rect 25134 19071 25190 19080
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24596 11354 24624 11630
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23846 8800 23902 8809
rect 23846 8735 23902 8744
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 22836 7336 22888 7342
rect 22836 7278 22888 7284
rect 22836 6452 22888 6458
rect 22836 6394 22888 6400
rect 22480 4126 22600 4154
rect 22480 3194 22508 4126
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 22848 2417 22876 6394
rect 23860 3641 23888 8735
rect 23952 7857 23980 9318
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 23938 7848 23994 7857
rect 23938 7783 23994 7792
rect 24044 7177 24072 8774
rect 24228 7313 24256 10406
rect 24768 10124 24820 10130
rect 24768 10066 24820 10072
rect 24780 9926 24808 10066
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24780 9722 24808 9862
rect 24768 9716 24820 9722
rect 24768 9658 24820 9664
rect 25148 9042 25176 19071
rect 25516 17882 25544 22879
rect 25504 17876 25556 17882
rect 25504 17818 25556 17824
rect 26252 13394 26280 27474
rect 27264 27443 27292 27474
rect 27618 22264 27674 22273
rect 27618 22199 27674 22208
rect 27632 15570 27660 22199
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27620 15088 27672 15094
rect 27620 15030 27672 15036
rect 27632 14657 27660 15030
rect 27618 14648 27674 14657
rect 27618 14583 27674 14592
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 25240 12617 25268 12650
rect 25226 12608 25282 12617
rect 25226 12543 25282 12552
rect 25778 10160 25834 10169
rect 25778 10095 25834 10104
rect 25792 9722 25820 10095
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25792 9518 25820 9658
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25136 9036 25188 9042
rect 25136 8978 25188 8984
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 25148 8634 25176 8978
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24214 7304 24270 7313
rect 24214 7239 24270 7248
rect 24030 7168 24086 7177
rect 24030 7103 24086 7112
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 27618 5672 27674 5681
rect 27618 5607 27674 5616
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 27632 4729 27660 5607
rect 27618 4720 27674 4729
rect 27618 4655 27674 4664
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23846 3632 23902 3641
rect 23846 3567 23902 3576
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 25412 2848 25464 2854
rect 25412 2790 25464 2796
rect 24216 2440 24268 2446
rect 22834 2408 22890 2417
rect 24216 2382 24268 2388
rect 22834 2343 22890 2352
rect 22652 2304 22704 2310
rect 22652 2246 22704 2252
rect 21638 82 21694 480
rect 21376 54 21694 82
rect 22664 82 22692 2246
rect 23018 82 23074 480
rect 22664 54 23074 82
rect 24228 82 24256 2382
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24398 82 24454 480
rect 24228 54 24454 82
rect 25424 82 25452 2790
rect 26884 2304 26936 2310
rect 26884 2246 26936 2252
rect 25778 82 25834 480
rect 25424 54 25834 82
rect 26896 82 26924 2246
rect 27158 82 27214 480
rect 26896 54 27214 82
rect 18786 0 18842 54
rect 20166 0 20222 54
rect 21638 0 21694 54
rect 23018 0 23074 54
rect 24398 0 24454 54
rect 25778 0 25834 54
rect 27158 0 27214 54
<< via2 >>
rect 110 24656 166 24712
rect 1122 25472 1178 25528
rect 110 19624 166 19680
rect 110 17040 166 17096
rect 110 13232 166 13288
rect 110 12008 166 12064
rect 110 10648 166 10704
rect 1674 22480 1730 22536
rect 1490 21664 1546 21720
rect 1582 20304 1638 20360
rect 1582 17992 1638 18048
rect 2226 26696 2282 26752
rect 110 8200 166 8256
rect 1582 8880 1638 8936
rect 110 4392 166 4448
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6550 23432 6606 23488
rect 6642 19216 6698 19272
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 4894 17176 4950 17232
rect 2226 6296 2282 6352
rect 1858 5208 1914 5264
rect 6366 18128 6422 18184
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5170 16496 5226 16552
rect 4894 16360 4950 16416
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6642 14320 6698 14376
rect 6550 13776 6606 13832
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 4986 10648 5042 10704
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 3974 6196 3976 6216
rect 3976 6196 4028 6216
rect 4028 6196 4030 6216
rect 3974 6160 4030 6196
rect 6918 12688 6974 12744
rect 6918 12144 6974 12200
rect 7286 13640 7342 13696
rect 6642 10512 6698 10568
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 2870 5072 2926 5128
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5446 3304 5502 3360
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5078 1808 5134 1864
rect 4894 1128 4950 1184
rect 7470 9968 7526 10024
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 12898 23704 12954 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 8666 16088 8722 16144
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 11794 17312 11850 17368
rect 7378 5072 7434 5128
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 13910 17176 13966 17232
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10046 14456 10102 14512
rect 9678 13640 9734 13696
rect 8850 10648 8906 10704
rect 9310 12144 9366 12200
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14646 17312 14702 17368
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14922 16088 14978 16144
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 9862 9288 9918 9344
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 8482 4140 8538 4176
rect 8482 4120 8484 4140
rect 8484 4120 8536 4140
rect 8536 4120 8538 4140
rect 8666 3440 8722 3496
rect 9034 4120 9090 4176
rect 9402 9016 9458 9072
rect 9954 9016 10010 9072
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 12530 9696 12586 9752
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10874 5752 10930 5808
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10138 4664 10194 4720
rect 7562 2352 7618 2408
rect 7562 1944 7618 2000
rect 6734 40 6790 96
rect 11886 7284 11888 7304
rect 11888 7284 11940 7304
rect 11940 7284 11942 7304
rect 11886 7248 11942 7284
rect 13542 11736 13598 11792
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 13818 10648 13874 10704
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 18050 22480 18106 22536
rect 16578 19216 16634 19272
rect 15658 13776 15714 13832
rect 16026 12688 16082 12744
rect 13726 9968 13782 10024
rect 14094 9968 14150 10024
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 13358 5208 13414 5264
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15382 4684 15438 4720
rect 15382 4664 15384 4684
rect 15384 4664 15436 4684
rect 15436 4664 15438 4684
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 22558 26696 22614 26752
rect 21362 25472 21418 25528
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19062 14456 19118 14512
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 17498 9016 17554 9072
rect 15750 4120 15806 4176
rect 15382 3576 15438 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 18234 8744 18290 8800
rect 18326 8472 18382 8528
rect 19706 13232 19762 13288
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19062 9560 19118 9616
rect 17222 5072 17278 5128
rect 18234 5752 18290 5808
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 16394 3440 16450 3496
rect 15566 1808 15622 1864
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 18786 1944 18842 2000
rect 20810 9560 20866 9616
rect 21086 10512 21142 10568
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 23976 24822 24032
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 22466 15408 22522 15464
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20994 3848 21050 3904
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22006 6160 22062 6216
rect 22650 15408 22706 15464
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 16496 24822 16552
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24122 14456 24178 14512
rect 23478 13912 23534 13968
rect 23202 9560 23258 9616
rect 23018 9016 23074 9072
rect 23294 8472 23350 8528
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24214 13912 24270 13968
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 25502 22888 25558 22944
rect 25134 20304 25190 20360
rect 25134 19080 25190 19136
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 23846 8744 23902 8800
rect 23938 7792 23994 7848
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 27618 22208 27674 22264
rect 27618 14592 27674 14648
rect 25226 12552 25282 12608
rect 25778 10104 25834 10160
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24214 7248 24270 7304
rect 24030 7112 24086 7168
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 27618 5616 27674 5672
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 27618 4664 27674 4720
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23846 3576 23902 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 22834 2352 22890 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
<< metal3 >>
rect 0 27208 480 27328
rect 27520 27208 28000 27328
rect 62 26754 122 27208
rect 2221 26754 2287 26757
rect 62 26752 2287 26754
rect 62 26696 2226 26752
rect 2282 26696 2287 26752
rect 62 26694 2287 26696
rect 2221 26691 2287 26694
rect 22553 26754 22619 26757
rect 27662 26754 27722 27208
rect 22553 26752 27722 26754
rect 22553 26696 22558 26752
rect 22614 26696 27722 26752
rect 22553 26694 27722 26696
rect 22553 26691 22619 26694
rect 0 25984 480 26104
rect 27520 25984 28000 26104
rect 62 25530 122 25984
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1117 25530 1183 25533
rect 62 25528 1183 25530
rect 62 25472 1122 25528
rect 1178 25472 1183 25528
rect 62 25470 1183 25472
rect 1117 25467 1183 25470
rect 21357 25530 21423 25533
rect 27662 25530 27722 25984
rect 21357 25528 27722 25530
rect 21357 25472 21362 25528
rect 21418 25472 27722 25528
rect 21357 25470 27722 25472
rect 21357 25467 21423 25470
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24712 480 24744
rect 0 24656 110 24712
rect 166 24656 480 24712
rect 0 24624 480 24656
rect 27520 24716 28000 24744
rect 27520 24652 27660 24716
rect 27724 24652 28000 24716
rect 27520 24624 28000 24652
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 24761 24034 24827 24037
rect 27654 24034 27660 24036
rect 24761 24032 27660 24034
rect 24761 23976 24766 24032
rect 24822 23976 27660 24032
rect 24761 23974 27660 23976
rect 24761 23971 24827 23974
rect 27654 23972 27660 23974
rect 27724 23972 27730 24036
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 12893 23762 12959 23765
rect 62 23760 12959 23762
rect 62 23704 12898 23760
rect 12954 23704 12959 23760
rect 62 23702 12959 23704
rect 62 23520 122 23702
rect 12893 23699 12959 23702
rect 0 23400 480 23520
rect 6545 23490 6611 23493
rect 6678 23490 6684 23492
rect 6545 23488 6684 23490
rect 6545 23432 6550 23488
rect 6606 23432 6684 23488
rect 6545 23430 6684 23432
rect 6545 23427 6611 23430
rect 6678 23428 6684 23430
rect 6748 23428 6754 23492
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 27520 23400 28000 23520
rect 19610 23359 19930 23360
rect 25497 22946 25563 22949
rect 27662 22946 27722 23400
rect 25497 22944 27722 22946
rect 25497 22888 25502 22944
rect 25558 22888 27722 22944
rect 25497 22886 27722 22888
rect 25497 22883 25563 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1669 22538 1735 22541
rect 18045 22538 18111 22541
rect 1669 22536 18111 22538
rect 1669 22480 1674 22536
rect 1730 22480 18050 22536
rect 18106 22480 18111 22536
rect 1669 22478 18111 22480
rect 1669 22475 1735 22478
rect 18045 22475 18111 22478
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 22264 28000 22296
rect 27520 22208 27618 22264
rect 27674 22208 28000 22264
rect 27520 22176 28000 22208
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1485 21722 1551 21725
rect 62 21720 1551 21722
rect 62 21664 1490 21720
rect 1546 21664 1551 21720
rect 62 21662 1551 21664
rect 1485 21659 1551 21662
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 0 20816 480 20936
rect 27520 20816 28000 20936
rect 62 20362 122 20816
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 1577 20362 1643 20365
rect 62 20360 1643 20362
rect 62 20304 1582 20360
rect 1638 20304 1643 20360
rect 62 20302 1643 20304
rect 1577 20299 1643 20302
rect 25129 20362 25195 20365
rect 27662 20362 27722 20816
rect 25129 20360 27722 20362
rect 25129 20304 25134 20360
rect 25190 20304 27722 20360
rect 25129 20302 27722 20304
rect 25129 20299 25195 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19680 480 19712
rect 0 19624 110 19680
rect 166 19624 480 19680
rect 0 19592 480 19624
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 27520 19592 28000 19712
rect 24277 19551 24597 19552
rect 6637 19274 6703 19277
rect 16573 19274 16639 19277
rect 6637 19272 16639 19274
rect 6637 19216 6642 19272
rect 6698 19216 16578 19272
rect 16634 19216 16639 19272
rect 6637 19214 16639 19216
rect 6637 19211 6703 19214
rect 16573 19211 16639 19214
rect 25129 19138 25195 19141
rect 27662 19138 27722 19592
rect 25129 19136 27722 19138
rect 25129 19080 25134 19136
rect 25190 19080 27722 19136
rect 25129 19078 27722 19080
rect 25129 19075 25195 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 5610 18528 5930 18529
rect 0 18368 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 27520 18368 28000 18488
rect 62 18050 122 18368
rect 6361 18186 6427 18189
rect 27662 18186 27722 18368
rect 6361 18184 27722 18186
rect 6361 18128 6366 18184
rect 6422 18128 27722 18184
rect 6361 18126 27722 18128
rect 6361 18123 6427 18126
rect 1577 18050 1643 18053
rect 62 18048 1643 18050
rect 62 17992 1582 18048
rect 1638 17992 1643 18048
rect 62 17990 1643 17992
rect 1577 17987 1643 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 11789 17370 11855 17373
rect 14641 17370 14707 17373
rect 11789 17368 14707 17370
rect 11789 17312 11794 17368
rect 11850 17312 14646 17368
rect 14702 17312 14707 17368
rect 11789 17310 14707 17312
rect 11789 17307 11855 17310
rect 14641 17307 14707 17310
rect 4889 17234 4955 17237
rect 13905 17234 13971 17237
rect 4889 17232 13971 17234
rect 4889 17176 4894 17232
rect 4950 17176 13910 17232
rect 13966 17176 13971 17232
rect 4889 17174 13971 17176
rect 4889 17171 4955 17174
rect 13905 17171 13971 17174
rect 0 17096 480 17128
rect 0 17040 110 17096
rect 166 17040 480 17096
rect 0 17008 480 17040
rect 27520 17008 28000 17128
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5165 16554 5231 16557
rect 10726 16554 10732 16556
rect 5165 16552 10732 16554
rect 5165 16496 5170 16552
rect 5226 16496 10732 16552
rect 5165 16494 10732 16496
rect 5165 16491 5231 16494
rect 10726 16492 10732 16494
rect 10796 16492 10802 16556
rect 24761 16554 24827 16557
rect 27662 16554 27722 17008
rect 24761 16552 27722 16554
rect 24761 16496 24766 16552
rect 24822 16496 27722 16552
rect 24761 16494 27722 16496
rect 24761 16491 24827 16494
rect 4889 16418 4955 16421
rect 62 16416 4955 16418
rect 62 16360 4894 16416
rect 4950 16360 4955 16416
rect 62 16358 4955 16360
rect 62 15904 122 16358
rect 4889 16355 4955 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 8661 16146 8727 16149
rect 14917 16146 14983 16149
rect 8661 16144 14983 16146
rect 8661 16088 8666 16144
rect 8722 16088 14922 16144
rect 14978 16088 14983 16144
rect 8661 16086 14983 16088
rect 8661 16083 8727 16086
rect 14917 16083 14983 16086
rect 0 15784 480 15904
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 27520 15784 28000 15904
rect 19610 15743 19930 15744
rect 10726 15404 10732 15468
rect 10796 15466 10802 15468
rect 22461 15466 22527 15469
rect 10796 15464 22527 15466
rect 10796 15408 22466 15464
rect 22522 15408 22527 15464
rect 10796 15406 22527 15408
rect 10796 15404 10802 15406
rect 22461 15403 22527 15406
rect 22645 15466 22711 15469
rect 27662 15466 27722 15784
rect 22645 15464 27722 15466
rect 22645 15408 22650 15464
rect 22706 15408 27722 15464
rect 22645 15406 27722 15408
rect 22645 15403 22711 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10277 14720 10597 14721
rect 0 14560 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 27520 14648 28000 14680
rect 27520 14592 27618 14648
rect 27674 14592 28000 14648
rect 27520 14560 28000 14592
rect 62 14378 122 14560
rect 10041 14514 10107 14517
rect 19057 14514 19123 14517
rect 24117 14514 24183 14517
rect 10041 14512 24183 14514
rect 10041 14456 10046 14512
rect 10102 14456 19062 14512
rect 19118 14456 24122 14512
rect 24178 14456 24183 14512
rect 10041 14454 24183 14456
rect 10041 14451 10107 14454
rect 19057 14451 19123 14454
rect 24117 14451 24183 14454
rect 6637 14378 6703 14381
rect 62 14376 6703 14378
rect 62 14320 6642 14376
rect 6698 14320 6703 14376
rect 62 14318 6703 14320
rect 6637 14315 6703 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 23473 13970 23539 13973
rect 24209 13970 24275 13973
rect 23473 13968 24275 13970
rect 23473 13912 23478 13968
rect 23534 13912 24214 13968
rect 24270 13912 24275 13968
rect 23473 13910 24275 13912
rect 23473 13907 23539 13910
rect 24209 13907 24275 13910
rect 6545 13834 6611 13837
rect 15653 13834 15719 13837
rect 6545 13832 15719 13834
rect 6545 13776 6550 13832
rect 6606 13776 15658 13832
rect 15714 13776 15719 13832
rect 6545 13774 15719 13776
rect 6545 13771 6611 13774
rect 15653 13771 15719 13774
rect 7281 13698 7347 13701
rect 9673 13698 9739 13701
rect 7281 13696 9739 13698
rect 7281 13640 7286 13696
rect 7342 13640 9678 13696
rect 9734 13640 9739 13696
rect 7281 13638 9739 13640
rect 7281 13635 7347 13638
rect 9673 13635 9739 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 0 13288 480 13320
rect 0 13232 110 13288
rect 166 13232 480 13288
rect 0 13200 480 13232
rect 19701 13290 19767 13293
rect 27520 13292 28000 13320
rect 27470 13290 27476 13292
rect 19701 13288 27476 13290
rect 19701 13232 19706 13288
rect 19762 13232 27476 13288
rect 19701 13230 27476 13232
rect 19701 13227 19767 13230
rect 27470 13228 27476 13230
rect 27540 13228 27660 13292
rect 27724 13228 28000 13292
rect 27520 13200 28000 13228
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6913 12746 6979 12749
rect 16021 12746 16087 12749
rect 6913 12744 16087 12746
rect 6913 12688 6918 12744
rect 6974 12688 16026 12744
rect 16082 12688 16087 12744
rect 6913 12686 16087 12688
rect 6913 12683 6979 12686
rect 16021 12683 16087 12686
rect 25221 12610 25287 12613
rect 25221 12608 27722 12610
rect 25221 12552 25226 12608
rect 25282 12552 27722 12608
rect 25221 12550 27722 12552
rect 25221 12547 25287 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 6913 12202 6979 12205
rect 9305 12202 9371 12205
rect 6913 12200 9371 12202
rect 6913 12144 6918 12200
rect 6974 12144 9310 12200
rect 9366 12144 9371 12200
rect 6913 12142 9371 12144
rect 6913 12139 6979 12142
rect 9305 12139 9371 12142
rect 27662 12096 27722 12550
rect 0 12064 480 12096
rect 0 12008 110 12064
rect 166 12008 480 12064
rect 0 11976 480 12008
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 27520 11976 28000 12096
rect 24277 11935 24597 11936
rect 6678 11732 6684 11796
rect 6748 11794 6754 11796
rect 13537 11794 13603 11797
rect 6748 11792 13603 11794
rect 6748 11736 13542 11792
rect 13598 11736 13603 11792
rect 6748 11734 13603 11736
rect 6748 11732 6754 11734
rect 13537 11731 13603 11734
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10704 480 10736
rect 0 10648 110 10704
rect 166 10648 480 10704
rect 0 10616 480 10648
rect 4981 10706 5047 10709
rect 8845 10706 8911 10709
rect 13813 10706 13879 10709
rect 4981 10704 13879 10706
rect 4981 10648 4986 10704
rect 5042 10648 8850 10704
rect 8906 10648 13818 10704
rect 13874 10648 13879 10704
rect 4981 10646 13879 10648
rect 4981 10643 5047 10646
rect 8845 10643 8911 10646
rect 13813 10643 13879 10646
rect 27520 10616 28000 10736
rect 6637 10570 6703 10573
rect 21081 10570 21147 10573
rect 6637 10568 21147 10570
rect 6637 10512 6642 10568
rect 6698 10512 21086 10568
rect 21142 10512 21147 10568
rect 6637 10510 21147 10512
rect 6637 10507 6703 10510
rect 21081 10507 21147 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 25773 10162 25839 10165
rect 27662 10162 27722 10616
rect 25773 10160 27722 10162
rect 25773 10104 25778 10160
rect 25834 10104 27722 10160
rect 25773 10102 27722 10104
rect 25773 10099 25839 10102
rect 7465 10026 7531 10029
rect 13721 10026 13787 10029
rect 14089 10026 14155 10029
rect 7465 10024 14155 10026
rect 7465 9968 7470 10024
rect 7526 9968 13726 10024
rect 13782 9968 14094 10024
rect 14150 9968 14155 10024
rect 7465 9966 14155 9968
rect 7465 9963 7531 9966
rect 13721 9963 13787 9966
rect 14089 9963 14155 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 12525 9754 12591 9757
rect 12750 9754 12756 9756
rect 12525 9752 12756 9754
rect 12525 9696 12530 9752
rect 12586 9696 12756 9752
rect 12525 9694 12756 9696
rect 12525 9691 12591 9694
rect 12750 9692 12756 9694
rect 12820 9692 12826 9756
rect 19057 9618 19123 9621
rect 20805 9618 20871 9621
rect 23197 9618 23263 9621
rect 19057 9616 23263 9618
rect 19057 9560 19062 9616
rect 19118 9560 20810 9616
rect 20866 9560 23202 9616
rect 23258 9560 23263 9616
rect 19057 9558 23263 9560
rect 19057 9555 19123 9558
rect 20805 9555 20871 9558
rect 23197 9555 23263 9558
rect 0 9392 480 9512
rect 27520 9392 28000 9512
rect 62 8938 122 9392
rect 9857 9346 9923 9349
rect 9990 9346 9996 9348
rect 9857 9344 9996 9346
rect 9857 9288 9862 9344
rect 9918 9288 9996 9344
rect 9857 9286 9996 9288
rect 9857 9283 9923 9286
rect 9990 9284 9996 9286
rect 10060 9284 10066 9348
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 9397 9074 9463 9077
rect 9949 9074 10015 9077
rect 17493 9074 17559 9077
rect 9397 9072 17559 9074
rect 9397 9016 9402 9072
rect 9458 9016 9954 9072
rect 10010 9016 17498 9072
rect 17554 9016 17559 9072
rect 9397 9014 17559 9016
rect 9397 9011 9463 9014
rect 9949 9011 10015 9014
rect 17493 9011 17559 9014
rect 23013 9074 23079 9077
rect 27662 9074 27722 9392
rect 23013 9072 27722 9074
rect 23013 9016 23018 9072
rect 23074 9016 27722 9072
rect 23013 9014 27722 9016
rect 23013 9011 23079 9014
rect 1577 8938 1643 8941
rect 62 8936 1643 8938
rect 62 8880 1582 8936
rect 1638 8880 1643 8936
rect 62 8878 1643 8880
rect 1577 8875 1643 8878
rect 18229 8802 18295 8805
rect 23841 8802 23907 8805
rect 18229 8800 23907 8802
rect 18229 8744 18234 8800
rect 18290 8744 23846 8800
rect 23902 8744 23907 8800
rect 18229 8742 23907 8744
rect 18229 8739 18295 8742
rect 23841 8739 23907 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 18321 8530 18387 8533
rect 23289 8530 23355 8533
rect 18321 8528 23355 8530
rect 18321 8472 18326 8528
rect 18382 8472 23294 8528
rect 23350 8472 23355 8528
rect 18321 8470 23355 8472
rect 18321 8467 18387 8470
rect 23289 8467 23355 8470
rect 0 8256 480 8288
rect 0 8200 110 8256
rect 166 8200 480 8256
rect 0 8168 480 8200
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8288
rect 19610 8127 19930 8128
rect 23422 7788 23428 7852
rect 23492 7850 23498 7852
rect 23933 7850 23999 7853
rect 23492 7848 23999 7850
rect 23492 7792 23938 7848
rect 23994 7792 23999 7848
rect 23492 7790 23999 7792
rect 23492 7788 23498 7790
rect 23933 7787 23999 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 11881 7306 11947 7309
rect 24209 7306 24275 7309
rect 27662 7306 27722 8168
rect 11881 7304 27722 7306
rect 11881 7248 11886 7304
rect 11942 7248 24214 7304
rect 24270 7248 27722 7304
rect 11881 7246 27722 7248
rect 11881 7243 11947 7246
rect 24209 7243 24275 7246
rect 23790 7108 23796 7172
rect 23860 7170 23866 7172
rect 24025 7170 24091 7173
rect 23860 7168 24091 7170
rect 23860 7112 24030 7168
rect 24086 7112 24091 7168
rect 23860 7110 24091 7112
rect 23860 7108 23866 7110
rect 24025 7107 24091 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6808 480 6928
rect 27520 6900 28000 6928
rect 27520 6836 27660 6900
rect 27724 6836 28000 6900
rect 27520 6808 28000 6836
rect 62 6354 122 6808
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 2221 6354 2287 6357
rect 62 6352 2287 6354
rect 62 6296 2226 6352
rect 2282 6296 2287 6352
rect 62 6294 2287 6296
rect 2221 6291 2287 6294
rect 3969 6218 4035 6221
rect 22001 6218 22067 6221
rect 3969 6216 22067 6218
rect 3969 6160 3974 6216
rect 4030 6160 22006 6216
rect 22062 6160 22067 6216
rect 3969 6158 22067 6160
rect 3969 6155 4035 6158
rect 22001 6155 22067 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 10869 5810 10935 5813
rect 18229 5810 18295 5813
rect 10869 5808 18295 5810
rect 10869 5752 10874 5808
rect 10930 5752 18234 5808
rect 18290 5752 18295 5808
rect 10869 5750 18295 5752
rect 10869 5747 10935 5750
rect 18229 5747 18295 5750
rect 0 5584 480 5704
rect 27520 5672 28000 5704
rect 27520 5616 27618 5672
rect 27674 5616 28000 5672
rect 27520 5584 28000 5616
rect 62 5266 122 5584
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 1853 5266 1919 5269
rect 13353 5266 13419 5269
rect 62 5264 1919 5266
rect 62 5208 1858 5264
rect 1914 5208 1919 5264
rect 62 5206 1919 5208
rect 1853 5203 1919 5206
rect 4110 5264 13419 5266
rect 4110 5208 13358 5264
rect 13414 5208 13419 5264
rect 4110 5206 13419 5208
rect 2865 5130 2931 5133
rect 4110 5130 4170 5206
rect 13353 5203 13419 5206
rect 2865 5128 4170 5130
rect 2865 5072 2870 5128
rect 2926 5072 4170 5128
rect 2865 5070 4170 5072
rect 7373 5130 7439 5133
rect 17217 5130 17283 5133
rect 7373 5128 17283 5130
rect 7373 5072 7378 5128
rect 7434 5072 17222 5128
rect 17278 5072 17283 5128
rect 7373 5070 17283 5072
rect 2865 5067 2931 5070
rect 7373 5067 7439 5070
rect 17217 5067 17283 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 10133 4722 10199 4725
rect 10726 4722 10732 4724
rect 10133 4720 10732 4722
rect 10133 4664 10138 4720
rect 10194 4664 10732 4720
rect 10133 4662 10732 4664
rect 10133 4659 10199 4662
rect 10726 4660 10732 4662
rect 10796 4660 10802 4724
rect 15377 4722 15443 4725
rect 27613 4722 27679 4725
rect 15377 4720 27679 4722
rect 15377 4664 15382 4720
rect 15438 4664 27618 4720
rect 27674 4664 27679 4720
rect 15377 4662 27679 4664
rect 15377 4659 15443 4662
rect 27613 4659 27679 4662
rect 0 4448 480 4480
rect 0 4392 110 4448
rect 166 4392 480 4448
rect 0 4360 480 4392
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4480
rect 24277 4319 24597 4320
rect 8477 4178 8543 4181
rect 9029 4178 9095 4181
rect 15745 4178 15811 4181
rect 8477 4176 15811 4178
rect 8477 4120 8482 4176
rect 8538 4120 9034 4176
rect 9090 4120 15750 4176
rect 15806 4120 15811 4176
rect 8477 4118 15811 4120
rect 8477 4115 8543 4118
rect 9029 4115 9095 4118
rect 15745 4115 15811 4118
rect 20989 3906 21055 3909
rect 27662 3906 27722 4360
rect 20989 3904 27722 3906
rect 20989 3848 20994 3904
rect 21050 3848 27722 3904
rect 20989 3846 27722 3848
rect 20989 3843 21055 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 27654 3770 27660 3772
rect 23430 3710 27660 3770
rect 15377 3634 15443 3637
rect 23430 3634 23490 3710
rect 27654 3708 27660 3710
rect 27724 3708 27730 3772
rect 15377 3632 23490 3634
rect 15377 3576 15382 3632
rect 15438 3576 23490 3632
rect 15377 3574 23490 3576
rect 23841 3634 23907 3637
rect 23841 3632 27722 3634
rect 23841 3576 23846 3632
rect 23902 3576 27722 3632
rect 23841 3574 27722 3576
rect 15377 3571 15443 3574
rect 23841 3571 23907 3574
rect 8661 3498 8727 3501
rect 16389 3498 16455 3501
rect 8661 3496 16455 3498
rect 8661 3440 8666 3496
rect 8722 3440 16394 3496
rect 16450 3440 16455 3496
rect 8661 3438 16455 3440
rect 8661 3435 8727 3438
rect 16389 3435 16455 3438
rect 5441 3362 5507 3365
rect 62 3360 5507 3362
rect 62 3304 5446 3360
rect 5502 3304 5507 3360
rect 62 3302 5507 3304
rect 62 3120 122 3302
rect 5441 3299 5507 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27662 3120 27722 3574
rect 0 3000 480 3120
rect 27520 3000 28000 3120
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 7557 2410 7623 2413
rect 62 2408 7623 2410
rect 62 2352 7562 2408
rect 7618 2352 7623 2408
rect 62 2350 7623 2352
rect 62 1896 122 2350
rect 7557 2347 7623 2350
rect 22829 2410 22895 2413
rect 22829 2408 27722 2410
rect 22829 2352 22834 2408
rect 22890 2352 27722 2408
rect 22829 2350 27722 2352
rect 22829 2347 22895 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 7557 2002 7623 2005
rect 18781 2002 18847 2005
rect 7557 2000 18847 2002
rect 7557 1944 7562 2000
rect 7618 1944 18786 2000
rect 18842 1944 18847 2000
rect 7557 1942 18847 1944
rect 7557 1939 7623 1942
rect 18781 1939 18847 1942
rect 27662 1896 27722 2350
rect 0 1776 480 1896
rect 5073 1866 5139 1869
rect 15561 1866 15627 1869
rect 5073 1864 15627 1866
rect 5073 1808 5078 1864
rect 5134 1808 15566 1864
rect 15622 1808 15627 1864
rect 5073 1806 15627 1808
rect 5073 1803 5139 1806
rect 15561 1803 15627 1806
rect 27520 1776 28000 1896
rect 4889 1186 4955 1189
rect 62 1184 4955 1186
rect 62 1128 4894 1184
rect 4950 1128 4955 1184
rect 62 1126 4955 1128
rect 62 672 122 1126
rect 4889 1123 4955 1126
rect 0 552 480 672
rect 27520 552 28000 672
rect 6729 98 6795 101
rect 27662 98 27722 552
rect 6729 96 27722 98
rect 6729 40 6734 96
rect 6790 40 27722 96
rect 6729 38 27722 40
rect 6729 35 6795 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 27660 24652 27724 24716
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 27660 23972 27724 24036
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 6684 23428 6748 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 10732 16492 10796 16556
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 10732 15404 10796 15468
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 27476 13228 27540 13292
rect 27660 13228 27724 13292
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 6684 11732 6748 11796
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 12756 9692 12820 9756
rect 9996 9284 10060 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 23428 7788 23492 7852
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 23796 7108 23860 7172
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 27660 6836 27724 6900
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 10732 4660 10796 4724
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 27660 3708 27724 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 6683 23492 6749 23493
rect 6683 23428 6684 23492
rect 6748 23428 6749 23492
rect 6683 23427 6749 23428
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 6686 11797 6746 23427
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 10731 16556 10797 16557
rect 10731 16492 10732 16556
rect 10796 16492 10797 16556
rect 10731 16491 10797 16492
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10734 15469 10794 16491
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 10731 15468 10797 15469
rect 10731 15404 10732 15468
rect 10796 15404 10797 15468
rect 10731 15403 10797 15404
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 6683 11796 6749 11797
rect 6683 11732 6684 11796
rect 6748 11732 6749 11796
rect 6683 11731 6749 11732
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9995 9348 10061 9349
rect 9995 9284 9996 9348
rect 10060 9284 10061 9348
rect 9995 9283 10061 9284
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 9998 7258 10058 9283
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10734 4725 10794 15403
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 12755 9756 12821 9757
rect 12755 9692 12756 9756
rect 12820 9692 12821 9756
rect 12755 9691 12821 9692
rect 12758 7938 12818 9691
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 10731 4724 10797 4725
rect 10731 4660 10732 4724
rect 10796 4660 10797 4724
rect 10731 4659 10797 4660
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 27659 24716 27725 24717
rect 27659 24652 27660 24716
rect 27724 24652 27725 24716
rect 27659 24651 27725 24652
rect 27662 24037 27722 24651
rect 27659 24036 27725 24037
rect 27659 23972 27660 24036
rect 27724 23972 27725 24036
rect 27659 23971 27725 23972
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 27475 13292 27541 13293
rect 27475 13228 27476 13292
rect 27540 13290 27541 13292
rect 27659 13292 27725 13293
rect 27659 13290 27660 13292
rect 27540 13230 27660 13290
rect 27540 13228 27541 13230
rect 27475 13227 27541 13228
rect 27659 13228 27660 13230
rect 27724 13228 27725 13292
rect 27659 13227 27725 13228
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 6560 24597 7584
rect 27659 6900 27725 6901
rect 27659 6836 27660 6900
rect 27724 6836 27725 6900
rect 27659 6835 27725 6836
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 27662 3773 27722 6835
rect 27659 3772 27725 3773
rect 27659 3708 27660 3772
rect 27724 3708 27725 3772
rect 27659 3707 27725 3708
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 9910 7022 10146 7258
rect 12670 7702 12906 7938
rect 23342 7852 23578 7938
rect 23342 7788 23428 7852
rect 23428 7788 23492 7852
rect 23492 7788 23578 7852
rect 23342 7702 23578 7788
rect 23710 7172 23946 7258
rect 23710 7108 23796 7172
rect 23796 7108 23860 7172
rect 23860 7108 23946 7172
rect 23710 7022 23946 7108
<< metal5 >>
rect 12628 7938 23620 7980
rect 12628 7702 12670 7938
rect 12906 7702 23342 7938
rect 23578 7702 23620 7938
rect 12628 7660 23620 7702
rect 9868 7258 23988 7300
rect 9868 7022 9910 7258
rect 10146 7022 23710 7258
rect 23946 7022 23988 7258
rect 9868 6980 23988 7022
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_1_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_34
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_46
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_68 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_71
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_63 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_72
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _178_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_85
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_83
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _084_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_96
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9844 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_100
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_139
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_139
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _186_
timestamp 1586364061
transform 1 0 13524 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_143
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_151
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_176
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_conb_1  _156_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_194
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_211
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_223
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_237
timestamp 1586364061
transform 1 0 22908 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_233
timestamp 1586364061
transform 1 0 22540 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_241
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_241
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_249
timestamp 1586364061
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23736 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_252
timestamp 1586364061
transform 1 0 24288 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_256
timestamp 1586364061
transform 1 0 24656 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_268
timestamp 1586364061
transform 1 0 25760 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_276
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 406 592
use scs8hd_or3_4  _089_
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_74
timestamp 1586364061
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 590 592
use scs8hd_conb_1  _155_
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_128
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_132
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_139
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 15732 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_157
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_161
timestamp 1586364061
transform 1 0 15916 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_183
timestamp 1586364061
transform 1 0 17940 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_191
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_230
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_242
timestamp 1586364061
transform 1 0 23368 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_254
timestamp 1586364061
transform 1 0 24472 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_decap_4  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_68
timestamp 1586364061
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_85
timestamp 1586364061
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _119_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_128
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_187
timestamp 1586364061
transform 1 0 18308 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_191
timestamp 1586364061
transform 1 0 18676 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_205
timestamp 1586364061
transform 1 0 19964 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_209
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_222
timestamp 1586364061
transform 1 0 21528 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_242
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_8  _058_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_139
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 15732 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_151
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_157
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_161
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_179
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_194
timestamp 1586364061
transform 1 0 18952 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_198
timestamp 1586364061
transform 1 0 19320 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_219
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_223
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_235
timestamp 1586364061
transform 1 0 22724 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_55
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_67
timestamp 1586364061
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _095_
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_131
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_148
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_213
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_230
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_6
timestamp 1586364061
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_17
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_10
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 314 592
use scs8hd_conb_1  _165_
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_21
timestamp 1586364061
transform 1 0 3036 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_28
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_40
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_36
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_40
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__C
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_50
timestamp 1586364061
transform 1 0 5704 0 -1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _073_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _060_
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_69
timestamp 1586364061
transform 1 0 7452 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_66
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _059_
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_76
timestamp 1586364061
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_80
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_97
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_90
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_101
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_99
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_139
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_147
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_143
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_155
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_168
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_176
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_173
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_1  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_183
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_194
timestamp 1586364061
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 18768 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 18124 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_198
timestamp 1586364061
transform 1 0 19320 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19688 0 1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_217
timestamp 1586364061
transform 1 0 21068 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_230
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_236
timestamp 1586364061
transform 1 0 22816 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_242
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_inv_8  _072_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_60
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _066_
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_73
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 590 592
use scs8hd_inv_8  _067_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_127
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_160
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_179
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_236
timestamp 1586364061
transform 1 0 22816 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_248
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _175_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_16
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_20
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__144__D
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_81
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_99
timestamp 1586364061
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_103
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_141
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_201
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_213
timestamp 1586364061
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_228
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_248
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_252
timestamp 1586364061
transform 1 0 24288 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_264
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _144_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_70
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 774 592
use scs8hd_or3_4  _130_
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_151
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_170
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_183
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_187
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_6  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_235
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_12
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_16
timestamp 1586364061
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _143_
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 1602 592
use scs8hd_buf_2  _177_
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_28
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_66
timestamp 1586364061
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_84
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _158_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_139
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_143
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_239
timestamp 1586364061
transform 1 0 23092 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_262
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_274
timestamp 1586364061
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_conb_1  _160_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_35
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _064_
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_39
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_52
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 406 592
use scs8hd_nor4_4  _137_
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_59
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_148
timestamp 1586364061
transform 1 0 14720 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_162
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_197
timestamp 1586364061
transform 1 0 19228 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_6  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_224
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_228
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 406 592
use scs8hd_conb_1  _167_
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_241
timestamp 1586364061
transform 1 0 23276 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_247
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_252
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _078_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_17
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_22
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_nor4_4  _149_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1602 592
use scs8hd_inv_8  _063_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _107_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_53
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_66
timestamp 1586364061
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__D
timestamp 1586364061
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _138_
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 1602 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _062_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__C
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_74
timestamp 1586364061
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_107
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_103
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_116
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use scs8hd_or2_4  _116_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 682 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13708 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_133
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_148
timestamp 1586364061
transform 1 0 14720 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_150
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 15364 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_164
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_182
timestamp 1586364061
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_226
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_243
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_260
timestamp 1586364061
transform 1 0 25024 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_272
timestamp 1586364061
transform 1 0 26128 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__D
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_29
timestamp 1586364061
transform 1 0 3772 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_34
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _108_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _139_
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_115
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_119
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 130 592
use scs8hd_or2_4  _087_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _085_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_212
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_252
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_259
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_275
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_11
timestamp 1586364061
transform 1 0 2116 0 -1 11424
box -38 -48 130 592
use scs8hd_nor4_4  _150_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__C
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_49
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_53
timestamp 1586364061
transform 1 0 5980 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 6164 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _061_
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__D
timestamp 1586364061
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__C
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_87
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _069_
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_138
timestamp 1586364061
transform 1 0 13800 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_194
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_204
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_222
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_226
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_250
timestamp 1586364061
transform 1 0 24104 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_262
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _172_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _079_
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 3956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_25
timestamp 1586364061
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_29
timestamp 1586364061
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _161_
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__D
timestamp 1586364061
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_47
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__C
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _140_
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 13340 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_129
timestamp 1586364061
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_142
timestamp 1586364061
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_250
timestamp 1586364061
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_2  _171_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_22
timestamp 1586364061
transform 1 0 3128 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _151_
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_62
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_66
timestamp 1586364061
transform 1 0 7176 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_81
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_85
timestamp 1586364061
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_108
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_119
timestamp 1586364061
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__C
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_165
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_184
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_188
timestamp 1586364061
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_205
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_208
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_8  FILLER_18_244
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_261
timestamp 1586364061
transform 1 0 25116 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_273
timestamp 1586364061
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_8  _082_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__D
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__D
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_nor4_4  _154_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1602 592
use scs8hd_nor4_4  _153_
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__C
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_44
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_48
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_52
timestamp 1586364061
transform 1 0 5888 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_71
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_75
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _123_
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_98
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__C
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_conb_1  _163_
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__D
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _148_
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1602 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__D
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__D
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_nor4_4  _152_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_127
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_195
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_20_204
timestamp 1586364061
transform 1 0 19872 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_202
timestamp 1586364061
transform 1 0 19688 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_212
timestamp 1586364061
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_244
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_20_252
timestamp 1586364061
transform 1 0 24288 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_258
timestamp 1586364061
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_270
timestamp 1586364061
transform 1 0 25944 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_274
timestamp 1586364061
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_12
timestamp 1586364061
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _141_
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 1602 592
use scs8hd_buf_2  _170_
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__142__D
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__C
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_24
timestamp 1586364061
transform 1 0 3312 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_21_60
timestamp 1586364061
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_88
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 314 592
use scs8hd_nor4_4  _147_
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _146_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_154
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_167
timestamp 1586364061
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 18952 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_190
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _168_
timestamp 1586364061
transform 1 0 20516 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_203
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_214
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_248
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_252
timestamp 1586364061
transform 1 0 24288 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_256
timestamp 1586364061
transform 1 0 24656 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_268
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_276
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_14
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _142_
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__C
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_18
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_49
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_67
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_71
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _145_
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1602 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_97
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_101
timestamp 1586364061
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_122
timestamp 1586364061
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_158
timestamp 1586364061
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_168
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_172
timestamp 1586364061
transform 1 0 16928 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 18952 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_185
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_193
timestamp 1586364061
transform 1 0 18860 0 -1 14688
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_203
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_207
timestamp 1586364061
transform 1 0 20148 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_211
timestamp 1586364061
transform 1 0 20516 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_228
timestamp 1586364061
transform 1 0 22080 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 23552 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_236
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_248
timestamp 1586364061
transform 1 0 23920 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_260
timestamp 1586364061
transform 1 0 25024 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_272
timestamp 1586364061
transform 1 0 26128 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _071_
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_26
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_44
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_79
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_83
timestamp 1586364061
transform 1 0 8740 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_116
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_151
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_195
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19964 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 21712 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_216
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_233
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_241
timestamp 1586364061
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 24380 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_43
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_47
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_50
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6624 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_75
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_104
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_108
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_123
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_127
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_131
timestamp 1586364061
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_24_157
timestamp 1586364061
transform 1 0 15548 0 -1 15776
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_161
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_164
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_183
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_24_186
timestamp 1586364061
transform 1 0 18216 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_225
timestamp 1586364061
transform 1 0 21804 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 1142 592
use scs8hd_buf_2  _179_
timestamp 1586364061
transform 1 0 24564 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_254
timestamp 1586364061
transform 1 0 24472 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_13
timestamp 1586364061
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_17
timestamp 1586364061
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_24
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_28
timestamp 1586364061
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_32
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_47
timestamp 1586364061
transform 1 0 5428 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_129
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_142
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_146
timestamp 1586364061
transform 1 0 14536 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_188
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_207
timestamp 1586364061
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_222
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_226
timestamp 1586364061
transform 1 0 21896 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_230
timestamp 1586364061
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_234
timestamp 1586364061
transform 1 0 22632 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_242
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_6
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_conb_1  _162_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_17
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_17
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_13
timestamp 1586364061
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 314 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 1472 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_25
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_25
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_28
timestamp 1586364061
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_78
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_88
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_84
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_85
timestamp 1586364061
transform 1 0 8924 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_81
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_105
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_101
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_104
timestamp 1586364061
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_112
timestamp 1586364061
transform 1 0 11408 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_108
timestamp 1586364061
transform 1 0 11040 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 1050 592
use scs8hd_inv_8  _077_
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_128
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 866 592
use scs8hd_or2_4  _100_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_149
timestamp 1586364061
transform 1 0 14812 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_166
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_177
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16652 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_187
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_184
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_194
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_191
timestamp 1586364061
transform 1 0 18676 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_198
timestamp 1586364061
transform 1 0 19320 0 1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_27_213
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_230
timestamp 1586364061
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_235
timestamp 1586364061
transform 1 0 22724 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_243
timestamp 1586364061
transform 1 0 23460 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 24288 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_259
timestamp 1586364061
transform 1 0 24932 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_251
timestamp 1586364061
transform 1 0 24196 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_266
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_271
timestamp 1586364061
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_274
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 314 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_28
timestamp 1586364061
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _070_
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_6  FILLER_28_49
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_63
timestamp 1586364061
transform 1 0 6900 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_75
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _159_
timestamp 1586364061
transform 1 0 11592 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_122
timestamp 1586364061
transform 1 0 12328 0 -1 17952
box -38 -48 314 592
use scs8hd_conb_1  _166_
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_134
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17204 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_171
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_209
timestamp 1586364061
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_28_223
timestamp 1586364061
transform 1 0 21620 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_231
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_236
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_248
timestamp 1586364061
transform 1 0 23920 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 24288 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_256
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_268
timestamp 1586364061
transform 1 0 25760 0 -1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_35
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 406 592
use scs8hd_conb_1  _164_
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_42
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_104
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_108
timestamp 1586364061
transform 1 0 11040 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_136
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_140
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_144
timestamp 1586364061
transform 1 0 14352 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_148
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_164
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_195
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_253
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_12
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_30_24
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4968 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_40
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12144 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_6  FILLER_30_114
timestamp 1586364061
transform 1 0 11592 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use scs8hd_conb_1  _169_
timestamp 1586364061
transform 1 0 17664 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_183
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_194
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_7
timestamp 1586364061
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_28
timestamp 1586364061
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_32
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_31_44
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _157_
timestamp 1586364061
transform 1 0 6900 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 130 592
use scs8hd_decap_6  FILLER_31_66
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 590 592
use scs8hd_buf_2  _183_
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 7728 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_78
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_89
timestamp 1586364061
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_93
timestamp 1586364061
transform 1 0 9660 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 590 592
use scs8hd_inv_8  _076_
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_144
timestamp 1586364061
transform 1 0 14352 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_180
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_253
timestamp 1586364061
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_262
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_274
timestamp 1586364061
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_62
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_6  FILLER_32_74
timestamp 1586364061
transform 1 0 7912 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_124
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_140
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_65
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_69
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_93
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_105
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_117
timestamp 1586364061
transform 1 0 11868 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_31
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_37_55
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 590 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_146
timestamp 1586364061
transform 1 0 14536 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_158
timestamp 1586364061
transform 1 0 15640 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_170
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_182
timestamp 1586364061
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_187
timestamp 1586364061
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_191
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_203
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_215
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_239
timestamp 1586364061
transform 1 0 23092 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_7
timestamp 1586364061
transform 1 0 1748 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_19
timestamp 1586364061
transform 1 0 2852 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_22
timestamp 1586364061
transform 1 0 3128 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_34
timestamp 1586364061
transform 1 0 4232 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_46
timestamp 1586364061
transform 1 0 5336 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _176_
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_39_80
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_85
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_89
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _174_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _173_
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_131
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_139
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_155
timestamp 1586364061
transform 1 0 15364 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_200
timestamp 1586364061
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_204
timestamp 1586364061
transform 1 0 19872 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_216
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_230
timestamp 1586364061
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_224
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_221
timestamp 1586364061
transform 1 0 21436 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_234
timestamp 1586364061
transform 1 0 22632 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_242
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_233
timestamp 1586364061
transform 1 0 22540 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_245
timestamp 1586364061
transform 1 0 23644 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_257
timestamp 1586364061
transform 1 0 24748 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_6  FILLER_40_269
timestamp 1586364061
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 552 480 672 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 1776 480 1896 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 3000 480 3120 6 address[2]
port 2 nsew default input
rlabel metal3 s 27520 552 28000 672 6 address[3]
port 3 nsew default input
rlabel metal2 s 754 27520 810 28000 6 address[4]
port 4 nsew default input
rlabel metal3 s 27520 1776 28000 1896 6 address[5]
port 5 nsew default input
rlabel metal3 s 27520 3000 28000 3120 6 address[6]
port 6 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 27520 6808 28000 6928 6 bottom_right_grid_pin_13_
port 9 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 bottom_right_grid_pin_15_
port 10 nsew default input
rlabel metal3 s 0 4360 480 4480 6 bottom_right_grid_pin_1_
port 11 nsew default input
rlabel metal3 s 0 5584 480 5704 6 bottom_right_grid_pin_3_
port 12 nsew default input
rlabel metal3 s 0 6808 480 6928 6 bottom_right_grid_pin_5_
port 13 nsew default input
rlabel metal3 s 27520 5584 28000 5704 6 bottom_right_grid_pin_7_
port 14 nsew default input
rlabel metal2 s 2226 27520 2282 28000 6 bottom_right_grid_pin_9_
port 15 nsew default input
rlabel metal2 s 4802 0 4858 480 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal2 s 5170 27520 5226 28000 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chanx_left_out[0]
port 25 nsew default tristate
rlabel metal3 s 0 8168 480 8288 6 chanx_left_out[1]
port 26 nsew default tristate
rlabel metal2 s 11058 27520 11114 28000 6 chanx_left_out[2]
port 27 nsew default tristate
rlabel metal3 s 0 9392 480 9512 6 chanx_left_out[3]
port 28 nsew default tristate
rlabel metal2 s 12530 27520 12586 28000 6 chanx_left_out[4]
port 29 nsew default tristate
rlabel metal2 s 14002 27520 14058 28000 6 chanx_left_out[5]
port 30 nsew default tristate
rlabel metal3 s 0 10616 480 10736 6 chanx_left_out[6]
port 31 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[7]
port 32 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[8]
port 33 nsew default tristate
rlabel metal2 s 15474 27520 15530 28000 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal3 s 27520 10616 28000 10736 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 16946 27520 17002 28000 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal3 s 27520 11976 28000 12096 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal3 s 27520 13200 28000 13320 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal3 s 0 20816 480 20936 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal3 s 27520 14560 28000 14680 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal3 s 27520 15784 28000 15904 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal3 s 27520 17008 28000 17128 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 16026 0 16082 480 6 chany_top_in[0]
port 52 nsew default input
rlabel metal3 s 27520 18368 28000 18488 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 18418 27520 18474 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal3 s 27520 19592 28000 19712 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 17406 0 17462 480 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 19890 27520 19946 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 18786 0 18842 480 6 chany_top_in[6]
port 58 nsew default input
rlabel metal3 s 0 22176 480 22296 6 chany_top_in[7]
port 59 nsew default input
rlabel metal3 s 27520 20816 28000 20936 6 chany_top_in[8]
port 60 nsew default input
rlabel metal3 s 27520 22176 28000 22296 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 22834 27520 22890 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal3 s 27520 24624 28000 24744 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 25778 27520 25834 28000 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 data_in
port 70 nsew default input
rlabel metal2 s 662 0 718 480 6 enable
port 71 nsew default input
rlabel metal3 s 0 25984 480 26104 6 left_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 0 27208 480 27328 6 left_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 20166 0 20222 480 6 top_left_grid_pin_13_
port 74 nsew default input
rlabel metal3 s 27520 27208 28000 27328 6 top_right_grid_pin_11_
port 75 nsew default input
rlabel metal2 s 25778 0 25834 480 6 top_right_grid_pin_13_
port 76 nsew default input
rlabel metal2 s 27158 0 27214 480 6 top_right_grid_pin_15_
port 77 nsew default input
rlabel metal2 s 21638 0 21694 480 6 top_right_grid_pin_1_
port 78 nsew default input
rlabel metal2 s 27250 27520 27306 28000 6 top_right_grid_pin_3_
port 79 nsew default input
rlabel metal2 s 23018 0 23074 480 6 top_right_grid_pin_5_
port 80 nsew default input
rlabel metal3 s 27520 25984 28000 26104 6 top_right_grid_pin_7_
port 81 nsew default input
rlabel metal2 s 24398 0 24454 480 6 top_right_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
