magic
tech sky130A
magscale 1 2
timestamp 1609023274
<< locali >>
rect 6871 5729 6963 5763
rect 6929 5627 6963 5729
<< viali >>
rect 4077 15113 4111 15147
rect 4721 15113 4755 15147
rect 5549 15113 5583 15147
rect 4353 15045 4387 15079
rect 4997 14977 5031 15011
rect 3893 14909 3927 14943
rect 4537 14909 4571 14943
rect 5365 14909 5399 14943
rect 5825 14773 5859 14807
rect 7481 14569 7515 14603
rect 9873 14569 9907 14603
rect 7297 14433 7331 14467
rect 9689 14433 9723 14467
rect 7757 14229 7791 14263
rect 10057 14229 10091 14263
rect 4169 14025 4203 14059
rect 4353 13821 4387 13855
rect 4609 13821 4643 13855
rect 5733 13685 5767 13719
rect 2789 13481 2823 13515
rect 4905 13481 4939 13515
rect 15485 13481 15519 13515
rect 2881 13345 2915 13379
rect 3249 13345 3283 13379
rect 5089 13345 5123 13379
rect 15301 13345 15335 13379
rect 3341 13141 3375 13175
rect 15025 13141 15059 13175
rect 7389 12393 7423 12427
rect 6101 12257 6135 12291
rect 7389 11645 7423 11679
rect 7634 11577 7668 11611
rect 7205 11509 7239 11543
rect 8769 11509 8803 11543
rect 7021 11305 7055 11339
rect 9229 11305 9263 11339
rect 9965 11237 9999 11271
rect 10241 11237 10275 11271
rect 7113 11169 7147 11203
rect 7757 11169 7791 11203
rect 8116 11169 8150 11203
rect 9321 11169 9355 11203
rect 7205 11101 7239 11135
rect 7849 11101 7883 11135
rect 6653 11033 6687 11067
rect 7573 11033 7607 11067
rect 3525 10761 3559 10795
rect 6653 10693 6687 10727
rect 3801 10625 3835 10659
rect 7389 10625 7423 10659
rect 7665 10625 7699 10659
rect 9781 10625 9815 10659
rect 10517 10625 10551 10659
rect 2932 10557 2966 10591
rect 7205 10557 7239 10591
rect 3019 10489 3053 10523
rect 3893 10489 3927 10523
rect 4813 10489 4847 10523
rect 7932 10489 7966 10523
rect 9597 10489 9631 10523
rect 10333 10489 10367 10523
rect 10793 10489 10827 10523
rect 6837 10421 6871 10455
rect 7297 10421 7331 10455
rect 9045 10421 9079 10455
rect 9137 10421 9171 10455
rect 9505 10421 9539 10455
rect 9965 10421 9999 10455
rect 10425 10421 10459 10455
rect 11069 10421 11103 10455
rect 10149 10217 10183 10251
rect 10793 10217 10827 10251
rect 1593 10149 1627 10183
rect 2513 10149 2547 10183
rect 6929 10081 6963 10115
rect 7389 10081 7423 10115
rect 7656 10081 7690 10115
rect 10057 10081 10091 10115
rect 1501 10013 1535 10047
rect 7021 10013 7055 10047
rect 7205 10013 7239 10047
rect 10241 10013 10275 10047
rect 6561 9877 6595 9911
rect 8769 9877 8803 9911
rect 9689 9877 9723 9911
rect 10609 9877 10643 9911
rect 7113 9673 7147 9707
rect 8125 9673 8159 9707
rect 7941 9605 7975 9639
rect 7573 9537 7607 9571
rect 7757 9537 7791 9571
rect 8677 9537 8711 9571
rect 9505 9537 9539 9571
rect 7481 9469 7515 9503
rect 8585 9469 8619 9503
rect 9413 9469 9447 9503
rect 8493 9401 8527 9435
rect 9321 9401 9355 9435
rect 1501 9333 1535 9367
rect 8953 9333 8987 9367
rect 9781 9333 9815 9367
rect 7021 9129 7055 9163
rect 6929 8993 6963 9027
rect 12633 8993 12667 9027
rect 7205 8925 7239 8959
rect 12817 8925 12851 8959
rect 6561 8789 6595 8823
rect 13553 8789 13587 8823
rect 3341 7293 3375 7327
rect 3617 7225 3651 7259
rect 7021 6409 7055 6443
rect 7849 6273 7883 6307
rect 7389 6205 7423 6239
rect 7941 5865 7975 5899
rect 9873 5865 9907 5899
rect 10885 5865 10919 5899
rect 11253 5865 11287 5899
rect 12265 5865 12299 5899
rect 12725 5865 12759 5899
rect 5089 5797 5123 5831
rect 5641 5797 5675 5831
rect 8861 5797 8895 5831
rect 4077 5729 4111 5763
rect 4445 5729 4479 5763
rect 5181 5729 5215 5763
rect 6561 5729 6595 5763
rect 6837 5729 6871 5763
rect 7021 5729 7055 5763
rect 7389 5729 7423 5763
rect 7757 5729 7791 5763
rect 8223 5729 8257 5763
rect 8677 5729 8711 5763
rect 9045 5729 9079 5763
rect 9413 5729 9447 5763
rect 9689 5729 9723 5763
rect 10057 5729 10091 5763
rect 10425 5729 10459 5763
rect 11621 5729 11655 5763
rect 12081 5729 12115 5763
rect 4813 5661 4847 5695
rect 12541 5661 12575 5695
rect 6745 5593 6779 5627
rect 6929 5593 6963 5627
rect 9229 5593 9263 5627
rect 11069 5593 11103 5627
rect 4261 5525 4295 5559
rect 4629 5525 4663 5559
rect 5365 5525 5399 5559
rect 7205 5525 7239 5559
rect 7573 5525 7607 5559
rect 8401 5525 8435 5559
rect 10241 5525 10275 5559
rect 10609 5525 10643 5559
rect 11805 5525 11839 5559
rect 5365 5321 5399 5355
rect 6009 5321 6043 5355
rect 7389 5321 7423 5355
rect 9321 5321 9355 5355
rect 9781 5321 9815 5355
rect 10241 5321 10275 5355
rect 10609 5321 10643 5355
rect 11069 5321 11103 5355
rect 13001 5321 13035 5355
rect 14013 5321 14047 5355
rect 11897 5253 11931 5287
rect 6653 5185 6687 5219
rect 12081 5185 12115 5219
rect 13645 5185 13679 5219
rect 4813 5117 4847 5151
rect 5181 5117 5215 5151
rect 5825 5117 5859 5151
rect 6193 5117 6227 5151
rect 6837 5117 6871 5151
rect 7205 5117 7239 5151
rect 7573 5117 7607 5151
rect 7941 5117 7975 5151
rect 8309 5117 8343 5151
rect 8677 5117 8711 5151
rect 9137 5117 9171 5151
rect 9597 5117 9631 5151
rect 10057 5117 10091 5151
rect 10425 5117 10459 5151
rect 10885 5117 10919 5151
rect 11253 5117 11287 5151
rect 11713 5117 11747 5151
rect 12449 5117 12483 5151
rect 12817 5117 12851 5151
rect 13185 5117 13219 5151
rect 4997 4981 5031 5015
rect 5641 4981 5675 5015
rect 6377 4981 6411 5015
rect 7021 4981 7055 5015
rect 7757 4981 7791 5015
rect 8125 4981 8159 5015
rect 8493 4981 8527 5015
rect 8861 4981 8895 5015
rect 11437 4981 11471 5015
rect 12633 4981 12667 5015
rect 13369 4981 13403 5015
rect 13829 4981 13863 5015
rect 9137 4777 9171 4811
rect 11621 4777 11655 4811
rect 8033 4641 8067 4675
rect 9229 4641 9263 4675
rect 10149 4641 10183 4675
rect 7665 4573 7699 4607
rect 9965 4573 9999 4607
rect 8769 4505 8803 4539
rect 10517 4505 10551 4539
rect 5273 4437 5307 4471
rect 6653 4437 6687 4471
rect 7297 4437 7331 4471
rect 8401 4437 8435 4471
rect 9413 4437 9447 4471
rect 9781 4437 9815 4471
rect 10885 4437 10919 4471
rect 12173 4437 12207 4471
<< metal1 >>
rect 5258 17892 5264 17944
rect 5316 17932 5322 17944
rect 5442 17932 5448 17944
rect 5316 17904 5448 17932
rect 5316 17892 5322 17904
rect 5442 17892 5448 17904
rect 5500 17892 5506 17944
rect 1104 17434 16008 17456
rect 1104 17382 3480 17434
rect 3532 17382 3544 17434
rect 3596 17382 3608 17434
rect 3660 17382 3672 17434
rect 3724 17382 8478 17434
rect 8530 17382 8542 17434
rect 8594 17382 8606 17434
rect 8658 17382 8670 17434
rect 8722 17382 13475 17434
rect 13527 17382 13539 17434
rect 13591 17382 13603 17434
rect 13655 17382 13667 17434
rect 13719 17382 16008 17434
rect 1104 17360 16008 17382
rect 1104 16890 16008 16912
rect 1104 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 10976 16890
rect 11028 16838 11040 16890
rect 11092 16838 11104 16890
rect 11156 16838 11168 16890
rect 11220 16838 16008 16890
rect 1104 16816 16008 16838
rect 7834 16532 7840 16584
rect 7892 16572 7898 16584
rect 10870 16572 10876 16584
rect 7892 16544 10876 16572
rect 7892 16532 7898 16544
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 1104 16346 16008 16368
rect 1104 16294 3480 16346
rect 3532 16294 3544 16346
rect 3596 16294 3608 16346
rect 3660 16294 3672 16346
rect 3724 16294 8478 16346
rect 8530 16294 8542 16346
rect 8594 16294 8606 16346
rect 8658 16294 8670 16346
rect 8722 16294 13475 16346
rect 13527 16294 13539 16346
rect 13591 16294 13603 16346
rect 13655 16294 13667 16346
rect 13719 16294 16008 16346
rect 1104 16272 16008 16294
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 10594 16096 10600 16108
rect 6512 16068 10600 16096
rect 6512 16056 6518 16068
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 9766 16028 9772 16040
rect 7156 16000 9772 16028
rect 7156 15988 7162 16000
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 9674 15960 9680 15972
rect 5684 15932 9680 15960
rect 5684 15920 5690 15932
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 13078 15920 13084 15972
rect 13136 15960 13142 15972
rect 15286 15960 15292 15972
rect 13136 15932 15292 15960
rect 13136 15920 13142 15932
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 3786 15852 3792 15904
rect 3844 15892 3850 15904
rect 3970 15892 3976 15904
rect 3844 15864 3976 15892
rect 3844 15852 3850 15864
rect 3970 15852 3976 15864
rect 4028 15852 4034 15904
rect 4338 15852 4344 15904
rect 4396 15892 4402 15904
rect 5350 15892 5356 15904
rect 4396 15864 5356 15892
rect 4396 15852 4402 15864
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 7742 15852 7748 15904
rect 7800 15892 7806 15904
rect 9766 15892 9772 15904
rect 7800 15864 9772 15892
rect 7800 15852 7806 15864
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 10134 15852 10140 15904
rect 10192 15892 10198 15904
rect 12342 15892 12348 15904
rect 10192 15864 12348 15892
rect 10192 15852 10198 15864
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 15654 15892 15660 15904
rect 13872 15864 15660 15892
rect 13872 15852 13878 15864
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 1104 15802 16008 15824
rect 1104 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 10976 15802
rect 11028 15750 11040 15802
rect 11092 15750 11104 15802
rect 11156 15750 11168 15802
rect 11220 15750 16008 15802
rect 1104 15728 16008 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 2682 15688 2688 15700
rect 1912 15660 2688 15688
rect 1912 15648 1918 15660
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3970 15688 3976 15700
rect 3108 15660 3976 15688
rect 3108 15648 3114 15660
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 13354 15688 13360 15700
rect 9088 15660 13360 15688
rect 9088 15648 9094 15660
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 9950 15620 9956 15632
rect 6328 15592 9956 15620
rect 6328 15580 6334 15592
rect 9950 15580 9956 15592
rect 10008 15580 10014 15632
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 13170 15620 13176 15632
rect 10836 15592 13176 15620
rect 10836 15580 10842 15592
rect 13170 15580 13176 15592
rect 13228 15580 13234 15632
rect 2222 15512 2228 15564
rect 2280 15552 2286 15564
rect 5534 15552 5540 15564
rect 2280 15524 5540 15552
rect 2280 15512 2286 15524
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 8846 15512 8852 15564
rect 8904 15552 8910 15564
rect 9398 15552 9404 15564
rect 8904 15524 9404 15552
rect 8904 15512 8910 15524
rect 9398 15512 9404 15524
rect 9456 15512 9462 15564
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 4706 15484 4712 15496
rect 1452 15456 4712 15484
rect 1452 15444 1458 15456
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 198 15376 204 15428
rect 256 15416 262 15428
rect 2866 15416 2872 15428
rect 256 15388 2872 15416
rect 256 15376 262 15388
rect 2866 15376 2872 15388
rect 2924 15376 2930 15428
rect 11974 15376 11980 15428
rect 12032 15416 12038 15428
rect 14458 15416 14464 15428
rect 12032 15388 14464 15416
rect 12032 15376 12038 15388
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 4798 15308 4804 15360
rect 4856 15348 4862 15360
rect 6730 15348 6736 15360
rect 4856 15320 6736 15348
rect 4856 15308 4862 15320
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 7282 15308 7288 15360
rect 7340 15348 7346 15360
rect 9582 15348 9588 15360
rect 7340 15320 9588 15348
rect 7340 15308 7346 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12710 15348 12716 15360
rect 11756 15320 12716 15348
rect 11756 15308 11762 15320
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 1104 15258 16008 15280
rect 1104 15206 3480 15258
rect 3532 15206 3544 15258
rect 3596 15206 3608 15258
rect 3660 15206 3672 15258
rect 3724 15206 8478 15258
rect 8530 15206 8542 15258
rect 8594 15206 8606 15258
rect 8658 15206 8670 15258
rect 8722 15206 13475 15258
rect 13527 15206 13539 15258
rect 13591 15206 13603 15258
rect 13655 15206 13667 15258
rect 13719 15206 16008 15258
rect 1104 15184 16008 15206
rect 566 15104 572 15156
rect 624 15144 630 15156
rect 4065 15147 4123 15153
rect 4065 15144 4077 15147
rect 624 15116 4077 15144
rect 624 15104 630 15116
rect 4065 15113 4077 15116
rect 4111 15113 4123 15147
rect 4706 15144 4712 15156
rect 4667 15116 4712 15144
rect 4065 15107 4123 15113
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 4341 15079 4399 15085
rect 4341 15045 4353 15079
rect 4387 15076 4399 15079
rect 7190 15076 7196 15088
rect 4387 15048 7196 15076
rect 4387 15045 4399 15048
rect 4341 15039 4399 15045
rect 3881 14943 3939 14949
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 4356 14940 4384 15039
rect 7190 15036 7196 15048
rect 7248 15036 7254 15088
rect 4985 15011 5043 15017
rect 4985 15008 4997 15011
rect 4540 14980 4997 15008
rect 4540 14949 4568 14980
rect 4985 14977 4997 14980
rect 5031 15008 5043 15011
rect 5534 15008 5540 15020
rect 5031 14980 5540 15008
rect 5031 14977 5043 14980
rect 4985 14971 5043 14977
rect 5534 14968 5540 14980
rect 5592 14968 5598 15020
rect 3927 14912 4384 14940
rect 4525 14943 4583 14949
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14909 5411 14943
rect 5353 14903 5411 14909
rect 5368 14804 5396 14903
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 5368 14776 5825 14804
rect 5813 14773 5825 14776
rect 5859 14804 5871 14807
rect 9858 14804 9864 14816
rect 5859 14776 9864 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 1104 14714 16008 14736
rect 1104 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 10976 14714
rect 11028 14662 11040 14714
rect 11092 14662 11104 14714
rect 11156 14662 11168 14714
rect 11220 14662 16008 14714
rect 1104 14640 16008 14662
rect 6730 14560 6736 14612
rect 6788 14600 6794 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 6788 14572 7481 14600
rect 6788 14560 6794 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 9640 14572 9873 14600
rect 9640 14560 9646 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 9861 14563 9919 14569
rect 7285 14467 7343 14473
rect 7285 14433 7297 14467
rect 7331 14464 7343 14467
rect 9677 14467 9735 14473
rect 7331 14436 7788 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 7760 14269 7788 14436
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 10042 14464 10048 14476
rect 9723 14436 10048 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 11514 14424 11520 14476
rect 11572 14464 11578 14476
rect 14826 14464 14832 14476
rect 11572 14436 14832 14464
rect 11572 14424 11578 14436
rect 14826 14424 14832 14436
rect 14884 14424 14890 14476
rect 7745 14263 7803 14269
rect 7745 14229 7757 14263
rect 7791 14260 7803 14263
rect 8846 14260 8852 14272
rect 7791 14232 8852 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 1104 14170 16008 14192
rect 1104 14118 3480 14170
rect 3532 14118 3544 14170
rect 3596 14118 3608 14170
rect 3660 14118 3672 14170
rect 3724 14118 8478 14170
rect 8530 14118 8542 14170
rect 8594 14118 8606 14170
rect 8658 14118 8670 14170
rect 8722 14118 13475 14170
rect 13527 14118 13539 14170
rect 13591 14118 13603 14170
rect 13655 14118 13667 14170
rect 13719 14118 16008 14170
rect 1104 14096 16008 14118
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 4120 14028 4169 14056
rect 4120 14016 4126 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4157 14019 4215 14025
rect 4172 13920 4200 14019
rect 4172 13892 4476 13920
rect 4338 13852 4344 13864
rect 4299 13824 4344 13852
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 4448 13852 4476 13892
rect 4597 13855 4655 13861
rect 4597 13852 4609 13855
rect 4448 13824 4609 13852
rect 4597 13821 4609 13824
rect 4643 13821 4655 13855
rect 4597 13815 4655 13821
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 1104 13626 16008 13648
rect 1104 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 10976 13626
rect 11028 13574 11040 13626
rect 11092 13574 11104 13626
rect 11156 13574 11168 13626
rect 11220 13574 16008 13626
rect 1104 13552 16008 13574
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 2866 13512 2872 13524
rect 2823 13484 2872 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4396 13484 4905 13512
rect 4396 13472 4402 13484
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 15470 13512 15476 13524
rect 15431 13484 15476 13512
rect 4893 13475 4951 13481
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 2884 13385 2912 13472
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13345 3295 13379
rect 3237 13339 3295 13345
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13376 5135 13379
rect 6270 13376 6276 13388
rect 5123 13348 6276 13376
rect 5123 13345 5135 13348
rect 5077 13339 5135 13345
rect 3252 13308 3280 13339
rect 6270 13336 6276 13348
rect 6328 13336 6334 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 15028 13348 15301 13376
rect 9306 13308 9312 13320
rect 3252 13280 9312 13308
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 3329 13175 3387 13181
rect 3329 13172 3341 13175
rect 3292 13144 3341 13172
rect 3292 13132 3298 13144
rect 3329 13141 3341 13144
rect 3375 13141 3387 13175
rect 3329 13135 3387 13141
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 15028 13181 15056 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14516 13144 15025 13172
rect 14516 13132 14522 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15013 13135 15071 13141
rect 1104 13082 16008 13104
rect 1104 13030 3480 13082
rect 3532 13030 3544 13082
rect 3596 13030 3608 13082
rect 3660 13030 3672 13082
rect 3724 13030 8478 13082
rect 8530 13030 8542 13082
rect 8594 13030 8606 13082
rect 8658 13030 8670 13082
rect 8722 13030 13475 13082
rect 13527 13030 13539 13082
rect 13591 13030 13603 13082
rect 13655 13030 13667 13082
rect 13719 13030 16008 13082
rect 1104 13008 16008 13030
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 13722 12628 13728 12640
rect 9364 12600 13728 12628
rect 9364 12588 9370 12600
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 1104 12538 16008 12560
rect 1104 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 10976 12538
rect 11028 12486 11040 12538
rect 11092 12486 11104 12538
rect 11156 12486 11168 12538
rect 11220 12486 16008 12538
rect 1104 12464 16008 12486
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6730 12424 6736 12436
rect 6328 12396 6736 12424
rect 6328 12384 6334 12396
rect 6730 12384 6736 12396
rect 6788 12424 6794 12436
rect 7377 12427 7435 12433
rect 7377 12424 7389 12427
rect 6788 12396 7389 12424
rect 6788 12384 6794 12396
rect 7377 12393 7389 12396
rect 7423 12393 7435 12427
rect 7377 12387 7435 12393
rect 11422 12384 11428 12436
rect 11480 12424 11486 12436
rect 11606 12424 11612 12436
rect 11480 12396 11612 12424
rect 11480 12384 11486 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 11330 12288 11336 12300
rect 6135 12260 11336 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 1104 11994 16008 12016
rect 1104 11942 3480 11994
rect 3532 11942 3544 11994
rect 3596 11942 3608 11994
rect 3660 11942 3672 11994
rect 3724 11942 8478 11994
rect 8530 11942 8542 11994
rect 8594 11942 8606 11994
rect 8658 11942 8670 11994
rect 8722 11942 13475 11994
rect 13527 11942 13539 11994
rect 13591 11942 13603 11994
rect 13655 11942 13667 11994
rect 13719 11942 16008 11994
rect 1104 11920 16008 11942
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 16942 11744 16948 11756
rect 15620 11716 16948 11744
rect 15620 11704 15626 11716
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11676 7435 11679
rect 7466 11676 7472 11688
rect 7423 11648 7472 11676
rect 7423 11645 7435 11648
rect 7377 11639 7435 11645
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 16482 11676 16488 11688
rect 15436 11648 16488 11676
rect 15436 11636 15442 11648
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 7282 11608 7288 11620
rect 5776 11580 7288 11608
rect 5776 11568 5782 11580
rect 7282 11568 7288 11580
rect 7340 11608 7346 11620
rect 7622 11611 7680 11617
rect 7622 11608 7634 11611
rect 7340 11580 7634 11608
rect 7340 11568 7346 11580
rect 7622 11577 7634 11580
rect 7668 11577 7680 11611
rect 7622 11571 7680 11577
rect 7190 11540 7196 11552
rect 7103 11512 7196 11540
rect 7190 11500 7196 11512
rect 7248 11540 7254 11552
rect 7466 11540 7472 11552
rect 7248 11512 7472 11540
rect 7248 11500 7254 11512
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 8352 11512 8769 11540
rect 8352 11500 8358 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 1104 11450 16008 11472
rect 1104 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 10976 11450
rect 11028 11398 11040 11450
rect 11092 11398 11104 11450
rect 11156 11398 11168 11450
rect 11220 11398 16008 11450
rect 1104 11376 16008 11398
rect 7009 11339 7067 11345
rect 7009 11305 7021 11339
rect 7055 11336 7067 11339
rect 9217 11339 9275 11345
rect 7055 11308 7972 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 7944 11268 7972 11308
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9306 11336 9312 11348
rect 9263 11308 9312 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 8938 11268 8944 11280
rect 6788 11240 7512 11268
rect 7944 11240 8944 11268
rect 6788 11228 6794 11240
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 7374 11200 7380 11212
rect 7147 11172 7380 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 7374 11160 7380 11172
rect 7432 11160 7438 11212
rect 7484 11200 7512 11240
rect 8938 11228 8944 11240
rect 8996 11268 9002 11280
rect 8996 11240 9352 11268
rect 8996 11228 9002 11240
rect 9324 11212 9352 11240
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 9953 11271 10011 11277
rect 9953 11268 9965 11271
rect 9916 11240 9965 11268
rect 9916 11228 9922 11240
rect 9953 11237 9965 11240
rect 9999 11237 10011 11271
rect 9953 11231 10011 11237
rect 10229 11271 10287 11277
rect 10229 11237 10241 11271
rect 10275 11268 10287 11271
rect 10686 11268 10692 11280
rect 10275 11240 10692 11268
rect 10275 11237 10287 11240
rect 10229 11231 10287 11237
rect 8110 11209 8116 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7484 11172 7757 11200
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 8104 11200 8116 11209
rect 8071 11172 8116 11200
rect 7745 11163 7803 11169
rect 8104 11163 8116 11172
rect 8110 11160 8116 11163
rect 8168 11160 8174 11212
rect 9306 11200 9312 11212
rect 9267 11172 9312 11200
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 6641 11067 6699 11073
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 7006 11064 7012 11076
rect 6687 11036 7012 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7208 10996 7236 11095
rect 7558 11064 7564 11076
rect 7519 11036 7564 11064
rect 7558 11024 7564 11036
rect 7616 11064 7622 11076
rect 7852 11064 7880 11095
rect 7616 11036 7880 11064
rect 7616 11024 7622 11036
rect 7282 10996 7288 11008
rect 7208 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 9490 10956 9496 11008
rect 9548 10996 9554 11008
rect 10244 10996 10272 11231
rect 10686 11228 10692 11240
rect 10744 11228 10750 11280
rect 9548 10968 10272 10996
rect 9548 10956 9554 10968
rect 1104 10906 16008 10928
rect 1104 10854 3480 10906
rect 3532 10854 3544 10906
rect 3596 10854 3608 10906
rect 3660 10854 3672 10906
rect 3724 10854 8478 10906
rect 8530 10854 8542 10906
rect 8594 10854 8606 10906
rect 8658 10854 8670 10906
rect 8722 10854 13475 10906
rect 13527 10854 13539 10906
rect 13591 10854 13603 10906
rect 13655 10854 13667 10906
rect 13719 10854 16008 10906
rect 1104 10832 16008 10854
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3384 10764 3525 10792
rect 3384 10752 3390 10764
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 3513 10755 3571 10761
rect 7392 10764 8708 10792
rect 3528 10656 3556 10755
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 6641 10727 6699 10733
rect 6641 10724 6653 10727
rect 5592 10696 6653 10724
rect 5592 10684 5598 10696
rect 6641 10693 6653 10696
rect 6687 10724 6699 10727
rect 7190 10724 7196 10736
rect 6687 10696 7196 10724
rect 6687 10693 6699 10696
rect 6641 10687 6699 10693
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3528 10628 3801 10656
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7392 10665 7420 10764
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7340 10628 7389 10656
rect 7340 10616 7346 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7616 10628 7665 10656
rect 7616 10616 7622 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 8680 10656 8708 10764
rect 10870 10752 10876 10804
rect 10928 10792 10934 10804
rect 13814 10792 13820 10804
rect 10928 10764 13820 10792
rect 10928 10752 10934 10764
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 8680 10628 9781 10656
rect 7653 10619 7711 10625
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 10042 10616 10048 10668
rect 10100 10656 10106 10668
rect 10318 10656 10324 10668
rect 10100 10628 10324 10656
rect 10100 10616 10106 10628
rect 10318 10616 10324 10628
rect 10376 10616 10382 10668
rect 10502 10656 10508 10668
rect 10463 10628 10508 10656
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 2920 10591 2978 10597
rect 2920 10588 2932 10591
rect 1544 10560 2932 10588
rect 1544 10548 1550 10560
rect 2920 10557 2932 10560
rect 2966 10588 2978 10591
rect 3234 10588 3240 10600
rect 2966 10560 3240 10588
rect 2966 10557 2978 10560
rect 2920 10551 2978 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 7156 10560 7205 10588
rect 7156 10548 7162 10560
rect 7193 10557 7205 10560
rect 7239 10588 7251 10591
rect 7466 10588 7472 10600
rect 7239 10560 7472 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7466 10548 7472 10560
rect 7524 10548 7530 10600
rect 7852 10560 12296 10588
rect 3007 10523 3065 10529
rect 3007 10489 3019 10523
rect 3053 10520 3065 10523
rect 3881 10523 3939 10529
rect 3053 10492 3740 10520
rect 3053 10489 3065 10492
rect 3007 10483 3065 10489
rect 3712 10452 3740 10492
rect 3881 10489 3893 10523
rect 3927 10489 3939 10523
rect 3881 10483 3939 10489
rect 4801 10523 4859 10529
rect 4801 10489 4813 10523
rect 4847 10520 4859 10523
rect 7852 10520 7880 10560
rect 4847 10492 7880 10520
rect 7920 10523 7978 10529
rect 4847 10489 4859 10492
rect 4801 10483 4859 10489
rect 7920 10489 7932 10523
rect 7966 10520 7978 10523
rect 8294 10520 8300 10532
rect 7966 10492 8300 10520
rect 7966 10489 7978 10492
rect 7920 10483 7978 10489
rect 3896 10452 3924 10483
rect 8294 10480 8300 10492
rect 8352 10480 8358 10532
rect 9585 10523 9643 10529
rect 9585 10489 9597 10523
rect 9631 10520 9643 10523
rect 9858 10520 9864 10532
rect 9631 10492 9864 10520
rect 9631 10489 9643 10492
rect 9585 10483 9643 10489
rect 9858 10480 9864 10492
rect 9916 10520 9922 10532
rect 10226 10520 10232 10532
rect 9916 10492 10232 10520
rect 9916 10480 9922 10492
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10321 10523 10379 10529
rect 10321 10489 10333 10523
rect 10367 10520 10379 10523
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 10367 10492 10793 10520
rect 10367 10489 10379 10492
rect 10321 10483 10379 10489
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 12268 10520 12296 10560
rect 14458 10520 14464 10532
rect 12268 10492 14464 10520
rect 10781 10483 10839 10489
rect 14458 10480 14464 10492
rect 14516 10480 14522 10532
rect 3712 10424 3924 10452
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 7098 10452 7104 10464
rect 6871 10424 7104 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 7248 10424 7297 10452
rect 7248 10412 7254 10424
rect 7285 10421 7297 10424
rect 7331 10452 7343 10455
rect 8386 10452 8392 10464
rect 7331 10424 8392 10452
rect 7331 10421 7343 10424
rect 7285 10415 7343 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 9030 10452 9036 10464
rect 8991 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9490 10452 9496 10464
rect 9180 10424 9225 10452
rect 9451 10424 9496 10452
rect 9180 10412 9186 10424
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9950 10452 9956 10464
rect 9911 10424 9956 10452
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10410 10452 10416 10464
rect 10371 10424 10416 10452
rect 10410 10412 10416 10424
rect 10468 10452 10474 10464
rect 10870 10452 10876 10464
rect 10468 10424 10876 10452
rect 10468 10412 10474 10424
rect 10870 10412 10876 10424
rect 10928 10452 10934 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 10928 10424 11069 10452
rect 10928 10412 10934 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 11057 10415 11115 10421
rect 1104 10362 16008 10384
rect 1104 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 10976 10362
rect 11028 10310 11040 10362
rect 11092 10310 11104 10362
rect 11156 10310 11168 10362
rect 11220 10310 16008 10362
rect 1104 10288 16008 10310
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7558 10248 7564 10260
rect 7064 10220 7564 10248
rect 7064 10208 7070 10220
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7650 10208 7656 10260
rect 7708 10208 7714 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9582 10248 9588 10260
rect 8444 10220 9588 10248
rect 8444 10208 8450 10220
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10778 10248 10784 10260
rect 10183 10220 10784 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 1486 10140 1492 10192
rect 1544 10180 1550 10192
rect 1581 10183 1639 10189
rect 1581 10180 1593 10183
rect 1544 10152 1593 10180
rect 1544 10140 1550 10152
rect 1581 10149 1593 10152
rect 1627 10149 1639 10183
rect 1581 10143 1639 10149
rect 2501 10183 2559 10189
rect 2501 10149 2513 10183
rect 2547 10180 2559 10183
rect 2774 10180 2780 10192
rect 2547 10152 2780 10180
rect 2547 10149 2559 10152
rect 2501 10143 2559 10149
rect 2774 10140 2780 10152
rect 2832 10140 2838 10192
rect 7668 10180 7696 10208
rect 7392 10152 7696 10180
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7282 10112 7288 10124
rect 6963 10084 7288 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7392 10121 7420 10152
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 10502 10180 10508 10192
rect 8352 10152 10508 10180
rect 8352 10140 8358 10152
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10081 7435 10115
rect 7644 10115 7702 10121
rect 7644 10112 7656 10115
rect 7377 10075 7435 10081
rect 7484 10084 7656 10112
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 1578 10044 1584 10056
rect 1535 10016 1584 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7484 10044 7512 10084
rect 7644 10081 7656 10084
rect 7690 10112 7702 10115
rect 9030 10112 9036 10124
rect 7690 10084 9036 10112
rect 7690 10081 7702 10084
rect 7644 10075 7702 10081
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 10091 10084 10180 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 7239 10016 7512 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 10152 9976 10180 10084
rect 10244 10053 10272 10152
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 10318 9976 10324 9988
rect 10152 9948 10324 9976
rect 10318 9936 10324 9948
rect 10376 9976 10382 9988
rect 10376 9948 10640 9976
rect 10376 9936 10382 9948
rect 6549 9911 6607 9917
rect 6549 9877 6561 9911
rect 6595 9908 6607 9911
rect 6914 9908 6920 9920
rect 6595 9880 6920 9908
rect 6595 9877 6607 9880
rect 6549 9871 6607 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 8110 9908 8116 9920
rect 7248 9880 8116 9908
rect 7248 9868 7254 9880
rect 8110 9868 8116 9880
rect 8168 9908 8174 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8168 9880 8769 9908
rect 8168 9868 8174 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 9674 9908 9680 9920
rect 9635 9880 9680 9908
rect 8757 9871 8815 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 10612 9917 10640 9948
rect 10597 9911 10655 9917
rect 10597 9877 10609 9911
rect 10643 9908 10655 9911
rect 10778 9908 10784 9920
rect 10643 9880 10784 9908
rect 10643 9877 10655 9880
rect 10597 9871 10655 9877
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 1104 9818 16008 9840
rect 1104 9766 3480 9818
rect 3532 9766 3544 9818
rect 3596 9766 3608 9818
rect 3660 9766 3672 9818
rect 3724 9766 8478 9818
rect 8530 9766 8542 9818
rect 8594 9766 8606 9818
rect 8658 9766 8670 9818
rect 8722 9766 13475 9818
rect 13527 9766 13539 9818
rect 13591 9766 13603 9818
rect 13655 9766 13667 9818
rect 13719 9766 16008 9818
rect 1104 9744 16008 9766
rect 7006 9664 7012 9716
rect 7064 9704 7070 9716
rect 7101 9707 7159 9713
rect 7101 9704 7113 9707
rect 7064 9676 7113 9704
rect 7064 9664 7070 9676
rect 7101 9673 7113 9676
rect 7147 9673 7159 9707
rect 7101 9667 7159 9673
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 8113 9707 8171 9713
rect 8113 9704 8125 9707
rect 7340 9676 8125 9704
rect 7340 9664 7346 9676
rect 8113 9673 8125 9676
rect 8159 9673 8171 9707
rect 8113 9667 8171 9673
rect 7466 9596 7472 9648
rect 7524 9636 7530 9648
rect 7929 9639 7987 9645
rect 7929 9636 7941 9639
rect 7524 9608 7941 9636
rect 7524 9596 7530 9608
rect 7929 9605 7941 9608
rect 7975 9605 7987 9639
rect 7929 9599 7987 9605
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 8294 9568 8300 9580
rect 7791 9540 8300 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 8294 9528 8300 9540
rect 8352 9568 8358 9580
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 8352 9540 8677 9568
rect 8352 9528 8358 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 9030 9528 9036 9580
rect 9088 9568 9094 9580
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 9088 9540 9505 9568
rect 9088 9528 9094 9540
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 7098 9460 7104 9512
rect 7156 9500 7162 9512
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 7156 9472 7481 9500
rect 7156 9460 7162 9472
rect 7469 9469 7481 9472
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9122 9500 9128 9512
rect 8619 9472 9128 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 9674 9500 9680 9512
rect 9447 9472 9680 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 8110 9432 8116 9444
rect 5500 9404 8116 9432
rect 5500 9392 5506 9404
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 8846 9432 8852 9444
rect 8527 9404 8852 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 8846 9392 8852 9404
rect 8904 9432 8910 9444
rect 9309 9435 9367 9441
rect 8904 9404 9260 9432
rect 8904 9392 8910 9404
rect 1489 9367 1547 9373
rect 1489 9333 1501 9367
rect 1535 9364 1547 9367
rect 1578 9364 1584 9376
rect 1535 9336 1584 9364
rect 1535 9333 1547 9336
rect 1489 9327 1547 9333
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 8938 9364 8944 9376
rect 8899 9336 8944 9364
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9232 9364 9260 9404
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9950 9432 9956 9444
rect 9355 9404 9956 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9950 9392 9956 9404
rect 10008 9392 10014 9444
rect 9769 9367 9827 9373
rect 9769 9364 9781 9367
rect 9232 9336 9781 9364
rect 9769 9333 9781 9336
rect 9815 9364 9827 9367
rect 12894 9364 12900 9376
rect 9815 9336 12900 9364
rect 9815 9333 9827 9336
rect 9769 9327 9827 9333
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 1104 9274 16008 9296
rect 1104 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 10976 9274
rect 11028 9222 11040 9274
rect 11092 9222 11104 9274
rect 11156 9222 11168 9274
rect 11220 9222 16008 9274
rect 1104 9200 16008 9222
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6972 9132 7021 9160
rect 6972 9120 6978 9132
rect 7009 9129 7021 9132
rect 7055 9129 7067 9163
rect 7009 9123 7067 9129
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 8938 9024 8944 9036
rect 6963 8996 8944 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 13354 9024 13360 9036
rect 12667 8996 13360 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 7190 8956 7196 8968
rect 7151 8928 7196 8956
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 11388 8928 12817 8956
rect 11388 8916 11394 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 4212 8792 6561 8820
rect 4212 8780 4218 8792
rect 6549 8789 6561 8792
rect 6595 8789 6607 8823
rect 6549 8783 6607 8789
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13412 8792 13553 8820
rect 13412 8780 13418 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 1104 8730 16008 8752
rect 1104 8678 3480 8730
rect 3532 8678 3544 8730
rect 3596 8678 3608 8730
rect 3660 8678 3672 8730
rect 3724 8678 8478 8730
rect 8530 8678 8542 8730
rect 8594 8678 8606 8730
rect 8658 8678 8670 8730
rect 8722 8678 13475 8730
rect 13527 8678 13539 8730
rect 13591 8678 13603 8730
rect 13655 8678 13667 8730
rect 13719 8678 16008 8730
rect 1104 8656 16008 8678
rect 1104 8186 16008 8208
rect 1104 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 10976 8186
rect 11028 8134 11040 8186
rect 11092 8134 11104 8186
rect 11156 8134 11168 8186
rect 11220 8134 16008 8186
rect 1104 8112 16008 8134
rect 1104 7642 16008 7664
rect 1104 7590 3480 7642
rect 3532 7590 3544 7642
rect 3596 7590 3608 7642
rect 3660 7590 3672 7642
rect 3724 7590 8478 7642
rect 8530 7590 8542 7642
rect 8594 7590 8606 7642
rect 8658 7590 8670 7642
rect 8722 7590 13475 7642
rect 13527 7590 13539 7642
rect 13591 7590 13603 7642
rect 13655 7590 13667 7642
rect 13719 7590 16008 7642
rect 1104 7568 16008 7590
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4154 7324 4160 7336
rect 3375 7296 4160 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 2958 7216 2964 7268
rect 3016 7256 3022 7268
rect 3605 7259 3663 7265
rect 3605 7256 3617 7259
rect 3016 7228 3617 7256
rect 3016 7216 3022 7228
rect 3605 7225 3617 7228
rect 3651 7225 3663 7259
rect 3605 7219 3663 7225
rect 1104 7098 16008 7120
rect 1104 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 10976 7098
rect 11028 7046 11040 7098
rect 11092 7046 11104 7098
rect 11156 7046 11168 7098
rect 11220 7046 16008 7098
rect 1104 7024 16008 7046
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 7282 6712 7288 6724
rect 4028 6684 7288 6712
rect 4028 6672 4034 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 9674 6644 9680 6656
rect 5684 6616 9680 6644
rect 5684 6604 5690 6616
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 1104 6554 16008 6576
rect 1104 6502 3480 6554
rect 3532 6502 3544 6554
rect 3596 6502 3608 6554
rect 3660 6502 3672 6554
rect 3724 6502 8478 6554
rect 8530 6502 8542 6554
rect 8594 6502 8606 6554
rect 8658 6502 8670 6554
rect 8722 6502 13475 6554
rect 13527 6502 13539 6554
rect 13591 6502 13603 6554
rect 13655 6502 13667 6554
rect 13719 6502 16008 6554
rect 1104 6480 16008 6502
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6972 6412 7021 6440
rect 6972 6400 6978 6412
rect 7009 6409 7021 6412
rect 7055 6440 7067 6443
rect 7834 6440 7840 6452
rect 7055 6412 7840 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 11422 6440 11428 6452
rect 7984 6412 11428 6440
rect 7984 6400 7990 6412
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 9306 6372 9312 6384
rect 4856 6344 9312 6372
rect 4856 6332 4862 6344
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7616 6276 7849 6304
rect 7616 6264 7622 6276
rect 7837 6273 7849 6276
rect 7883 6304 7895 6307
rect 11882 6304 11888 6316
rect 7883 6276 11888 6304
rect 7883 6273 7895 6276
rect 7837 6267 7895 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7156 6208 7389 6236
rect 7156 6196 7162 6208
rect 7377 6205 7389 6208
rect 7423 6236 7435 6239
rect 7926 6236 7932 6248
rect 7423 6208 7932 6236
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 7926 6196 7932 6208
rect 7984 6196 7990 6248
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 11698 6236 11704 6248
rect 8904 6208 11704 6236
rect 8904 6196 8910 6208
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 7466 6168 7472 6180
rect 5132 6140 7472 6168
rect 5132 6128 5138 6140
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 7834 6128 7840 6180
rect 7892 6168 7898 6180
rect 12250 6168 12256 6180
rect 7892 6140 12256 6168
rect 7892 6128 7898 6140
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 8662 6100 8668 6112
rect 7800 6072 8668 6100
rect 7800 6060 7806 6072
rect 8662 6060 8668 6072
rect 8720 6100 8726 6112
rect 10686 6100 10692 6112
rect 8720 6072 10692 6100
rect 8720 6060 8726 6072
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 13998 6100 14004 6112
rect 10928 6072 14004 6100
rect 10928 6060 10934 6072
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 1104 6010 16008 6032
rect 1104 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 10976 6010
rect 11028 5958 11040 6010
rect 11092 5958 11104 6010
rect 11156 5958 11168 6010
rect 11220 5958 16008 6010
rect 1104 5936 16008 5958
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 4488 5868 7941 5896
rect 4488 5856 4494 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 9180 5868 9873 5896
rect 9180 5856 9186 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 10870 5896 10876 5908
rect 10831 5868 10876 5896
rect 9861 5859 9919 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11514 5896 11520 5908
rect 11287 5868 11520 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 5074 5828 5080 5840
rect 4448 5800 5080 5828
rect 4448 5769 4476 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5626 5828 5632 5840
rect 5184 5800 5632 5828
rect 5184 5769 5212 5800
rect 5626 5788 5632 5800
rect 5684 5788 5690 5840
rect 8846 5828 8852 5840
rect 8220 5800 8852 5828
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5729 4123 5763
rect 4065 5723 4123 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5729 4491 5763
rect 4433 5723 4491 5729
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6595 5732 6837 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7098 5760 7104 5772
rect 7055 5732 7104 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 4080 5692 4108 5723
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 7558 5760 7564 5772
rect 7423 5732 7564 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7742 5760 7748 5772
rect 7703 5732 7748 5760
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 8220 5769 8248 5800
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 10888 5828 10916 5856
rect 9692 5800 10916 5828
rect 8211 5763 8269 5769
rect 8211 5729 8223 5763
rect 8257 5729 8269 5763
rect 8662 5760 8668 5772
rect 8623 5732 8668 5760
rect 8211 5723 8269 5729
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 9030 5760 9036 5772
rect 8991 5732 9036 5760
rect 9030 5720 9036 5732
rect 9088 5760 9094 5772
rect 9692 5769 9720 5800
rect 9401 5763 9459 5769
rect 9401 5760 9413 5763
rect 9088 5732 9413 5760
rect 9088 5720 9094 5732
rect 9401 5729 9413 5732
rect 9447 5729 9459 5763
rect 9401 5723 9459 5729
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 11256 5760 11284 5859
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 12250 5896 12256 5908
rect 12211 5868 12256 5896
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12713 5899 12771 5905
rect 12713 5865 12725 5899
rect 12759 5896 12771 5899
rect 15378 5896 15384 5908
rect 12759 5868 15384 5896
rect 12759 5865 12771 5868
rect 12713 5859 12771 5865
rect 10459 5732 11284 5760
rect 11609 5763 11667 5769
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 11609 5729 11621 5763
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 12069 5763 12127 5769
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12728 5760 12756 5859
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 12115 5732 12756 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 4798 5692 4804 5704
rect 4080 5664 4804 5692
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 4890 5652 4896 5704
rect 4948 5692 4954 5704
rect 10060 5692 10088 5723
rect 11624 5692 11652 5723
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 4948 5664 9260 5692
rect 10060 5664 11100 5692
rect 11624 5664 12541 5692
rect 4948 5652 4954 5664
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 6733 5627 6791 5633
rect 6733 5624 6745 5627
rect 4764 5596 6745 5624
rect 4764 5584 4770 5596
rect 6733 5593 6745 5596
rect 6779 5593 6791 5627
rect 6914 5624 6920 5636
rect 6875 5596 6920 5624
rect 6733 5587 6791 5593
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 9232 5633 9260 5664
rect 11072 5633 11100 5664
rect 12529 5661 12541 5664
rect 12575 5692 12587 5695
rect 15286 5692 15292 5704
rect 12575 5664 15292 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 9217 5627 9275 5633
rect 7524 5596 8892 5624
rect 7524 5584 7530 5596
rect 4246 5556 4252 5568
rect 4207 5528 4252 5556
rect 4246 5516 4252 5528
rect 4304 5516 4310 5568
rect 4614 5556 4620 5568
rect 4575 5528 4620 5556
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7190 5556 7196 5568
rect 7151 5528 7196 5556
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 7558 5556 7564 5568
rect 7519 5528 7564 5556
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 8389 5559 8447 5565
rect 8389 5556 8401 5559
rect 7708 5528 8401 5556
rect 7708 5516 7714 5528
rect 8389 5525 8401 5528
rect 8435 5525 8447 5559
rect 8864 5556 8892 5596
rect 9217 5593 9229 5627
rect 9263 5593 9275 5627
rect 11057 5627 11115 5633
rect 9217 5587 9275 5593
rect 9324 5596 10732 5624
rect 9324 5556 9352 5596
rect 8864 5528 9352 5556
rect 8389 5519 8447 5525
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10229 5559 10287 5565
rect 10229 5556 10241 5559
rect 10008 5528 10241 5556
rect 10008 5516 10014 5528
rect 10229 5525 10241 5528
rect 10275 5525 10287 5559
rect 10229 5519 10287 5525
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 10376 5528 10609 5556
rect 10376 5516 10382 5528
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10704 5556 10732 5596
rect 11057 5593 11069 5627
rect 11103 5624 11115 5627
rect 11974 5624 11980 5636
rect 11103 5596 11980 5624
rect 11103 5593 11115 5596
rect 11057 5587 11115 5593
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 10704 5528 11805 5556
rect 10597 5519 10655 5525
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 1104 5466 16008 5488
rect 1104 5414 3480 5466
rect 3532 5414 3544 5466
rect 3596 5414 3608 5466
rect 3660 5414 3672 5466
rect 3724 5414 8478 5466
rect 8530 5414 8542 5466
rect 8594 5414 8606 5466
rect 8658 5414 8670 5466
rect 8722 5414 13475 5466
rect 13527 5414 13539 5466
rect 13591 5414 13603 5466
rect 13655 5414 13667 5466
rect 13719 5414 16008 5466
rect 1104 5392 16008 5414
rect 934 5312 940 5364
rect 992 5352 998 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 992 5324 5365 5352
rect 992 5312 998 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5997 5355 6055 5361
rect 5997 5352 6009 5355
rect 5353 5315 5411 5321
rect 5460 5324 6009 5352
rect 2682 5244 2688 5296
rect 2740 5284 2746 5296
rect 5460 5284 5488 5324
rect 5997 5321 6009 5324
rect 6043 5321 6055 5355
rect 5997 5315 6055 5321
rect 7282 5312 7288 5364
rect 7340 5352 7346 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7340 5324 7389 5352
rect 7340 5312 7346 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 7377 5315 7435 5321
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 8168 5324 9321 5352
rect 8168 5312 8174 5324
rect 9309 5321 9321 5324
rect 9355 5321 9367 5355
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 9309 5315 9367 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 10100 5324 10241 5352
rect 10100 5312 10106 5324
rect 10229 5321 10241 5324
rect 10275 5321 10287 5355
rect 10594 5352 10600 5364
rect 10555 5324 10600 5352
rect 10229 5315 10287 5321
rect 10594 5312 10600 5324
rect 10652 5312 10658 5364
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12894 5312 12900 5364
rect 12952 5352 12958 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12952 5324 13001 5352
rect 12952 5312 12958 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 14001 5355 14059 5361
rect 14001 5352 14013 5355
rect 13228 5324 14013 5352
rect 13228 5312 13234 5324
rect 14001 5321 14013 5324
rect 14047 5352 14059 5355
rect 15562 5352 15568 5364
rect 14047 5324 15568 5352
rect 14047 5321 14059 5324
rect 14001 5315 14059 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 8294 5284 8300 5296
rect 2740 5256 5488 5284
rect 7484 5256 8300 5284
rect 2740 5244 2746 5256
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 5828 5188 6653 5216
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 5074 5148 5080 5160
rect 4847 5120 5080 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5169 5151 5227 5157
rect 5169 5117 5181 5151
rect 5215 5148 5227 5151
rect 5626 5148 5632 5160
rect 5215 5120 5632 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 5626 5108 5632 5120
rect 5684 5108 5690 5160
rect 5828 5157 5856 5188
rect 6641 5185 6653 5188
rect 6687 5216 6699 5219
rect 6914 5216 6920 5228
rect 6687 5188 6920 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7282 5216 7288 5228
rect 7116 5188 7288 5216
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5117 5871 5151
rect 5813 5111 5871 5117
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6546 5148 6552 5160
rect 6227 5120 6552 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7116 5148 7144 5188
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 6871 5120 7144 5148
rect 7193 5151 7251 5157
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7484 5148 7512 5256
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 9858 5244 9864 5296
rect 9916 5284 9922 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 9916 5256 11897 5284
rect 9916 5244 9922 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 15194 5284 15200 5296
rect 11885 5247 11943 5253
rect 12084 5256 15200 5284
rect 9674 5216 9680 5228
rect 8312 5188 9680 5216
rect 7239 5120 7512 5148
rect 7561 5151 7619 5157
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7561 5117 7573 5151
rect 7607 5148 7619 5151
rect 7742 5148 7748 5160
rect 7607 5120 7748 5148
rect 7607 5117 7619 5120
rect 7561 5111 7619 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 7926 5148 7932 5160
rect 7887 5120 7932 5148
rect 7926 5108 7932 5120
rect 7984 5108 7990 5160
rect 8312 5157 8340 5188
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 12084 5225 12112 5256
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 12069 5219 12127 5225
rect 12069 5216 12081 5219
rect 10888 5188 12081 5216
rect 8297 5151 8355 5157
rect 8297 5117 8309 5151
rect 8343 5117 8355 5151
rect 8662 5148 8668 5160
rect 8623 5120 8668 5148
rect 8297 5111 8355 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5117 9183 5151
rect 9582 5148 9588 5160
rect 9543 5120 9588 5148
rect 9125 5111 9183 5117
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 9140 5080 9168 5111
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 10042 5148 10048 5160
rect 10003 5120 10048 5148
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10888 5157 10916 5188
rect 12069 5185 12081 5188
rect 12115 5185 12127 5219
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 12069 5179 12127 5185
rect 12452 5188 13645 5216
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 11606 5148 11612 5160
rect 11287 5120 11612 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 9766 5080 9772 5092
rect 4212 5052 8892 5080
rect 9140 5052 9772 5080
rect 4212 5040 4218 5052
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5626 5012 5632 5024
rect 5587 4984 5632 5012
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 7156 4984 7757 5012
rect 7156 4972 7162 4984
rect 7745 4981 7757 4984
rect 7791 4981 7803 5015
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 7745 4975 7803 4981
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 8478 5012 8484 5024
rect 8439 4984 8484 5012
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 8864 5021 8892 5052
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 10428 5080 10456 5111
rect 11606 5108 11612 5120
rect 11664 5108 11670 5160
rect 11701 5151 11759 5157
rect 11701 5117 11713 5151
rect 11747 5148 11759 5151
rect 12342 5148 12348 5160
rect 11747 5120 12348 5148
rect 11747 5117 11759 5120
rect 11701 5111 11759 5117
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12452 5157 12480 5188
rect 13633 5185 13645 5188
rect 13679 5216 13691 5219
rect 16482 5216 16488 5228
rect 13679 5188 16488 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5117 12863 5151
rect 13170 5148 13176 5160
rect 13131 5120 13176 5148
rect 12805 5111 12863 5117
rect 11330 5080 11336 5092
rect 10428 5052 11336 5080
rect 11330 5040 11336 5052
rect 11388 5040 11394 5092
rect 12820 5080 12848 5111
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 12820 5052 13860 5080
rect 13832 5024 13860 5052
rect 8849 5015 8907 5021
rect 8849 4981 8861 5015
rect 8895 4981 8907 5015
rect 11422 5012 11428 5024
rect 11383 4984 11428 5012
rect 8849 4975 8907 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 13354 5012 13360 5024
rect 13315 4984 13360 5012
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13814 5012 13820 5024
rect 13775 4984 13820 5012
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 1104 4922 16008 4944
rect 1104 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 10976 4922
rect 11028 4870 11040 4922
rect 11092 4870 11104 4922
rect 11156 4870 11168 4922
rect 11220 4870 16008 4922
rect 1104 4848 16008 4870
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 8478 4808 8484 4820
rect 5316 4780 8484 4808
rect 5316 4768 5322 4780
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 8720 4780 9137 4808
rect 8720 4768 8726 4780
rect 9125 4777 9137 4780
rect 9171 4808 9183 4811
rect 10134 4808 10140 4820
rect 9171 4780 10140 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11606 4808 11612 4820
rect 11567 4780 11612 4808
rect 11606 4768 11612 4780
rect 11664 4808 11670 4820
rect 13078 4808 13084 4820
rect 11664 4780 13084 4808
rect 11664 4768 11670 4780
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 3878 4700 3884 4752
rect 3936 4740 3942 4752
rect 7098 4740 7104 4752
rect 3936 4712 7104 4740
rect 3936 4700 3942 4712
rect 7098 4700 7104 4712
rect 7156 4700 7162 4752
rect 8110 4740 8116 4752
rect 7668 4712 8116 4740
rect 3786 4632 3792 4684
rect 3844 4672 3850 4684
rect 7668 4672 7696 4712
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 15654 4740 15660 4752
rect 10836 4712 15660 4740
rect 10836 4700 10842 4712
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 3844 4644 7696 4672
rect 3844 4632 3850 4644
rect 7742 4632 7748 4684
rect 7800 4672 7806 4684
rect 8021 4675 8079 4681
rect 8021 4672 8033 4675
rect 7800 4644 8033 4672
rect 7800 4632 7806 4644
rect 8021 4641 8033 4644
rect 8067 4672 8079 4675
rect 8846 4672 8852 4684
rect 8067 4644 8852 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8846 4632 8852 4644
rect 8904 4632 8910 4684
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 10137 4675 10195 4681
rect 10137 4672 10149 4675
rect 9263 4644 10149 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 10137 4641 10149 4644
rect 10183 4672 10195 4675
rect 10410 4672 10416 4684
rect 10183 4644 10416 4672
rect 10183 4641 10195 4644
rect 10137 4635 10195 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8294 4604 8300 4616
rect 7699 4576 8300 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9640 4576 9965 4604
rect 9640 4564 9646 4576
rect 9953 4573 9965 4576
rect 9999 4604 10011 4607
rect 13906 4604 13912 4616
rect 9999 4576 13912 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 2498 4496 2504 4548
rect 2556 4536 2562 4548
rect 7006 4536 7012 4548
rect 2556 4508 7012 4536
rect 2556 4496 2562 4508
rect 7006 4496 7012 4508
rect 7064 4496 7070 4548
rect 8757 4539 8815 4545
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 9674 4536 9680 4548
rect 8803 4508 9680 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 10505 4539 10563 4545
rect 10505 4536 10517 4539
rect 10100 4508 10517 4536
rect 10100 4496 10106 4508
rect 10505 4505 10517 4508
rect 10551 4536 10563 4539
rect 11054 4536 11060 4548
rect 10551 4508 11060 4536
rect 10551 4505 10563 4508
rect 10505 4499 10563 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 5258 4468 5264 4480
rect 5219 4440 5264 4468
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 7282 4468 7288 4480
rect 7243 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 7926 4428 7932 4480
rect 7984 4468 7990 4480
rect 8389 4471 8447 4477
rect 8389 4468 8401 4471
rect 7984 4440 8401 4468
rect 7984 4428 7990 4440
rect 8389 4437 8401 4440
rect 8435 4468 8447 4471
rect 8938 4468 8944 4480
rect 8435 4440 8944 4468
rect 8435 4437 8447 4440
rect 8389 4431 8447 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9398 4468 9404 4480
rect 9359 4440 9404 4468
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 9766 4468 9772 4480
rect 9727 4440 9772 4468
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 11146 4468 11152 4480
rect 10919 4440 11152 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 12161 4471 12219 4477
rect 12161 4437 12173 4471
rect 12207 4468 12219 4471
rect 12434 4468 12440 4480
rect 12207 4440 12440 4468
rect 12207 4437 12219 4440
rect 12161 4431 12219 4437
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 1104 4378 16008 4400
rect 1104 4326 3480 4378
rect 3532 4326 3544 4378
rect 3596 4326 3608 4378
rect 3660 4326 3672 4378
rect 3724 4326 8478 4378
rect 8530 4326 8542 4378
rect 8594 4326 8606 4378
rect 8658 4326 8670 4378
rect 8722 4326 13475 4378
rect 13527 4326 13539 4378
rect 13591 4326 13603 4378
rect 13655 4326 13667 4378
rect 13719 4326 16008 4378
rect 1104 4304 16008 4326
rect 5258 4224 5264 4276
rect 5316 4264 5322 4276
rect 9214 4264 9220 4276
rect 5316 4236 9220 4264
rect 5316 4224 5322 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 6638 4156 6644 4208
rect 6696 4196 6702 4208
rect 10502 4196 10508 4208
rect 6696 4168 10508 4196
rect 6696 4156 6702 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 7190 4128 7196 4140
rect 2832 4100 7196 4128
rect 2832 4088 2838 4100
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 13262 4128 13268 4140
rect 9824 4100 13268 4128
rect 9824 4088 9830 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 16942 4128 16948 4140
rect 13872 4100 16948 4128
rect 13872 4088 13878 4100
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 7558 4060 7564 4072
rect 3200 4032 7564 4060
rect 3200 4020 3206 4032
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 11054 4020 11060 4072
rect 11112 4060 11118 4072
rect 14366 4060 14372 4072
rect 11112 4032 14372 4060
rect 11112 4020 11118 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 9214 3992 9220 4004
rect 5684 3964 9220 3992
rect 5684 3952 5690 3964
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 14734 3992 14740 4004
rect 11204 3964 14740 3992
rect 11204 3952 11210 3964
rect 14734 3952 14740 3964
rect 14792 3952 14798 4004
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 11422 3924 11428 3936
rect 6696 3896 11428 3924
rect 6696 3884 6702 3896
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 1104 3834 16008 3856
rect 1104 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 10976 3834
rect 11028 3782 11040 3834
rect 11092 3782 11104 3834
rect 11156 3782 11168 3834
rect 11220 3782 16008 3834
rect 1104 3760 16008 3782
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 10042 3720 10048 3732
rect 6972 3692 10048 3720
rect 6972 3680 6978 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 9398 3652 9404 3664
rect 7064 3624 9404 3652
rect 7064 3612 7070 3624
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 10870 3584 10876 3596
rect 7340 3556 10876 3584
rect 7340 3544 7346 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 7650 3516 7656 3528
rect 4120 3488 7656 3516
rect 4120 3476 4126 3488
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 11330 3516 11336 3528
rect 8352 3488 11336 3516
rect 8352 3476 8358 3488
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 8846 3408 8852 3460
rect 8904 3448 8910 3460
rect 11790 3448 11796 3460
rect 8904 3420 11796 3448
rect 8904 3408 8910 3420
rect 11790 3408 11796 3420
rect 11848 3408 11854 3460
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 12158 3380 12164 3392
rect 8996 3352 12164 3380
rect 8996 3340 9002 3352
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 1104 3290 16008 3312
rect 1104 3238 3480 3290
rect 3532 3238 3544 3290
rect 3596 3238 3608 3290
rect 3660 3238 3672 3290
rect 3724 3238 8478 3290
rect 8530 3238 8542 3290
rect 8594 3238 8606 3290
rect 8658 3238 8670 3290
rect 8722 3238 13475 3290
rect 13527 3238 13539 3290
rect 13591 3238 13603 3290
rect 13655 3238 13667 3290
rect 13719 3238 16008 3290
rect 1104 3216 16008 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 4706 3176 4712 3188
rect 2372 3148 4712 3176
rect 2372 3136 2378 3148
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 9950 3176 9956 3188
rect 5776 3148 9956 3176
rect 5776 3136 5782 3148
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 16022 3176 16028 3188
rect 12492 3148 16028 3176
rect 12492 3136 12498 3148
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 5350 3108 5356 3120
rect 1912 3080 5356 3108
rect 1912 3068 1918 3080
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 8846 3108 8852 3120
rect 7432 3080 8852 3108
rect 7432 3068 7438 3080
rect 8846 3068 8852 3080
rect 8904 3068 8910 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 12618 3108 12624 3120
rect 9732 3080 12624 3108
rect 9732 3068 9738 3080
rect 12618 3068 12624 3080
rect 12676 3068 12682 3120
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 6362 3040 6368 3052
rect 1544 3012 6368 3040
rect 1544 3000 1550 3012
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 566 2932 572 2984
rect 624 2972 630 2984
rect 4982 2972 4988 2984
rect 624 2944 4988 2972
rect 624 2932 630 2944
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 10318 2972 10324 2984
rect 6328 2944 10324 2972
rect 6328 2932 6334 2944
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 4246 2904 4252 2916
rect 256 2876 4252 2904
rect 256 2864 262 2876
rect 4246 2864 4252 2876
rect 4304 2864 4310 2916
rect 1026 2796 1032 2848
rect 1084 2836 1090 2848
rect 4614 2836 4620 2848
rect 1084 2808 4620 2836
rect 1084 2796 1090 2808
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 13354 2836 13360 2848
rect 8352 2808 13360 2836
rect 8352 2796 8358 2808
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 1104 2746 16008 2768
rect 1104 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 10976 2746
rect 11028 2694 11040 2746
rect 11092 2694 11104 2746
rect 11156 2694 11168 2746
rect 11220 2694 16008 2746
rect 1104 2672 16008 2694
rect 1104 2202 16008 2224
rect 1104 2150 3480 2202
rect 3532 2150 3544 2202
rect 3596 2150 3608 2202
rect 3660 2150 3672 2202
rect 3724 2150 8478 2202
rect 8530 2150 8542 2202
rect 8594 2150 8606 2202
rect 8658 2150 8670 2202
rect 8722 2150 13475 2202
rect 13527 2150 13539 2202
rect 13591 2150 13603 2202
rect 13655 2150 13667 2202
rect 13719 2150 16008 2202
rect 1104 2128 16008 2150
<< via1 >>
rect 5264 17892 5316 17944
rect 5448 17892 5500 17944
rect 3480 17382 3532 17434
rect 3544 17382 3596 17434
rect 3608 17382 3660 17434
rect 3672 17382 3724 17434
rect 8478 17382 8530 17434
rect 8542 17382 8594 17434
rect 8606 17382 8658 17434
rect 8670 17382 8722 17434
rect 13475 17382 13527 17434
rect 13539 17382 13591 17434
rect 13603 17382 13655 17434
rect 13667 17382 13719 17434
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 10976 16838 11028 16890
rect 11040 16838 11092 16890
rect 11104 16838 11156 16890
rect 11168 16838 11220 16890
rect 7840 16532 7892 16584
rect 10876 16532 10928 16584
rect 3480 16294 3532 16346
rect 3544 16294 3596 16346
rect 3608 16294 3660 16346
rect 3672 16294 3724 16346
rect 8478 16294 8530 16346
rect 8542 16294 8594 16346
rect 8606 16294 8658 16346
rect 8670 16294 8722 16346
rect 13475 16294 13527 16346
rect 13539 16294 13591 16346
rect 13603 16294 13655 16346
rect 13667 16294 13719 16346
rect 6460 16056 6512 16108
rect 10600 16056 10652 16108
rect 7104 15988 7156 16040
rect 9772 15988 9824 16040
rect 5632 15920 5684 15972
rect 9680 15920 9732 15972
rect 13084 15920 13136 15972
rect 15292 15920 15344 15972
rect 3792 15852 3844 15904
rect 3976 15852 4028 15904
rect 4344 15852 4396 15904
rect 5356 15852 5408 15904
rect 7748 15852 7800 15904
rect 9772 15852 9824 15904
rect 10140 15852 10192 15904
rect 12348 15852 12400 15904
rect 13820 15852 13872 15904
rect 15660 15852 15712 15904
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 10976 15750 11028 15802
rect 11040 15750 11092 15802
rect 11104 15750 11156 15802
rect 11168 15750 11220 15802
rect 1860 15648 1912 15700
rect 2688 15648 2740 15700
rect 3056 15648 3108 15700
rect 3976 15648 4028 15700
rect 9036 15648 9088 15700
rect 13360 15648 13412 15700
rect 6276 15580 6328 15632
rect 9956 15580 10008 15632
rect 10784 15580 10836 15632
rect 13176 15580 13228 15632
rect 2228 15512 2280 15564
rect 5540 15512 5592 15564
rect 8852 15512 8904 15564
rect 9404 15512 9456 15564
rect 1400 15444 1452 15496
rect 4712 15444 4764 15496
rect 204 15376 256 15428
rect 2872 15376 2924 15428
rect 11980 15376 12032 15428
rect 14464 15376 14516 15428
rect 4804 15308 4856 15360
rect 6736 15308 6788 15360
rect 7288 15308 7340 15360
rect 9588 15308 9640 15360
rect 11704 15308 11756 15360
rect 12716 15308 12768 15360
rect 3480 15206 3532 15258
rect 3544 15206 3596 15258
rect 3608 15206 3660 15258
rect 3672 15206 3724 15258
rect 8478 15206 8530 15258
rect 8542 15206 8594 15258
rect 8606 15206 8658 15258
rect 8670 15206 8722 15258
rect 13475 15206 13527 15258
rect 13539 15206 13591 15258
rect 13603 15206 13655 15258
rect 13667 15206 13719 15258
rect 572 15104 624 15156
rect 4712 15147 4764 15156
rect 4712 15113 4721 15147
rect 4721 15113 4755 15147
rect 4755 15113 4764 15147
rect 4712 15104 4764 15113
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 7196 15036 7248 15088
rect 5540 14968 5592 15020
rect 9864 14764 9916 14816
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 10976 14662 11028 14714
rect 11040 14662 11092 14714
rect 11104 14662 11156 14714
rect 11168 14662 11220 14714
rect 6736 14560 6788 14612
rect 9588 14560 9640 14612
rect 10048 14424 10100 14476
rect 11520 14424 11572 14476
rect 14832 14424 14884 14476
rect 8852 14220 8904 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 3480 14118 3532 14170
rect 3544 14118 3596 14170
rect 3608 14118 3660 14170
rect 3672 14118 3724 14170
rect 8478 14118 8530 14170
rect 8542 14118 8594 14170
rect 8606 14118 8658 14170
rect 8670 14118 8722 14170
rect 13475 14118 13527 14170
rect 13539 14118 13591 14170
rect 13603 14118 13655 14170
rect 13667 14118 13719 14170
rect 4068 14016 4120 14068
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 10976 13574 11028 13626
rect 11040 13574 11092 13626
rect 11104 13574 11156 13626
rect 11168 13574 11220 13626
rect 2872 13472 2924 13524
rect 4344 13472 4396 13524
rect 15476 13515 15528 13524
rect 15476 13481 15485 13515
rect 15485 13481 15519 13515
rect 15519 13481 15528 13515
rect 15476 13472 15528 13481
rect 6276 13336 6328 13388
rect 9312 13268 9364 13320
rect 3240 13132 3292 13184
rect 14464 13132 14516 13184
rect 3480 13030 3532 13082
rect 3544 13030 3596 13082
rect 3608 13030 3660 13082
rect 3672 13030 3724 13082
rect 8478 13030 8530 13082
rect 8542 13030 8594 13082
rect 8606 13030 8658 13082
rect 8670 13030 8722 13082
rect 13475 13030 13527 13082
rect 13539 13030 13591 13082
rect 13603 13030 13655 13082
rect 13667 13030 13719 13082
rect 9312 12588 9364 12640
rect 13728 12588 13780 12640
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 10976 12486 11028 12538
rect 11040 12486 11092 12538
rect 11104 12486 11156 12538
rect 11168 12486 11220 12538
rect 6276 12384 6328 12436
rect 6736 12384 6788 12436
rect 11428 12384 11480 12436
rect 11612 12384 11664 12436
rect 11336 12248 11388 12300
rect 3480 11942 3532 11994
rect 3544 11942 3596 11994
rect 3608 11942 3660 11994
rect 3672 11942 3724 11994
rect 8478 11942 8530 11994
rect 8542 11942 8594 11994
rect 8606 11942 8658 11994
rect 8670 11942 8722 11994
rect 13475 11942 13527 11994
rect 13539 11942 13591 11994
rect 13603 11942 13655 11994
rect 13667 11942 13719 11994
rect 15568 11704 15620 11756
rect 16948 11704 17000 11756
rect 7472 11636 7524 11688
rect 15384 11636 15436 11688
rect 16488 11636 16540 11688
rect 5724 11568 5776 11620
rect 7288 11568 7340 11620
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 7472 11500 7524 11552
rect 8300 11500 8352 11552
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 10976 11398 11028 11450
rect 11040 11398 11092 11450
rect 11104 11398 11156 11450
rect 11168 11398 11220 11450
rect 6736 11228 6788 11280
rect 9312 11296 9364 11348
rect 7380 11160 7432 11212
rect 8944 11228 8996 11280
rect 9864 11228 9916 11280
rect 8116 11203 8168 11212
rect 8116 11169 8150 11203
rect 8150 11169 8168 11203
rect 8116 11160 8168 11169
rect 9312 11203 9364 11212
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 7012 11024 7064 11076
rect 7564 11067 7616 11076
rect 7564 11033 7573 11067
rect 7573 11033 7607 11067
rect 7607 11033 7616 11067
rect 7564 11024 7616 11033
rect 7288 10956 7340 11008
rect 9496 10956 9548 11008
rect 10692 11228 10744 11280
rect 3480 10854 3532 10906
rect 3544 10854 3596 10906
rect 3608 10854 3660 10906
rect 3672 10854 3724 10906
rect 8478 10854 8530 10906
rect 8542 10854 8594 10906
rect 8606 10854 8658 10906
rect 8670 10854 8722 10906
rect 13475 10854 13527 10906
rect 13539 10854 13591 10906
rect 13603 10854 13655 10906
rect 13667 10854 13719 10906
rect 3332 10752 3384 10804
rect 5540 10684 5592 10736
rect 7196 10684 7248 10736
rect 7288 10616 7340 10668
rect 7564 10616 7616 10668
rect 10876 10752 10928 10804
rect 13820 10752 13872 10804
rect 10048 10616 10100 10668
rect 10324 10616 10376 10668
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 1492 10548 1544 10600
rect 3240 10548 3292 10600
rect 7104 10548 7156 10600
rect 7472 10548 7524 10600
rect 8300 10480 8352 10532
rect 9864 10480 9916 10532
rect 10232 10480 10284 10532
rect 14464 10480 14516 10532
rect 7104 10412 7156 10464
rect 7196 10412 7248 10464
rect 8392 10412 8444 10464
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9496 10455 9548 10464
rect 9128 10412 9180 10421
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 10416 10455 10468 10464
rect 10416 10421 10425 10455
rect 10425 10421 10459 10455
rect 10459 10421 10468 10455
rect 10416 10412 10468 10421
rect 10876 10412 10928 10464
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 10976 10310 11028 10362
rect 11040 10310 11092 10362
rect 11104 10310 11156 10362
rect 11168 10310 11220 10362
rect 7012 10208 7064 10260
rect 7564 10208 7616 10260
rect 7656 10208 7708 10260
rect 8392 10208 8444 10260
rect 9588 10208 9640 10260
rect 10784 10251 10836 10260
rect 10784 10217 10793 10251
rect 10793 10217 10827 10251
rect 10827 10217 10836 10251
rect 10784 10208 10836 10217
rect 1492 10140 1544 10192
rect 2780 10140 2832 10192
rect 7288 10072 7340 10124
rect 8300 10140 8352 10192
rect 1584 10004 1636 10056
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 9036 10072 9088 10124
rect 10508 10140 10560 10192
rect 10324 9936 10376 9988
rect 6920 9868 6972 9920
rect 7196 9868 7248 9920
rect 8116 9868 8168 9920
rect 9680 9911 9732 9920
rect 9680 9877 9689 9911
rect 9689 9877 9723 9911
rect 9723 9877 9732 9911
rect 9680 9868 9732 9877
rect 10784 9868 10836 9920
rect 3480 9766 3532 9818
rect 3544 9766 3596 9818
rect 3608 9766 3660 9818
rect 3672 9766 3724 9818
rect 8478 9766 8530 9818
rect 8542 9766 8594 9818
rect 8606 9766 8658 9818
rect 8670 9766 8722 9818
rect 13475 9766 13527 9818
rect 13539 9766 13591 9818
rect 13603 9766 13655 9818
rect 13667 9766 13719 9818
rect 7012 9664 7064 9716
rect 7288 9664 7340 9716
rect 7472 9596 7524 9648
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 8300 9528 8352 9580
rect 9036 9528 9088 9580
rect 7104 9460 7156 9512
rect 9128 9460 9180 9512
rect 9680 9460 9732 9512
rect 5448 9392 5500 9444
rect 8116 9392 8168 9444
rect 8852 9392 8904 9444
rect 1584 9324 1636 9376
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 9956 9392 10008 9444
rect 12900 9324 12952 9376
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 10976 9222 11028 9274
rect 11040 9222 11092 9274
rect 11104 9222 11156 9274
rect 11168 9222 11220 9274
rect 6920 9120 6972 9172
rect 8944 8984 8996 9036
rect 13360 8984 13412 9036
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 11336 8916 11388 8968
rect 4160 8780 4212 8832
rect 13360 8780 13412 8832
rect 3480 8678 3532 8730
rect 3544 8678 3596 8730
rect 3608 8678 3660 8730
rect 3672 8678 3724 8730
rect 8478 8678 8530 8730
rect 8542 8678 8594 8730
rect 8606 8678 8658 8730
rect 8670 8678 8722 8730
rect 13475 8678 13527 8730
rect 13539 8678 13591 8730
rect 13603 8678 13655 8730
rect 13667 8678 13719 8730
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 10976 8134 11028 8186
rect 11040 8134 11092 8186
rect 11104 8134 11156 8186
rect 11168 8134 11220 8186
rect 3480 7590 3532 7642
rect 3544 7590 3596 7642
rect 3608 7590 3660 7642
rect 3672 7590 3724 7642
rect 8478 7590 8530 7642
rect 8542 7590 8594 7642
rect 8606 7590 8658 7642
rect 8670 7590 8722 7642
rect 13475 7590 13527 7642
rect 13539 7590 13591 7642
rect 13603 7590 13655 7642
rect 13667 7590 13719 7642
rect 4160 7284 4212 7336
rect 2964 7216 3016 7268
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 10976 7046 11028 7098
rect 11040 7046 11092 7098
rect 11104 7046 11156 7098
rect 11168 7046 11220 7098
rect 3976 6672 4028 6724
rect 7288 6672 7340 6724
rect 5632 6604 5684 6656
rect 9680 6604 9732 6656
rect 3480 6502 3532 6554
rect 3544 6502 3596 6554
rect 3608 6502 3660 6554
rect 3672 6502 3724 6554
rect 8478 6502 8530 6554
rect 8542 6502 8594 6554
rect 8606 6502 8658 6554
rect 8670 6502 8722 6554
rect 13475 6502 13527 6554
rect 13539 6502 13591 6554
rect 13603 6502 13655 6554
rect 13667 6502 13719 6554
rect 6920 6400 6972 6452
rect 7840 6400 7892 6452
rect 7932 6400 7984 6452
rect 11428 6400 11480 6452
rect 4804 6332 4856 6384
rect 9312 6332 9364 6384
rect 7564 6264 7616 6316
rect 11888 6264 11940 6316
rect 7104 6196 7156 6248
rect 7932 6196 7984 6248
rect 8852 6196 8904 6248
rect 11704 6196 11756 6248
rect 5080 6128 5132 6180
rect 7472 6128 7524 6180
rect 7840 6128 7892 6180
rect 12256 6128 12308 6180
rect 7748 6060 7800 6112
rect 8668 6060 8720 6112
rect 10692 6060 10744 6112
rect 10876 6060 10928 6112
rect 14004 6060 14056 6112
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 10976 5958 11028 6010
rect 11040 5958 11092 6010
rect 11104 5958 11156 6010
rect 11168 5958 11220 6010
rect 4436 5856 4488 5908
rect 9128 5856 9180 5908
rect 10876 5899 10928 5908
rect 10876 5865 10885 5899
rect 10885 5865 10919 5899
rect 10919 5865 10928 5899
rect 10876 5856 10928 5865
rect 5080 5831 5132 5840
rect 5080 5797 5089 5831
rect 5089 5797 5123 5831
rect 5123 5797 5132 5831
rect 5080 5788 5132 5797
rect 5632 5831 5684 5840
rect 5632 5797 5641 5831
rect 5641 5797 5675 5831
rect 5675 5797 5684 5831
rect 5632 5788 5684 5797
rect 8852 5831 8904 5840
rect 7104 5720 7156 5772
rect 7564 5720 7616 5772
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 8852 5797 8861 5831
rect 8861 5797 8895 5831
rect 8895 5797 8904 5831
rect 8852 5788 8904 5797
rect 8668 5763 8720 5772
rect 8668 5729 8677 5763
rect 8677 5729 8711 5763
rect 8711 5729 8720 5763
rect 8668 5720 8720 5729
rect 9036 5763 9088 5772
rect 9036 5729 9045 5763
rect 9045 5729 9079 5763
rect 9079 5729 9088 5763
rect 9036 5720 9088 5729
rect 11520 5856 11572 5908
rect 12256 5899 12308 5908
rect 12256 5865 12265 5899
rect 12265 5865 12299 5899
rect 12299 5865 12308 5899
rect 12256 5856 12308 5865
rect 15384 5856 15436 5908
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 4896 5652 4948 5704
rect 4712 5584 4764 5636
rect 6920 5627 6972 5636
rect 6920 5593 6929 5627
rect 6929 5593 6963 5627
rect 6963 5593 6972 5627
rect 6920 5584 6972 5593
rect 7472 5584 7524 5636
rect 15292 5652 15344 5704
rect 4252 5559 4304 5568
rect 4252 5525 4261 5559
rect 4261 5525 4295 5559
rect 4295 5525 4304 5559
rect 4252 5516 4304 5525
rect 4620 5559 4672 5568
rect 4620 5525 4629 5559
rect 4629 5525 4663 5559
rect 4663 5525 4672 5559
rect 4620 5516 4672 5525
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 7656 5516 7708 5568
rect 9956 5516 10008 5568
rect 10324 5516 10376 5568
rect 11980 5584 12032 5636
rect 3480 5414 3532 5466
rect 3544 5414 3596 5466
rect 3608 5414 3660 5466
rect 3672 5414 3724 5466
rect 8478 5414 8530 5466
rect 8542 5414 8594 5466
rect 8606 5414 8658 5466
rect 8670 5414 8722 5466
rect 13475 5414 13527 5466
rect 13539 5414 13591 5466
rect 13603 5414 13655 5466
rect 13667 5414 13719 5466
rect 940 5312 992 5364
rect 2688 5244 2740 5296
rect 7288 5312 7340 5364
rect 8116 5312 8168 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 10048 5312 10100 5364
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 12900 5312 12952 5364
rect 13176 5312 13228 5364
rect 15568 5312 15620 5364
rect 5080 5108 5132 5160
rect 5632 5108 5684 5160
rect 6920 5176 6972 5228
rect 6552 5108 6604 5160
rect 7288 5176 7340 5228
rect 8300 5244 8352 5296
rect 9864 5244 9916 5296
rect 7748 5108 7800 5160
rect 7932 5151 7984 5160
rect 7932 5117 7941 5151
rect 7941 5117 7975 5151
rect 7975 5117 7984 5151
rect 7932 5108 7984 5117
rect 9680 5176 9732 5228
rect 15200 5244 15252 5296
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 9588 5151 9640 5160
rect 4160 5040 4212 5092
rect 9588 5117 9597 5151
rect 9597 5117 9631 5151
rect 9631 5117 9640 5151
rect 9588 5108 9640 5117
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 7104 4972 7156 5024
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 9772 5040 9824 5092
rect 11612 5108 11664 5160
rect 12348 5108 12400 5160
rect 16488 5176 16540 5228
rect 13176 5151 13228 5160
rect 11336 5040 11388 5092
rect 13176 5117 13185 5151
rect 13185 5117 13219 5151
rect 13219 5117 13228 5151
rect 13176 5108 13228 5117
rect 11428 5015 11480 5024
rect 11428 4981 11437 5015
rect 11437 4981 11471 5015
rect 11471 4981 11480 5015
rect 11428 4972 11480 4981
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 13820 4972 13872 4981
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 10976 4870 11028 4922
rect 11040 4870 11092 4922
rect 11104 4870 11156 4922
rect 11168 4870 11220 4922
rect 5264 4768 5316 4820
rect 8484 4768 8536 4820
rect 8668 4768 8720 4820
rect 10140 4768 10192 4820
rect 11612 4811 11664 4820
rect 11612 4777 11621 4811
rect 11621 4777 11655 4811
rect 11655 4777 11664 4811
rect 11612 4768 11664 4777
rect 13084 4768 13136 4820
rect 3884 4700 3936 4752
rect 7104 4700 7156 4752
rect 3792 4632 3844 4684
rect 8116 4700 8168 4752
rect 10784 4700 10836 4752
rect 15660 4700 15712 4752
rect 7748 4632 7800 4684
rect 8852 4632 8904 4684
rect 10416 4632 10468 4684
rect 8300 4564 8352 4616
rect 9588 4564 9640 4616
rect 13912 4564 13964 4616
rect 2504 4496 2556 4548
rect 7012 4496 7064 4548
rect 9680 4496 9732 4548
rect 10048 4496 10100 4548
rect 11060 4496 11112 4548
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 7932 4428 7984 4480
rect 8944 4428 8996 4480
rect 9404 4471 9456 4480
rect 9404 4437 9413 4471
rect 9413 4437 9447 4471
rect 9447 4437 9456 4471
rect 9404 4428 9456 4437
rect 9772 4471 9824 4480
rect 9772 4437 9781 4471
rect 9781 4437 9815 4471
rect 9815 4437 9824 4471
rect 9772 4428 9824 4437
rect 11152 4428 11204 4480
rect 12440 4428 12492 4480
rect 3480 4326 3532 4378
rect 3544 4326 3596 4378
rect 3608 4326 3660 4378
rect 3672 4326 3724 4378
rect 8478 4326 8530 4378
rect 8542 4326 8594 4378
rect 8606 4326 8658 4378
rect 8670 4326 8722 4378
rect 13475 4326 13527 4378
rect 13539 4326 13591 4378
rect 13603 4326 13655 4378
rect 13667 4326 13719 4378
rect 5264 4224 5316 4276
rect 9220 4224 9272 4276
rect 6644 4156 6696 4208
rect 10508 4156 10560 4208
rect 2780 4088 2832 4140
rect 7196 4088 7248 4140
rect 9772 4088 9824 4140
rect 13268 4088 13320 4140
rect 13820 4088 13872 4140
rect 16948 4088 17000 4140
rect 3148 4020 3200 4072
rect 7564 4020 7616 4072
rect 11060 4020 11112 4072
rect 14372 4020 14424 4072
rect 5632 3952 5684 4004
rect 9220 3952 9272 4004
rect 11152 3952 11204 4004
rect 14740 3952 14792 4004
rect 6644 3884 6696 3936
rect 11428 3884 11480 3936
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 10976 3782 11028 3834
rect 11040 3782 11092 3834
rect 11104 3782 11156 3834
rect 11168 3782 11220 3834
rect 6920 3680 6972 3732
rect 10048 3680 10100 3732
rect 7012 3612 7064 3664
rect 9404 3612 9456 3664
rect 7288 3544 7340 3596
rect 10876 3544 10928 3596
rect 4068 3476 4120 3528
rect 7656 3476 7708 3528
rect 8300 3476 8352 3528
rect 11336 3476 11388 3528
rect 8852 3408 8904 3460
rect 11796 3408 11848 3460
rect 8944 3340 8996 3392
rect 12164 3340 12216 3392
rect 3480 3238 3532 3290
rect 3544 3238 3596 3290
rect 3608 3238 3660 3290
rect 3672 3238 3724 3290
rect 8478 3238 8530 3290
rect 8542 3238 8594 3290
rect 8606 3238 8658 3290
rect 8670 3238 8722 3290
rect 13475 3238 13527 3290
rect 13539 3238 13591 3290
rect 13603 3238 13655 3290
rect 13667 3238 13719 3290
rect 2320 3136 2372 3188
rect 4712 3136 4764 3188
rect 5724 3136 5776 3188
rect 9956 3136 10008 3188
rect 12440 3136 12492 3188
rect 16028 3136 16080 3188
rect 1860 3068 1912 3120
rect 5356 3068 5408 3120
rect 7380 3068 7432 3120
rect 8852 3068 8904 3120
rect 9680 3068 9732 3120
rect 12624 3068 12676 3120
rect 1492 3000 1544 3052
rect 6368 3000 6420 3052
rect 572 2932 624 2984
rect 4988 2932 5040 2984
rect 6276 2932 6328 2984
rect 10324 2932 10376 2984
rect 204 2864 256 2916
rect 4252 2864 4304 2916
rect 1032 2796 1084 2848
rect 4620 2796 4672 2848
rect 8300 2796 8352 2848
rect 13360 2796 13412 2848
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 10976 2694 11028 2746
rect 11040 2694 11092 2746
rect 11104 2694 11156 2746
rect 11168 2694 11220 2746
rect 3480 2150 3532 2202
rect 3544 2150 3596 2202
rect 3608 2150 3660 2202
rect 3672 2150 3724 2202
rect 8478 2150 8530 2202
rect 8542 2150 8594 2202
rect 8606 2150 8658 2202
rect 8670 2150 8722 2202
rect 13475 2150 13527 2202
rect 13539 2150 13591 2202
rect 13603 2150 13655 2202
rect 13667 2150 13719 2202
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1858 19200 1914 20000
rect 2226 19200 2282 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3514 19200 3570 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4802 19200 4858 20000
rect 5170 19200 5226 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6458 19200 6514 20000
rect 6826 19200 6882 20000
rect 7286 19200 7342 20000
rect 7746 19200 7802 20000
rect 8114 19200 8170 20000
rect 8574 19200 8630 20000
rect 8942 19200 8998 20000
rect 9402 19200 9458 20000
rect 9770 19200 9826 20000
rect 10230 19200 10286 20000
rect 10690 19200 10746 20000
rect 11058 19200 11114 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12346 19200 12402 20000
rect 12714 19200 12770 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 14002 19200 14058 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15290 19200 15346 20000
rect 15658 19200 15714 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16946 19200 17002 20000
rect 216 15434 244 19200
rect 204 15428 256 15434
rect 204 15370 256 15376
rect 584 15162 612 19200
rect 572 15156 624 15162
rect 572 15098 624 15104
rect 1044 12458 1072 19200
rect 1412 15502 1440 19200
rect 1872 15706 1900 19200
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 2240 15570 2268 19200
rect 2700 15994 2728 19200
rect 2516 15966 2728 15994
rect 2228 15564 2280 15570
rect 2228 15506 2280 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 952 12430 1072 12458
rect 952 5370 980 12430
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 10198 1532 10542
rect 1492 10192 1544 10198
rect 1492 10134 1544 10140
rect 1504 8401 1532 10134
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1596 9382 1624 9998
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1490 8392 1546 8401
rect 1490 8327 1546 8336
rect 940 5364 992 5370
rect 940 5306 992 5312
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 800 244 2858
rect 584 800 612 2926
rect 1032 2848 1084 2854
rect 1032 2790 1084 2796
rect 1044 800 1072 2790
rect 1504 800 1532 2994
rect 1596 1737 1624 9318
rect 2516 4554 2544 15966
rect 3068 15706 3096 19200
rect 3528 17626 3556 19200
rect 3528 17598 3924 17626
rect 3454 17436 3750 17456
rect 3510 17434 3534 17436
rect 3590 17434 3614 17436
rect 3670 17434 3694 17436
rect 3532 17382 3534 17434
rect 3596 17382 3608 17434
rect 3670 17382 3672 17434
rect 3510 17380 3534 17382
rect 3590 17380 3614 17382
rect 3670 17380 3694 17382
rect 3454 17360 3750 17380
rect 3454 16348 3750 16368
rect 3510 16346 3534 16348
rect 3590 16346 3614 16348
rect 3670 16346 3694 16348
rect 3532 16294 3534 16346
rect 3596 16294 3608 16346
rect 3670 16294 3672 16346
rect 3510 16292 3534 16294
rect 3590 16292 3614 16294
rect 3670 16292 3694 16294
rect 3454 16272 3750 16292
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2700 5302 2728 15642
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2778 15056 2834 15065
rect 2778 14991 2834 15000
rect 2792 10198 2820 14991
rect 2884 13530 2912 15370
rect 3454 15260 3750 15280
rect 3510 15258 3534 15260
rect 3590 15258 3614 15260
rect 3670 15258 3694 15260
rect 3532 15206 3534 15258
rect 3596 15206 3608 15258
rect 3670 15206 3672 15258
rect 3510 15204 3534 15206
rect 3590 15204 3614 15206
rect 3670 15204 3694 15206
rect 3454 15184 3750 15204
rect 3454 14172 3750 14192
rect 3510 14170 3534 14172
rect 3590 14170 3614 14172
rect 3670 14170 3694 14172
rect 3532 14118 3534 14170
rect 3596 14118 3608 14170
rect 3670 14118 3672 14170
rect 3510 14116 3534 14118
rect 3590 14116 3614 14118
rect 3670 14116 3694 14118
rect 3454 14096 3750 14116
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 10606 3280 13126
rect 3454 13084 3750 13104
rect 3510 13082 3534 13084
rect 3590 13082 3614 13084
rect 3670 13082 3694 13084
rect 3532 13030 3534 13082
rect 3596 13030 3608 13082
rect 3670 13030 3672 13082
rect 3510 13028 3534 13030
rect 3590 13028 3614 13030
rect 3670 13028 3694 13030
rect 3454 13008 3750 13028
rect 3454 11996 3750 12016
rect 3510 11994 3534 11996
rect 3590 11994 3614 11996
rect 3670 11994 3694 11996
rect 3532 11942 3534 11994
rect 3596 11942 3608 11994
rect 3670 11942 3672 11994
rect 3510 11940 3534 11942
rect 3590 11940 3614 11942
rect 3670 11940 3694 11942
rect 3454 11920 3750 11940
rect 3330 11656 3386 11665
rect 3330 11591 3386 11600
rect 3344 10810 3372 11591
rect 3454 10908 3750 10928
rect 3510 10906 3534 10908
rect 3590 10906 3614 10908
rect 3670 10906 3694 10908
rect 3532 10854 3534 10906
rect 3596 10854 3608 10906
rect 3670 10854 3672 10906
rect 3510 10852 3534 10854
rect 3590 10852 3614 10854
rect 3670 10852 3694 10854
rect 3454 10832 3750 10852
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 3454 9820 3750 9840
rect 3510 9818 3534 9820
rect 3590 9818 3614 9820
rect 3670 9818 3694 9820
rect 3532 9766 3534 9818
rect 3596 9766 3608 9818
rect 3670 9766 3672 9818
rect 3510 9764 3534 9766
rect 3590 9764 3614 9766
rect 3670 9764 3694 9766
rect 3454 9744 3750 9764
rect 3454 8732 3750 8752
rect 3510 8730 3534 8732
rect 3590 8730 3614 8732
rect 3670 8730 3694 8732
rect 3532 8678 3534 8730
rect 3596 8678 3608 8730
rect 3670 8678 3672 8730
rect 3510 8676 3534 8678
rect 3590 8676 3614 8678
rect 3670 8676 3694 8678
rect 3454 8656 3750 8676
rect 3454 7644 3750 7664
rect 3510 7642 3534 7644
rect 3590 7642 3614 7644
rect 3670 7642 3694 7644
rect 3532 7590 3534 7642
rect 3596 7590 3608 7642
rect 3670 7590 3672 7642
rect 3510 7588 3534 7590
rect 3590 7588 3614 7590
rect 3670 7588 3694 7590
rect 3454 7568 3750 7588
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2688 5296 2740 5302
rect 2688 5238 2740 5244
rect 2976 5001 3004 7210
rect 3454 6556 3750 6576
rect 3510 6554 3534 6556
rect 3590 6554 3614 6556
rect 3670 6554 3694 6556
rect 3532 6502 3534 6554
rect 3596 6502 3608 6554
rect 3670 6502 3672 6554
rect 3510 6500 3534 6502
rect 3590 6500 3614 6502
rect 3670 6500 3694 6502
rect 3454 6480 3750 6500
rect 3454 5468 3750 5488
rect 3510 5466 3534 5468
rect 3590 5466 3614 5468
rect 3670 5466 3694 5468
rect 3532 5414 3534 5466
rect 3596 5414 3608 5466
rect 3670 5414 3672 5466
rect 3510 5412 3534 5414
rect 3590 5412 3614 5414
rect 3670 5412 3694 5414
rect 3454 5392 3750 5412
rect 2962 4992 3018 5001
rect 2962 4927 3018 4936
rect 3804 4690 3832 15846
rect 3896 4758 3924 17598
rect 3988 15910 4016 19200
rect 4066 18320 4122 18329
rect 4066 18255 4122 18264
rect 3976 15904 4028 15910
rect 3976 15846 4028 15852
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3988 6730 4016 15642
rect 4080 14074 4108 18255
rect 4356 15910 4384 19200
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4724 15162 4752 15438
rect 4816 15366 4844 19200
rect 5184 19122 5212 19200
rect 5184 19094 5304 19122
rect 5276 17950 5304 19094
rect 5264 17944 5316 17950
rect 5264 17886 5316 17892
rect 5448 17944 5500 17950
rect 5448 17886 5500 17892
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4356 13530 4384 13806
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 7342 4200 8774
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 3454 4380 3750 4400
rect 3510 4378 3534 4380
rect 3590 4378 3614 4380
rect 3670 4378 3694 4380
rect 3532 4326 3534 4378
rect 3596 4326 3608 4378
rect 3670 4326 3672 4378
rect 3510 4324 3534 4326
rect 3590 4324 3614 4326
rect 3670 4324 3694 4326
rect 3454 4304 3750 4324
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1582 1728 1638 1737
rect 1582 1663 1638 1672
rect 1872 800 1900 3062
rect 2332 800 2360 3130
rect 2792 800 2820 4082
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3160 800 3188 4014
rect 4172 3890 4200 5034
rect 3804 3862 4200 3890
rect 3454 3292 3750 3312
rect 3510 3290 3534 3292
rect 3590 3290 3614 3292
rect 3670 3290 3694 3292
rect 3532 3238 3534 3290
rect 3596 3238 3608 3290
rect 3670 3238 3672 3290
rect 3510 3236 3534 3238
rect 3590 3236 3614 3238
rect 3670 3236 3694 3238
rect 3454 3216 3750 3236
rect 3454 2204 3750 2224
rect 3510 2202 3534 2204
rect 3590 2202 3614 2204
rect 3670 2202 3694 2204
rect 3532 2150 3534 2202
rect 3596 2150 3608 2202
rect 3670 2150 3672 2202
rect 3510 2148 3534 2150
rect 3590 2148 3614 2150
rect 3670 2148 3694 2150
rect 3454 2128 3750 2148
rect 3804 1986 3832 3862
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3620 1958 3832 1986
rect 3620 800 3648 1958
rect 4080 800 4108 3470
rect 4264 2922 4292 5510
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4448 800 4476 5850
rect 4816 5710 4844 6326
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5846 5120 6122
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4896 5704 4948 5710
rect 5368 5658 5396 15846
rect 5460 9450 5488 17886
rect 5644 15978 5672 19200
rect 6012 17082 6040 19200
rect 6012 17054 6316 17082
rect 5953 16892 6249 16912
rect 6009 16890 6033 16892
rect 6089 16890 6113 16892
rect 6169 16890 6193 16892
rect 6031 16838 6033 16890
rect 6095 16838 6107 16890
rect 6169 16838 6171 16890
rect 6009 16836 6033 16838
rect 6089 16836 6113 16838
rect 6169 16836 6193 16838
rect 5953 16816 6249 16836
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5953 15804 6249 15824
rect 6009 15802 6033 15804
rect 6089 15802 6113 15804
rect 6169 15802 6193 15804
rect 6031 15750 6033 15802
rect 6095 15750 6107 15802
rect 6169 15750 6171 15802
rect 6009 15748 6033 15750
rect 6089 15748 6113 15750
rect 6169 15748 6193 15750
rect 5953 15728 6249 15748
rect 6288 15638 6316 17054
rect 6472 16114 6500 19200
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 15162 5580 15506
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5552 10742 5580 14962
rect 5953 14716 6249 14736
rect 6009 14714 6033 14716
rect 6089 14714 6113 14716
rect 6169 14714 6193 14716
rect 6031 14662 6033 14714
rect 6095 14662 6107 14714
rect 6169 14662 6171 14714
rect 6009 14660 6033 14662
rect 6089 14660 6113 14662
rect 6169 14660 6193 14662
rect 5953 14640 6249 14660
rect 6748 14618 6776 15302
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 11626 5764 13670
rect 5953 13628 6249 13648
rect 6009 13626 6033 13628
rect 6089 13626 6113 13628
rect 6169 13626 6193 13628
rect 6031 13574 6033 13626
rect 6095 13574 6107 13626
rect 6169 13574 6171 13626
rect 6009 13572 6033 13574
rect 6089 13572 6113 13574
rect 6169 13572 6193 13574
rect 5953 13552 6249 13572
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 5953 12540 6249 12560
rect 6009 12538 6033 12540
rect 6089 12538 6113 12540
rect 6169 12538 6193 12540
rect 6031 12486 6033 12538
rect 6095 12486 6107 12538
rect 6169 12486 6171 12538
rect 6009 12484 6033 12486
rect 6089 12484 6113 12486
rect 6169 12484 6193 12486
rect 5953 12464 6249 12484
rect 6288 12442 6316 13330
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5953 11452 6249 11472
rect 6009 11450 6033 11452
rect 6089 11450 6113 11452
rect 6169 11450 6193 11452
rect 6031 11398 6033 11450
rect 6095 11398 6107 11450
rect 6169 11398 6171 11450
rect 6009 11396 6033 11398
rect 6089 11396 6113 11398
rect 6169 11396 6193 11398
rect 5953 11376 6249 11396
rect 6748 11286 6776 12378
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5953 10364 6249 10384
rect 6009 10362 6033 10364
rect 6089 10362 6113 10364
rect 6169 10362 6193 10364
rect 6031 10310 6033 10362
rect 6095 10310 6107 10362
rect 6169 10310 6171 10362
rect 6009 10308 6033 10310
rect 6089 10308 6113 10310
rect 6169 10308 6193 10310
rect 5953 10288 6249 10308
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5953 9276 6249 9296
rect 6009 9274 6033 9276
rect 6089 9274 6113 9276
rect 6169 9274 6193 9276
rect 6031 9222 6033 9274
rect 6095 9222 6107 9274
rect 6169 9222 6171 9274
rect 6009 9220 6033 9222
rect 6089 9220 6113 9222
rect 6169 9220 6193 9222
rect 5953 9200 6249 9220
rect 5953 8188 6249 8208
rect 6009 8186 6033 8188
rect 6089 8186 6113 8188
rect 6169 8186 6193 8188
rect 6031 8134 6033 8186
rect 6095 8134 6107 8186
rect 6169 8134 6171 8186
rect 6009 8132 6033 8134
rect 6089 8132 6113 8134
rect 6169 8132 6193 8134
rect 5953 8112 6249 8132
rect 5953 7100 6249 7120
rect 6009 7098 6033 7100
rect 6089 7098 6113 7100
rect 6169 7098 6193 7100
rect 6031 7046 6033 7098
rect 6095 7046 6107 7098
rect 6169 7046 6171 7098
rect 6009 7044 6033 7046
rect 6089 7044 6113 7046
rect 6169 7044 6193 7046
rect 5953 7024 6249 7044
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5644 5846 5672 6598
rect 5953 6012 6249 6032
rect 6009 6010 6033 6012
rect 6089 6010 6113 6012
rect 6169 6010 6193 6012
rect 6031 5958 6033 6010
rect 6095 5958 6107 6010
rect 6169 5958 6171 6010
rect 6009 5956 6033 5958
rect 6089 5956 6113 5958
rect 6169 5956 6193 5958
rect 5953 5936 6249 5956
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 4896 5646 4948 5652
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4632 2854 4660 5510
rect 4724 3194 4752 5578
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4908 800 4936 5646
rect 5276 5630 5396 5658
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5000 2990 5028 4966
rect 5092 4468 5120 5102
rect 5276 4826 5304 5630
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5264 4480 5316 4486
rect 5092 4440 5264 4468
rect 5264 4422 5316 4428
rect 5276 4282 5304 4422
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5368 3126 5396 5510
rect 6840 5273 6868 19200
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7024 10266 7052 11018
rect 7116 10606 7144 15982
rect 7300 15366 7328 19200
rect 7760 15910 7788 19200
rect 8128 19122 8156 19200
rect 8128 19094 8248 19122
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7196 15088 7248 15094
rect 7196 15030 7248 15036
rect 7208 11558 7236 15030
rect 7472 11688 7524 11694
rect 7524 11636 7604 11642
rect 7472 11630 7604 11636
rect 7288 11620 7340 11626
rect 7484 11614 7604 11630
rect 7288 11562 7340 11568
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7300 11014 7328 11562
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11234 7512 11494
rect 7392 11218 7512 11234
rect 7380 11212 7512 11218
rect 7432 11206 7512 11212
rect 7380 11154 7432 11160
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7208 10470 7236 10678
rect 7300 10674 7328 10950
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9178 6960 9862
rect 7024 9722 7052 9998
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7116 9518 7144 10406
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 7208 8974 7236 9862
rect 7300 9722 7328 10066
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6932 5642 6960 6394
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7116 5778 7144 6190
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6826 5264 6882 5273
rect 6826 5199 6882 5208
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 6552 5160 6604 5166
rect 6604 5108 6684 5114
rect 6552 5102 6684 5108
rect 5644 5030 5672 5102
rect 6564 5086 6684 5102
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 5644 4010 5672 4966
rect 5953 4924 6249 4944
rect 6009 4922 6033 4924
rect 6089 4922 6113 4924
rect 6169 4922 6193 4924
rect 6031 4870 6033 4922
rect 6095 4870 6107 4922
rect 6169 4870 6171 4922
rect 6009 4868 6033 4870
rect 6089 4868 6113 4870
rect 6169 4868 6193 4870
rect 5953 4848 6249 4868
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5953 3836 6249 3856
rect 6009 3834 6033 3836
rect 6089 3834 6113 3836
rect 6169 3834 6193 3836
rect 6031 3782 6033 3834
rect 6095 3782 6107 3834
rect 6169 3782 6171 3834
rect 6009 3780 6033 3782
rect 6089 3780 6113 3782
rect 6169 3780 6193 3782
rect 5953 3760 6249 3780
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5354 912 5410 921
rect 5354 847 5410 856
rect 5368 800 5396 847
rect 5736 800 5764 3130
rect 6380 3058 6408 4966
rect 6656 4486 6684 5086
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6656 4214 6684 4422
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 5953 2748 6249 2768
rect 6009 2746 6033 2748
rect 6089 2746 6113 2748
rect 6169 2746 6193 2748
rect 6031 2694 6033 2746
rect 6095 2694 6107 2746
rect 6169 2694 6171 2746
rect 6009 2692 6033 2694
rect 6089 2692 6113 2694
rect 6169 2692 6193 2694
rect 5953 2672 6249 2692
rect 6288 1850 6316 2926
rect 6196 1822 6316 1850
rect 6196 800 6224 1822
rect 6656 800 6684 3878
rect 6932 3738 6960 5170
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7024 4554 7052 4966
rect 7116 4758 7144 4966
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7208 4146 7236 5510
rect 7300 5370 7328 6666
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7300 4486 7328 5170
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7024 800 7052 3606
rect 7300 3602 7328 4422
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7392 3126 7420 11154
rect 7576 11082 7604 11614
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 7576 10674 7604 11018
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 7484 9654 7512 10542
rect 7576 10418 7604 10610
rect 7576 10390 7696 10418
rect 7668 10266 7696 10390
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7484 6186 7512 9590
rect 7576 9586 7604 10202
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7852 6458 7880 16526
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8128 9926 8156 11154
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7576 5778 7604 6258
rect 7944 6254 7972 6394
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7840 6180 7892 6186
rect 7840 6122 7892 6128
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5778 7788 6054
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7484 800 7512 5578
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7576 4078 7604 5510
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7668 3534 7696 5510
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7760 4690 7788 5102
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7852 898 7880 6122
rect 8128 5370 8156 9386
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7932 5160 7984 5166
rect 8220 5137 8248 19094
rect 8588 17626 8616 19200
rect 8588 17598 8892 17626
rect 8452 17436 8748 17456
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8530 17382 8532 17434
rect 8594 17382 8606 17434
rect 8668 17382 8670 17434
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8452 17360 8748 17380
rect 8452 16348 8748 16368
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8530 16294 8532 16346
rect 8594 16294 8606 16346
rect 8668 16294 8670 16346
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8452 16272 8748 16292
rect 8864 15570 8892 17598
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8452 15260 8748 15280
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8530 15206 8532 15258
rect 8594 15206 8606 15258
rect 8668 15206 8670 15258
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8452 15184 8748 15204
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8452 14172 8748 14192
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8530 14118 8532 14170
rect 8594 14118 8606 14170
rect 8668 14118 8670 14170
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8452 14096 8748 14116
rect 8452 13084 8748 13104
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8530 13030 8532 13082
rect 8594 13030 8606 13082
rect 8668 13030 8670 13082
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8452 13008 8748 13028
rect 8452 11996 8748 12016
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8530 11942 8532 11994
rect 8594 11942 8606 11994
rect 8668 11942 8670 11994
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8452 11920 8748 11940
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 10538 8340 11494
rect 8452 10908 8748 10928
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8530 10854 8532 10906
rect 8594 10854 8606 10906
rect 8668 10854 8670 10906
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8452 10832 8748 10852
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8312 10198 8340 10474
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8312 9586 8340 10134
rect 8452 9820 8748 9840
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8530 9766 8532 9818
rect 8594 9766 8606 9818
rect 8668 9766 8670 9818
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8452 9744 8748 9764
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8864 9450 8892 14214
rect 8956 11286 8984 19200
rect 9416 15858 9444 19200
rect 9784 16046 9812 19200
rect 10244 19145 10272 19200
rect 10230 19136 10286 19145
rect 10230 19071 10286 19080
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9232 15830 9444 15858
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 9048 10554 9076 15642
rect 8956 10526 9076 10554
rect 8956 9466 8984 10526
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9048 10130 9076 10406
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9048 9586 9076 10066
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9140 9518 9168 10406
rect 9128 9512 9180 9518
rect 8852 9444 8904 9450
rect 8956 9438 9076 9466
rect 9128 9454 9180 9460
rect 8852 9386 8904 9392
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 9042 8984 9318
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8452 8732 8748 8752
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8530 8678 8532 8730
rect 8594 8678 8606 8730
rect 8668 8678 8670 8730
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8452 8656 8748 8676
rect 8452 7644 8748 7664
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8530 7590 8532 7642
rect 8594 7590 8606 7642
rect 8668 7590 8670 7642
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8452 7568 8748 7588
rect 8452 6556 8748 6576
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8530 6502 8532 6554
rect 8594 6502 8606 6554
rect 8668 6502 8670 6554
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8452 6480 8748 6500
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5778 8708 6054
rect 8864 5846 8892 6190
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 9048 5778 9076 9438
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 9036 5772 9088 5778
rect 9036 5714 9088 5720
rect 8452 5468 8748 5488
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8530 5414 8532 5466
rect 8594 5414 8606 5466
rect 8668 5414 8670 5466
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8452 5392 8748 5412
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 7932 5102 7984 5108
rect 8206 5128 8262 5137
rect 7944 4486 7972 5102
rect 8206 5063 8262 5072
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8128 4758 8156 4966
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8312 4622 8340 5238
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4826 8524 4966
rect 8680 4826 8708 5102
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 8312 3534 8340 4558
rect 8452 4380 8748 4400
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8530 4326 8532 4378
rect 8594 4326 8606 4378
rect 8668 4326 8670 4378
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8452 4304 8748 4324
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8864 3466 8892 4626
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8956 3398 8984 4422
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8452 3292 8748 3312
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8530 3238 8532 3290
rect 8594 3238 8606 3290
rect 8668 3238 8670 3290
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8452 3216 8748 3236
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7852 870 7972 898
rect 7944 800 7972 870
rect 8312 800 8340 2790
rect 8452 2204 8748 2224
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8530 2150 8532 2202
rect 8594 2150 8606 2202
rect 8668 2150 8670 2202
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8452 2128 8748 2148
rect 8864 1986 8892 3062
rect 8772 1958 8892 1986
rect 8772 800 8800 1958
rect 9140 921 9168 5850
rect 9232 4282 9260 15830
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12646 9352 13262
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 11354 9352 12582
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9324 6390 9352 11154
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9416 5409 9444 15506
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9600 14618 9628 15302
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9508 10470 9536 10950
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 9625 9536 10406
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9494 9616 9550 9625
rect 9494 9551 9550 9560
rect 9600 9489 9628 10202
rect 9692 10010 9720 15914
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 9784 10146 9812 15846
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 11286 9904 14758
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 10538 9904 11222
rect 9968 10554 9996 15574
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 14278 10088 14418
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 10674 10088 14214
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9864 10532 9916 10538
rect 9968 10526 10088 10554
rect 9864 10474 9916 10480
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9784 10118 9904 10146
rect 9692 9982 9812 10010
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9518 9720 9862
rect 9680 9512 9732 9518
rect 9586 9480 9642 9489
rect 9680 9454 9732 9460
rect 9586 9415 9642 9424
rect 9586 9344 9642 9353
rect 9642 9302 9720 9330
rect 9586 9279 9642 9288
rect 9692 6662 9720 9302
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9402 5400 9458 5409
rect 9784 5370 9812 9982
rect 9402 5335 9458 5344
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9876 5302 9904 10118
rect 9968 9450 9996 10406
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 4622 9628 5102
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9692 4554 9720 5170
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9126 912 9182 921
rect 9126 847 9182 856
rect 9232 800 9260 3946
rect 9416 3670 9444 4422
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9692 3126 9720 4490
rect 9784 4486 9812 5034
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 4146 9812 4422
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9968 3194 9996 5510
rect 10060 5370 10088 10526
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10060 4554 10088 5102
rect 10152 4826 10180 15846
rect 10612 10962 10640 16050
rect 10704 11286 10732 19200
rect 11072 17082 11100 19200
rect 10888 17054 11100 17082
rect 10888 16590 10916 17054
rect 10950 16892 11246 16912
rect 11006 16890 11030 16892
rect 11086 16890 11110 16892
rect 11166 16890 11190 16892
rect 11028 16838 11030 16890
rect 11092 16838 11104 16890
rect 11166 16838 11168 16890
rect 11006 16836 11030 16838
rect 11086 16836 11110 16838
rect 11166 16836 11190 16838
rect 10950 16816 11246 16836
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10950 15804 11246 15824
rect 11006 15802 11030 15804
rect 11086 15802 11110 15804
rect 11166 15802 11190 15804
rect 11028 15750 11030 15802
rect 11092 15750 11104 15802
rect 11166 15750 11168 15802
rect 11006 15748 11030 15750
rect 11086 15748 11110 15750
rect 11166 15748 11190 15750
rect 10950 15728 11246 15748
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10612 10934 10732 10962
rect 10704 10724 10732 10934
rect 10612 10696 10732 10724
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10244 9625 10272 10474
rect 10336 9994 10364 10610
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9586 912 9642 921
rect 9586 847 9642 856
rect 9600 800 9628 847
rect 10060 800 10088 3674
rect 10336 2990 10364 5510
rect 10428 4690 10456 10406
rect 10520 10198 10548 10610
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10506 10024 10562 10033
rect 10506 9959 10562 9968
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10520 4214 10548 9959
rect 10612 5370 10640 10696
rect 10796 10266 10824 15574
rect 10950 14716 11246 14736
rect 11006 14714 11030 14716
rect 11086 14714 11110 14716
rect 11166 14714 11190 14716
rect 11028 14662 11030 14714
rect 11092 14662 11104 14714
rect 11166 14662 11168 14714
rect 11006 14660 11030 14662
rect 11086 14660 11110 14662
rect 11166 14660 11190 14662
rect 10950 14640 11246 14660
rect 11532 14600 11560 19200
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11532 14572 11652 14600
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 10950 13628 11246 13648
rect 11006 13626 11030 13628
rect 11086 13626 11110 13628
rect 11166 13626 11190 13628
rect 11028 13574 11030 13626
rect 11092 13574 11104 13626
rect 11166 13574 11168 13626
rect 11006 13572 11030 13574
rect 11086 13572 11110 13574
rect 11166 13572 11190 13574
rect 10950 13552 11246 13572
rect 10950 12540 11246 12560
rect 11006 12538 11030 12540
rect 11086 12538 11110 12540
rect 11166 12538 11190 12540
rect 11028 12486 11030 12538
rect 11092 12486 11104 12538
rect 11166 12486 11168 12538
rect 11006 12484 11030 12486
rect 11086 12484 11110 12486
rect 11166 12484 11190 12486
rect 10950 12464 11246 12484
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10950 11452 11246 11472
rect 11006 11450 11030 11452
rect 11086 11450 11110 11452
rect 11166 11450 11190 11452
rect 11028 11398 11030 11450
rect 11092 11398 11104 11450
rect 11166 11398 11168 11450
rect 11006 11396 11030 11398
rect 11086 11396 11110 11398
rect 11166 11396 11190 11398
rect 10950 11376 11246 11396
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10470 10916 10746
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10950 10364 11246 10384
rect 11006 10362 11030 10364
rect 11086 10362 11110 10364
rect 11166 10362 11190 10364
rect 11028 10310 11030 10362
rect 11092 10310 11104 10362
rect 11166 10310 11168 10362
rect 11006 10308 11030 10310
rect 11086 10308 11110 10310
rect 11166 10308 11190 10310
rect 10950 10288 11246 10308
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10796 10010 10824 10202
rect 10704 9982 10824 10010
rect 10704 6118 10732 9982
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10796 4758 10824 9862
rect 10950 9276 11246 9296
rect 11006 9274 11030 9276
rect 11086 9274 11110 9276
rect 11166 9274 11190 9276
rect 11028 9222 11030 9274
rect 11092 9222 11104 9274
rect 11166 9222 11168 9274
rect 11006 9220 11030 9222
rect 11086 9220 11110 9222
rect 11166 9220 11190 9222
rect 10950 9200 11246 9220
rect 11348 8974 11376 12242
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 10950 8188 11246 8208
rect 11006 8186 11030 8188
rect 11086 8186 11110 8188
rect 11166 8186 11190 8188
rect 11028 8134 11030 8186
rect 11092 8134 11104 8186
rect 11166 8134 11168 8186
rect 11006 8132 11030 8134
rect 11086 8132 11110 8134
rect 11166 8132 11190 8134
rect 10950 8112 11246 8132
rect 10950 7100 11246 7120
rect 11006 7098 11030 7100
rect 11086 7098 11110 7100
rect 11166 7098 11190 7100
rect 11028 7046 11030 7098
rect 11092 7046 11104 7098
rect 11166 7046 11168 7098
rect 11006 7044 11030 7046
rect 11086 7044 11110 7046
rect 11166 7044 11190 7046
rect 10950 7024 11246 7044
rect 11440 6458 11468 12378
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5914 10916 6054
rect 10950 6012 11246 6032
rect 11006 6010 11030 6012
rect 11086 6010 11110 6012
rect 11166 6010 11190 6012
rect 11028 5958 11030 6010
rect 11092 5958 11104 6010
rect 11166 5958 11168 6010
rect 11006 5956 11030 5958
rect 11086 5956 11110 5958
rect 11166 5956 11190 5958
rect 10950 5936 11246 5956
rect 11532 5914 11560 14418
rect 11624 12442 11652 14572
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11716 6254 11744 15302
rect 11900 6322 11928 19200
rect 12360 15910 12388 19200
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11992 5642 12020 15370
rect 12728 15366 12756 19200
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12268 5914 12296 6122
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 12912 5522 12940 9318
rect 12912 5494 13032 5522
rect 12898 5400 12954 5409
rect 11060 5364 11112 5370
rect 12898 5335 12900 5344
rect 11060 5306 11112 5312
rect 12952 5335 12954 5344
rect 12900 5306 12952 5312
rect 11072 5273 11100 5306
rect 11058 5264 11114 5273
rect 11058 5199 11114 5208
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 12348 5160 12400 5166
rect 12622 5128 12678 5137
rect 12400 5108 12480 5114
rect 12348 5102 12480 5108
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 10950 4924 11246 4944
rect 11006 4922 11030 4924
rect 11086 4922 11110 4924
rect 11166 4922 11190 4924
rect 11028 4870 11030 4922
rect 11092 4870 11104 4922
rect 11166 4870 11168 4922
rect 11006 4868 11030 4870
rect 11086 4868 11110 4870
rect 11166 4868 11190 4870
rect 10950 4848 11246 4868
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 11072 4078 11100 4490
rect 11152 4480 11204 4486
rect 11348 4468 11376 5034
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11204 4440 11376 4468
rect 11152 4422 11204 4428
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 11164 4010 11192 4422
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11440 3942 11468 4966
rect 11624 4826 11652 5102
rect 12360 5086 12480 5102
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 12452 4486 12480 5086
rect 12622 5063 12678 5072
rect 12636 5030 12664 5063
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 10950 3836 11246 3856
rect 11006 3834 11030 3836
rect 11086 3834 11110 3836
rect 11166 3834 11190 3836
rect 11028 3782 11030 3834
rect 11092 3782 11104 3834
rect 11166 3782 11168 3834
rect 11006 3780 11030 3782
rect 11086 3780 11110 3782
rect 11166 3780 11190 3782
rect 10950 3760 11246 3780
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 10506 912 10562 921
rect 10506 847 10562 856
rect 10520 800 10548 847
rect 10888 800 10916 3538
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 10950 2748 11246 2768
rect 11006 2746 11030 2748
rect 11086 2746 11110 2748
rect 11166 2746 11190 2748
rect 11028 2694 11030 2746
rect 11092 2694 11104 2746
rect 11166 2694 11168 2746
rect 11006 2692 11030 2694
rect 11086 2692 11110 2694
rect 11166 2692 11190 2694
rect 10950 2672 11246 2692
rect 11348 800 11376 3470
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11808 800 11836 3402
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12176 800 12204 3334
rect 12452 3194 12480 4422
rect 13004 3482 13032 5494
rect 13096 4826 13124 15914
rect 13188 15638 13216 19200
rect 13556 17626 13584 19200
rect 13372 17598 13584 17626
rect 13372 15706 13400 17598
rect 13449 17436 13745 17456
rect 13505 17434 13529 17436
rect 13585 17434 13609 17436
rect 13665 17434 13689 17436
rect 13527 17382 13529 17434
rect 13591 17382 13603 17434
rect 13665 17382 13667 17434
rect 13505 17380 13529 17382
rect 13585 17380 13609 17382
rect 13665 17380 13689 17382
rect 13449 17360 13745 17380
rect 13449 16348 13745 16368
rect 13505 16346 13529 16348
rect 13585 16346 13609 16348
rect 13665 16346 13689 16348
rect 13527 16294 13529 16346
rect 13591 16294 13603 16346
rect 13665 16294 13667 16346
rect 13505 16292 13529 16294
rect 13585 16292 13609 16294
rect 13665 16292 13689 16294
rect 13449 16272 13745 16292
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13449 15260 13745 15280
rect 13505 15258 13529 15260
rect 13585 15258 13609 15260
rect 13665 15258 13689 15260
rect 13527 15206 13529 15258
rect 13591 15206 13603 15258
rect 13665 15206 13667 15258
rect 13505 15204 13529 15206
rect 13585 15204 13609 15206
rect 13665 15204 13689 15206
rect 13449 15184 13745 15204
rect 13449 14172 13745 14192
rect 13505 14170 13529 14172
rect 13585 14170 13609 14172
rect 13665 14170 13689 14172
rect 13527 14118 13529 14170
rect 13591 14118 13603 14170
rect 13665 14118 13667 14170
rect 13505 14116 13529 14118
rect 13585 14116 13609 14118
rect 13665 14116 13689 14118
rect 13449 14096 13745 14116
rect 13449 13084 13745 13104
rect 13505 13082 13529 13084
rect 13585 13082 13609 13084
rect 13665 13082 13689 13084
rect 13527 13030 13529 13082
rect 13591 13030 13603 13082
rect 13665 13030 13667 13082
rect 13505 13028 13529 13030
rect 13585 13028 13609 13030
rect 13665 13028 13689 13030
rect 13449 13008 13745 13028
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12481 13768 12582
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13449 11996 13745 12016
rect 13505 11994 13529 11996
rect 13585 11994 13609 11996
rect 13665 11994 13689 11996
rect 13527 11942 13529 11994
rect 13591 11942 13603 11994
rect 13665 11942 13667 11994
rect 13505 11940 13529 11942
rect 13585 11940 13609 11942
rect 13665 11940 13689 11942
rect 13449 11920 13745 11940
rect 13449 10908 13745 10928
rect 13505 10906 13529 10908
rect 13585 10906 13609 10908
rect 13665 10906 13689 10908
rect 13527 10854 13529 10906
rect 13591 10854 13603 10906
rect 13665 10854 13667 10906
rect 13505 10852 13529 10854
rect 13585 10852 13609 10854
rect 13665 10852 13689 10854
rect 13449 10832 13745 10852
rect 13832 10810 13860 15846
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13449 9820 13745 9840
rect 13505 9818 13529 9820
rect 13585 9818 13609 9820
rect 13665 9818 13689 9820
rect 13527 9766 13529 9818
rect 13591 9766 13603 9818
rect 13665 9766 13667 9818
rect 13505 9764 13529 9766
rect 13585 9764 13609 9766
rect 13665 9764 13689 9766
rect 13449 9744 13745 9764
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13372 8838 13400 8978
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 7449 13400 8774
rect 13449 8732 13745 8752
rect 13505 8730 13529 8732
rect 13585 8730 13609 8732
rect 13665 8730 13689 8732
rect 13527 8678 13529 8730
rect 13591 8678 13603 8730
rect 13665 8678 13667 8730
rect 13505 8676 13529 8678
rect 13585 8676 13609 8678
rect 13665 8676 13689 8678
rect 13449 8656 13745 8676
rect 13449 7644 13745 7664
rect 13505 7642 13529 7644
rect 13585 7642 13609 7644
rect 13665 7642 13689 7644
rect 13527 7590 13529 7642
rect 13591 7590 13603 7642
rect 13665 7590 13667 7642
rect 13505 7588 13529 7590
rect 13585 7588 13609 7590
rect 13665 7588 13689 7590
rect 13449 7568 13745 7588
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13449 6556 13745 6576
rect 13505 6554 13529 6556
rect 13585 6554 13609 6556
rect 13665 6554 13689 6556
rect 13527 6502 13529 6554
rect 13591 6502 13603 6554
rect 13665 6502 13667 6554
rect 13505 6500 13529 6502
rect 13585 6500 13609 6502
rect 13665 6500 13689 6502
rect 13449 6480 13745 6500
rect 14016 6118 14044 19200
rect 14476 15434 14504 19200
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14844 14482 14872 19200
rect 15304 15978 15332 19200
rect 15474 17504 15530 17513
rect 15474 17439 15530 17448
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 15488 13530 15516 17439
rect 15672 15910 15700 19200
rect 15660 15904 15712 15910
rect 16132 15858 16160 19200
rect 15660 15846 15712 15852
rect 15764 15830 16160 15858
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 10538 14504 13126
rect 15764 11914 15792 15830
rect 15304 11886 15792 11914
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13449 5468 13745 5488
rect 13505 5466 13529 5468
rect 13585 5466 13609 5468
rect 13665 5466 13689 5468
rect 13527 5414 13529 5466
rect 13591 5414 13603 5466
rect 13665 5414 13667 5466
rect 13505 5412 13529 5414
rect 13585 5412 13609 5414
rect 13665 5412 13689 5414
rect 13449 5392 13745 5412
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13188 5166 13216 5306
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13004 3454 13124 3482
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12636 800 12664 3062
rect 13096 800 13124 3454
rect 13280 1986 13308 4082
rect 13372 2854 13400 4966
rect 13449 4380 13745 4400
rect 13505 4378 13529 4380
rect 13585 4378 13609 4380
rect 13665 4378 13689 4380
rect 13527 4326 13529 4378
rect 13591 4326 13603 4378
rect 13665 4326 13667 4378
rect 13505 4324 13529 4326
rect 13585 4324 13609 4326
rect 13665 4324 13689 4326
rect 13449 4304 13745 4324
rect 13832 4146 13860 4966
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13449 3292 13745 3312
rect 13505 3290 13529 3292
rect 13585 3290 13609 3292
rect 13665 3290 13689 3292
rect 13527 3238 13529 3290
rect 13591 3238 13603 3290
rect 13665 3238 13667 3290
rect 13505 3236 13529 3238
rect 13585 3236 13609 3238
rect 13665 3236 13689 3238
rect 13449 3216 13745 3236
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13449 2204 13745 2224
rect 13505 2202 13529 2204
rect 13585 2202 13609 2204
rect 13665 2202 13689 2204
rect 13527 2150 13529 2202
rect 13591 2150 13603 2202
rect 13665 2150 13667 2202
rect 13505 2148 13529 2150
rect 13585 2148 13609 2150
rect 13665 2148 13689 2150
rect 13449 2128 13745 2148
rect 13280 1958 13492 1986
rect 13464 800 13492 1958
rect 13924 800 13952 4558
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14384 800 14412 4014
rect 14476 2553 14504 10474
rect 15304 5710 15332 11886
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 5914 15424 11630
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15580 5370 15608 11698
rect 16500 11694 16528 19200
rect 16960 11762 16988 19200
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14462 2544 14518 2553
rect 14462 2479 14518 2488
rect 14752 800 14780 3946
rect 15212 800 15240 5238
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15672 800 15700 4694
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16040 800 16068 3130
rect 16500 800 16528 5170
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16960 800 16988 4082
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< via2 >>
rect 1490 8336 1546 8392
rect 3454 17434 3510 17436
rect 3534 17434 3590 17436
rect 3614 17434 3670 17436
rect 3694 17434 3750 17436
rect 3454 17382 3480 17434
rect 3480 17382 3510 17434
rect 3534 17382 3544 17434
rect 3544 17382 3590 17434
rect 3614 17382 3660 17434
rect 3660 17382 3670 17434
rect 3694 17382 3724 17434
rect 3724 17382 3750 17434
rect 3454 17380 3510 17382
rect 3534 17380 3590 17382
rect 3614 17380 3670 17382
rect 3694 17380 3750 17382
rect 3454 16346 3510 16348
rect 3534 16346 3590 16348
rect 3614 16346 3670 16348
rect 3694 16346 3750 16348
rect 3454 16294 3480 16346
rect 3480 16294 3510 16346
rect 3534 16294 3544 16346
rect 3544 16294 3590 16346
rect 3614 16294 3660 16346
rect 3660 16294 3670 16346
rect 3694 16294 3724 16346
rect 3724 16294 3750 16346
rect 3454 16292 3510 16294
rect 3534 16292 3590 16294
rect 3614 16292 3670 16294
rect 3694 16292 3750 16294
rect 2778 15000 2834 15056
rect 3454 15258 3510 15260
rect 3534 15258 3590 15260
rect 3614 15258 3670 15260
rect 3694 15258 3750 15260
rect 3454 15206 3480 15258
rect 3480 15206 3510 15258
rect 3534 15206 3544 15258
rect 3544 15206 3590 15258
rect 3614 15206 3660 15258
rect 3660 15206 3670 15258
rect 3694 15206 3724 15258
rect 3724 15206 3750 15258
rect 3454 15204 3510 15206
rect 3534 15204 3590 15206
rect 3614 15204 3670 15206
rect 3694 15204 3750 15206
rect 3454 14170 3510 14172
rect 3534 14170 3590 14172
rect 3614 14170 3670 14172
rect 3694 14170 3750 14172
rect 3454 14118 3480 14170
rect 3480 14118 3510 14170
rect 3534 14118 3544 14170
rect 3544 14118 3590 14170
rect 3614 14118 3660 14170
rect 3660 14118 3670 14170
rect 3694 14118 3724 14170
rect 3724 14118 3750 14170
rect 3454 14116 3510 14118
rect 3534 14116 3590 14118
rect 3614 14116 3670 14118
rect 3694 14116 3750 14118
rect 3454 13082 3510 13084
rect 3534 13082 3590 13084
rect 3614 13082 3670 13084
rect 3694 13082 3750 13084
rect 3454 13030 3480 13082
rect 3480 13030 3510 13082
rect 3534 13030 3544 13082
rect 3544 13030 3590 13082
rect 3614 13030 3660 13082
rect 3660 13030 3670 13082
rect 3694 13030 3724 13082
rect 3724 13030 3750 13082
rect 3454 13028 3510 13030
rect 3534 13028 3590 13030
rect 3614 13028 3670 13030
rect 3694 13028 3750 13030
rect 3454 11994 3510 11996
rect 3534 11994 3590 11996
rect 3614 11994 3670 11996
rect 3694 11994 3750 11996
rect 3454 11942 3480 11994
rect 3480 11942 3510 11994
rect 3534 11942 3544 11994
rect 3544 11942 3590 11994
rect 3614 11942 3660 11994
rect 3660 11942 3670 11994
rect 3694 11942 3724 11994
rect 3724 11942 3750 11994
rect 3454 11940 3510 11942
rect 3534 11940 3590 11942
rect 3614 11940 3670 11942
rect 3694 11940 3750 11942
rect 3330 11600 3386 11656
rect 3454 10906 3510 10908
rect 3534 10906 3590 10908
rect 3614 10906 3670 10908
rect 3694 10906 3750 10908
rect 3454 10854 3480 10906
rect 3480 10854 3510 10906
rect 3534 10854 3544 10906
rect 3544 10854 3590 10906
rect 3614 10854 3660 10906
rect 3660 10854 3670 10906
rect 3694 10854 3724 10906
rect 3724 10854 3750 10906
rect 3454 10852 3510 10854
rect 3534 10852 3590 10854
rect 3614 10852 3670 10854
rect 3694 10852 3750 10854
rect 3454 9818 3510 9820
rect 3534 9818 3590 9820
rect 3614 9818 3670 9820
rect 3694 9818 3750 9820
rect 3454 9766 3480 9818
rect 3480 9766 3510 9818
rect 3534 9766 3544 9818
rect 3544 9766 3590 9818
rect 3614 9766 3660 9818
rect 3660 9766 3670 9818
rect 3694 9766 3724 9818
rect 3724 9766 3750 9818
rect 3454 9764 3510 9766
rect 3534 9764 3590 9766
rect 3614 9764 3670 9766
rect 3694 9764 3750 9766
rect 3454 8730 3510 8732
rect 3534 8730 3590 8732
rect 3614 8730 3670 8732
rect 3694 8730 3750 8732
rect 3454 8678 3480 8730
rect 3480 8678 3510 8730
rect 3534 8678 3544 8730
rect 3544 8678 3590 8730
rect 3614 8678 3660 8730
rect 3660 8678 3670 8730
rect 3694 8678 3724 8730
rect 3724 8678 3750 8730
rect 3454 8676 3510 8678
rect 3534 8676 3590 8678
rect 3614 8676 3670 8678
rect 3694 8676 3750 8678
rect 3454 7642 3510 7644
rect 3534 7642 3590 7644
rect 3614 7642 3670 7644
rect 3694 7642 3750 7644
rect 3454 7590 3480 7642
rect 3480 7590 3510 7642
rect 3534 7590 3544 7642
rect 3544 7590 3590 7642
rect 3614 7590 3660 7642
rect 3660 7590 3670 7642
rect 3694 7590 3724 7642
rect 3724 7590 3750 7642
rect 3454 7588 3510 7590
rect 3534 7588 3590 7590
rect 3614 7588 3670 7590
rect 3694 7588 3750 7590
rect 3454 6554 3510 6556
rect 3534 6554 3590 6556
rect 3614 6554 3670 6556
rect 3694 6554 3750 6556
rect 3454 6502 3480 6554
rect 3480 6502 3510 6554
rect 3534 6502 3544 6554
rect 3544 6502 3590 6554
rect 3614 6502 3660 6554
rect 3660 6502 3670 6554
rect 3694 6502 3724 6554
rect 3724 6502 3750 6554
rect 3454 6500 3510 6502
rect 3534 6500 3590 6502
rect 3614 6500 3670 6502
rect 3694 6500 3750 6502
rect 3454 5466 3510 5468
rect 3534 5466 3590 5468
rect 3614 5466 3670 5468
rect 3694 5466 3750 5468
rect 3454 5414 3480 5466
rect 3480 5414 3510 5466
rect 3534 5414 3544 5466
rect 3544 5414 3590 5466
rect 3614 5414 3660 5466
rect 3660 5414 3670 5466
rect 3694 5414 3724 5466
rect 3724 5414 3750 5466
rect 3454 5412 3510 5414
rect 3534 5412 3590 5414
rect 3614 5412 3670 5414
rect 3694 5412 3750 5414
rect 2962 4936 3018 4992
rect 4066 18264 4122 18320
rect 3454 4378 3510 4380
rect 3534 4378 3590 4380
rect 3614 4378 3670 4380
rect 3694 4378 3750 4380
rect 3454 4326 3480 4378
rect 3480 4326 3510 4378
rect 3534 4326 3544 4378
rect 3544 4326 3590 4378
rect 3614 4326 3660 4378
rect 3660 4326 3670 4378
rect 3694 4326 3724 4378
rect 3724 4326 3750 4378
rect 3454 4324 3510 4326
rect 3534 4324 3590 4326
rect 3614 4324 3670 4326
rect 3694 4324 3750 4326
rect 1582 1672 1638 1728
rect 3454 3290 3510 3292
rect 3534 3290 3590 3292
rect 3614 3290 3670 3292
rect 3694 3290 3750 3292
rect 3454 3238 3480 3290
rect 3480 3238 3510 3290
rect 3534 3238 3544 3290
rect 3544 3238 3590 3290
rect 3614 3238 3660 3290
rect 3660 3238 3670 3290
rect 3694 3238 3724 3290
rect 3724 3238 3750 3290
rect 3454 3236 3510 3238
rect 3534 3236 3590 3238
rect 3614 3236 3670 3238
rect 3694 3236 3750 3238
rect 3454 2202 3510 2204
rect 3534 2202 3590 2204
rect 3614 2202 3670 2204
rect 3694 2202 3750 2204
rect 3454 2150 3480 2202
rect 3480 2150 3510 2202
rect 3534 2150 3544 2202
rect 3544 2150 3590 2202
rect 3614 2150 3660 2202
rect 3660 2150 3670 2202
rect 3694 2150 3724 2202
rect 3724 2150 3750 2202
rect 3454 2148 3510 2150
rect 3534 2148 3590 2150
rect 3614 2148 3670 2150
rect 3694 2148 3750 2150
rect 5953 16890 6009 16892
rect 6033 16890 6089 16892
rect 6113 16890 6169 16892
rect 6193 16890 6249 16892
rect 5953 16838 5979 16890
rect 5979 16838 6009 16890
rect 6033 16838 6043 16890
rect 6043 16838 6089 16890
rect 6113 16838 6159 16890
rect 6159 16838 6169 16890
rect 6193 16838 6223 16890
rect 6223 16838 6249 16890
rect 5953 16836 6009 16838
rect 6033 16836 6089 16838
rect 6113 16836 6169 16838
rect 6193 16836 6249 16838
rect 5953 15802 6009 15804
rect 6033 15802 6089 15804
rect 6113 15802 6169 15804
rect 6193 15802 6249 15804
rect 5953 15750 5979 15802
rect 5979 15750 6009 15802
rect 6033 15750 6043 15802
rect 6043 15750 6089 15802
rect 6113 15750 6159 15802
rect 6159 15750 6169 15802
rect 6193 15750 6223 15802
rect 6223 15750 6249 15802
rect 5953 15748 6009 15750
rect 6033 15748 6089 15750
rect 6113 15748 6169 15750
rect 6193 15748 6249 15750
rect 5953 14714 6009 14716
rect 6033 14714 6089 14716
rect 6113 14714 6169 14716
rect 6193 14714 6249 14716
rect 5953 14662 5979 14714
rect 5979 14662 6009 14714
rect 6033 14662 6043 14714
rect 6043 14662 6089 14714
rect 6113 14662 6159 14714
rect 6159 14662 6169 14714
rect 6193 14662 6223 14714
rect 6223 14662 6249 14714
rect 5953 14660 6009 14662
rect 6033 14660 6089 14662
rect 6113 14660 6169 14662
rect 6193 14660 6249 14662
rect 5953 13626 6009 13628
rect 6033 13626 6089 13628
rect 6113 13626 6169 13628
rect 6193 13626 6249 13628
rect 5953 13574 5979 13626
rect 5979 13574 6009 13626
rect 6033 13574 6043 13626
rect 6043 13574 6089 13626
rect 6113 13574 6159 13626
rect 6159 13574 6169 13626
rect 6193 13574 6223 13626
rect 6223 13574 6249 13626
rect 5953 13572 6009 13574
rect 6033 13572 6089 13574
rect 6113 13572 6169 13574
rect 6193 13572 6249 13574
rect 5953 12538 6009 12540
rect 6033 12538 6089 12540
rect 6113 12538 6169 12540
rect 6193 12538 6249 12540
rect 5953 12486 5979 12538
rect 5979 12486 6009 12538
rect 6033 12486 6043 12538
rect 6043 12486 6089 12538
rect 6113 12486 6159 12538
rect 6159 12486 6169 12538
rect 6193 12486 6223 12538
rect 6223 12486 6249 12538
rect 5953 12484 6009 12486
rect 6033 12484 6089 12486
rect 6113 12484 6169 12486
rect 6193 12484 6249 12486
rect 5953 11450 6009 11452
rect 6033 11450 6089 11452
rect 6113 11450 6169 11452
rect 6193 11450 6249 11452
rect 5953 11398 5979 11450
rect 5979 11398 6009 11450
rect 6033 11398 6043 11450
rect 6043 11398 6089 11450
rect 6113 11398 6159 11450
rect 6159 11398 6169 11450
rect 6193 11398 6223 11450
rect 6223 11398 6249 11450
rect 5953 11396 6009 11398
rect 6033 11396 6089 11398
rect 6113 11396 6169 11398
rect 6193 11396 6249 11398
rect 5953 10362 6009 10364
rect 6033 10362 6089 10364
rect 6113 10362 6169 10364
rect 6193 10362 6249 10364
rect 5953 10310 5979 10362
rect 5979 10310 6009 10362
rect 6033 10310 6043 10362
rect 6043 10310 6089 10362
rect 6113 10310 6159 10362
rect 6159 10310 6169 10362
rect 6193 10310 6223 10362
rect 6223 10310 6249 10362
rect 5953 10308 6009 10310
rect 6033 10308 6089 10310
rect 6113 10308 6169 10310
rect 6193 10308 6249 10310
rect 5953 9274 6009 9276
rect 6033 9274 6089 9276
rect 6113 9274 6169 9276
rect 6193 9274 6249 9276
rect 5953 9222 5979 9274
rect 5979 9222 6009 9274
rect 6033 9222 6043 9274
rect 6043 9222 6089 9274
rect 6113 9222 6159 9274
rect 6159 9222 6169 9274
rect 6193 9222 6223 9274
rect 6223 9222 6249 9274
rect 5953 9220 6009 9222
rect 6033 9220 6089 9222
rect 6113 9220 6169 9222
rect 6193 9220 6249 9222
rect 5953 8186 6009 8188
rect 6033 8186 6089 8188
rect 6113 8186 6169 8188
rect 6193 8186 6249 8188
rect 5953 8134 5979 8186
rect 5979 8134 6009 8186
rect 6033 8134 6043 8186
rect 6043 8134 6089 8186
rect 6113 8134 6159 8186
rect 6159 8134 6169 8186
rect 6193 8134 6223 8186
rect 6223 8134 6249 8186
rect 5953 8132 6009 8134
rect 6033 8132 6089 8134
rect 6113 8132 6169 8134
rect 6193 8132 6249 8134
rect 5953 7098 6009 7100
rect 6033 7098 6089 7100
rect 6113 7098 6169 7100
rect 6193 7098 6249 7100
rect 5953 7046 5979 7098
rect 5979 7046 6009 7098
rect 6033 7046 6043 7098
rect 6043 7046 6089 7098
rect 6113 7046 6159 7098
rect 6159 7046 6169 7098
rect 6193 7046 6223 7098
rect 6223 7046 6249 7098
rect 5953 7044 6009 7046
rect 6033 7044 6089 7046
rect 6113 7044 6169 7046
rect 6193 7044 6249 7046
rect 5953 6010 6009 6012
rect 6033 6010 6089 6012
rect 6113 6010 6169 6012
rect 6193 6010 6249 6012
rect 5953 5958 5979 6010
rect 5979 5958 6009 6010
rect 6033 5958 6043 6010
rect 6043 5958 6089 6010
rect 6113 5958 6159 6010
rect 6159 5958 6169 6010
rect 6193 5958 6223 6010
rect 6223 5958 6249 6010
rect 5953 5956 6009 5958
rect 6033 5956 6089 5958
rect 6113 5956 6169 5958
rect 6193 5956 6249 5958
rect 6826 5208 6882 5264
rect 5953 4922 6009 4924
rect 6033 4922 6089 4924
rect 6113 4922 6169 4924
rect 6193 4922 6249 4924
rect 5953 4870 5979 4922
rect 5979 4870 6009 4922
rect 6033 4870 6043 4922
rect 6043 4870 6089 4922
rect 6113 4870 6159 4922
rect 6159 4870 6169 4922
rect 6193 4870 6223 4922
rect 6223 4870 6249 4922
rect 5953 4868 6009 4870
rect 6033 4868 6089 4870
rect 6113 4868 6169 4870
rect 6193 4868 6249 4870
rect 5953 3834 6009 3836
rect 6033 3834 6089 3836
rect 6113 3834 6169 3836
rect 6193 3834 6249 3836
rect 5953 3782 5979 3834
rect 5979 3782 6009 3834
rect 6033 3782 6043 3834
rect 6043 3782 6089 3834
rect 6113 3782 6159 3834
rect 6159 3782 6169 3834
rect 6193 3782 6223 3834
rect 6223 3782 6249 3834
rect 5953 3780 6009 3782
rect 6033 3780 6089 3782
rect 6113 3780 6169 3782
rect 6193 3780 6249 3782
rect 5354 856 5410 912
rect 5953 2746 6009 2748
rect 6033 2746 6089 2748
rect 6113 2746 6169 2748
rect 6193 2746 6249 2748
rect 5953 2694 5979 2746
rect 5979 2694 6009 2746
rect 6033 2694 6043 2746
rect 6043 2694 6089 2746
rect 6113 2694 6159 2746
rect 6159 2694 6169 2746
rect 6193 2694 6223 2746
rect 6223 2694 6249 2746
rect 5953 2692 6009 2694
rect 6033 2692 6089 2694
rect 6113 2692 6169 2694
rect 6193 2692 6249 2694
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8478 17434
rect 8478 17382 8508 17434
rect 8532 17382 8542 17434
rect 8542 17382 8588 17434
rect 8612 17382 8658 17434
rect 8658 17382 8668 17434
rect 8692 17382 8722 17434
rect 8722 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8478 16346
rect 8478 16294 8508 16346
rect 8532 16294 8542 16346
rect 8542 16294 8588 16346
rect 8612 16294 8658 16346
rect 8658 16294 8668 16346
rect 8692 16294 8722 16346
rect 8722 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8478 15258
rect 8478 15206 8508 15258
rect 8532 15206 8542 15258
rect 8542 15206 8588 15258
rect 8612 15206 8658 15258
rect 8658 15206 8668 15258
rect 8692 15206 8722 15258
rect 8722 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8478 14170
rect 8478 14118 8508 14170
rect 8532 14118 8542 14170
rect 8542 14118 8588 14170
rect 8612 14118 8658 14170
rect 8658 14118 8668 14170
rect 8692 14118 8722 14170
rect 8722 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8478 13082
rect 8478 13030 8508 13082
rect 8532 13030 8542 13082
rect 8542 13030 8588 13082
rect 8612 13030 8658 13082
rect 8658 13030 8668 13082
rect 8692 13030 8722 13082
rect 8722 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8478 11994
rect 8478 11942 8508 11994
rect 8532 11942 8542 11994
rect 8542 11942 8588 11994
rect 8612 11942 8658 11994
rect 8658 11942 8668 11994
rect 8692 11942 8722 11994
rect 8722 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8478 10906
rect 8478 10854 8508 10906
rect 8532 10854 8542 10906
rect 8542 10854 8588 10906
rect 8612 10854 8658 10906
rect 8658 10854 8668 10906
rect 8692 10854 8722 10906
rect 8722 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8478 9818
rect 8478 9766 8508 9818
rect 8532 9766 8542 9818
rect 8542 9766 8588 9818
rect 8612 9766 8658 9818
rect 8658 9766 8668 9818
rect 8692 9766 8722 9818
rect 8722 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 10230 19080 10286 19136
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8478 8730
rect 8478 8678 8508 8730
rect 8532 8678 8542 8730
rect 8542 8678 8588 8730
rect 8612 8678 8658 8730
rect 8658 8678 8668 8730
rect 8692 8678 8722 8730
rect 8722 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8478 7642
rect 8478 7590 8508 7642
rect 8532 7590 8542 7642
rect 8542 7590 8588 7642
rect 8612 7590 8658 7642
rect 8658 7590 8668 7642
rect 8692 7590 8722 7642
rect 8722 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8478 6554
rect 8478 6502 8508 6554
rect 8532 6502 8542 6554
rect 8542 6502 8588 6554
rect 8612 6502 8658 6554
rect 8658 6502 8668 6554
rect 8692 6502 8722 6554
rect 8722 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8478 5466
rect 8478 5414 8508 5466
rect 8532 5414 8542 5466
rect 8542 5414 8588 5466
rect 8612 5414 8658 5466
rect 8658 5414 8668 5466
rect 8692 5414 8722 5466
rect 8722 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8206 5072 8262 5128
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8478 4378
rect 8478 4326 8508 4378
rect 8532 4326 8542 4378
rect 8542 4326 8588 4378
rect 8612 4326 8658 4378
rect 8658 4326 8668 4378
rect 8692 4326 8722 4378
rect 8722 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8478 3290
rect 8478 3238 8508 3290
rect 8532 3238 8542 3290
rect 8542 3238 8588 3290
rect 8612 3238 8658 3290
rect 8658 3238 8668 3290
rect 8692 3238 8722 3290
rect 8722 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8478 2202
rect 8478 2150 8508 2202
rect 8532 2150 8542 2202
rect 8542 2150 8588 2202
rect 8612 2150 8658 2202
rect 8658 2150 8668 2202
rect 8692 2150 8722 2202
rect 8722 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9494 9560 9550 9616
rect 9586 9424 9642 9480
rect 9586 9288 9642 9344
rect 9402 5344 9458 5400
rect 9126 856 9182 912
rect 10950 16890 11006 16892
rect 11030 16890 11086 16892
rect 11110 16890 11166 16892
rect 11190 16890 11246 16892
rect 10950 16838 10976 16890
rect 10976 16838 11006 16890
rect 11030 16838 11040 16890
rect 11040 16838 11086 16890
rect 11110 16838 11156 16890
rect 11156 16838 11166 16890
rect 11190 16838 11220 16890
rect 11220 16838 11246 16890
rect 10950 16836 11006 16838
rect 11030 16836 11086 16838
rect 11110 16836 11166 16838
rect 11190 16836 11246 16838
rect 10950 15802 11006 15804
rect 11030 15802 11086 15804
rect 11110 15802 11166 15804
rect 11190 15802 11246 15804
rect 10950 15750 10976 15802
rect 10976 15750 11006 15802
rect 11030 15750 11040 15802
rect 11040 15750 11086 15802
rect 11110 15750 11156 15802
rect 11156 15750 11166 15802
rect 11190 15750 11220 15802
rect 11220 15750 11246 15802
rect 10950 15748 11006 15750
rect 11030 15748 11086 15750
rect 11110 15748 11166 15750
rect 11190 15748 11246 15750
rect 10230 9560 10286 9616
rect 9586 856 9642 912
rect 10506 9968 10562 10024
rect 10950 14714 11006 14716
rect 11030 14714 11086 14716
rect 11110 14714 11166 14716
rect 11190 14714 11246 14716
rect 10950 14662 10976 14714
rect 10976 14662 11006 14714
rect 11030 14662 11040 14714
rect 11040 14662 11086 14714
rect 11110 14662 11156 14714
rect 11156 14662 11166 14714
rect 11190 14662 11220 14714
rect 11220 14662 11246 14714
rect 10950 14660 11006 14662
rect 11030 14660 11086 14662
rect 11110 14660 11166 14662
rect 11190 14660 11246 14662
rect 10950 13626 11006 13628
rect 11030 13626 11086 13628
rect 11110 13626 11166 13628
rect 11190 13626 11246 13628
rect 10950 13574 10976 13626
rect 10976 13574 11006 13626
rect 11030 13574 11040 13626
rect 11040 13574 11086 13626
rect 11110 13574 11156 13626
rect 11156 13574 11166 13626
rect 11190 13574 11220 13626
rect 11220 13574 11246 13626
rect 10950 13572 11006 13574
rect 11030 13572 11086 13574
rect 11110 13572 11166 13574
rect 11190 13572 11246 13574
rect 10950 12538 11006 12540
rect 11030 12538 11086 12540
rect 11110 12538 11166 12540
rect 11190 12538 11246 12540
rect 10950 12486 10976 12538
rect 10976 12486 11006 12538
rect 11030 12486 11040 12538
rect 11040 12486 11086 12538
rect 11110 12486 11156 12538
rect 11156 12486 11166 12538
rect 11190 12486 11220 12538
rect 11220 12486 11246 12538
rect 10950 12484 11006 12486
rect 11030 12484 11086 12486
rect 11110 12484 11166 12486
rect 11190 12484 11246 12486
rect 10950 11450 11006 11452
rect 11030 11450 11086 11452
rect 11110 11450 11166 11452
rect 11190 11450 11246 11452
rect 10950 11398 10976 11450
rect 10976 11398 11006 11450
rect 11030 11398 11040 11450
rect 11040 11398 11086 11450
rect 11110 11398 11156 11450
rect 11156 11398 11166 11450
rect 11190 11398 11220 11450
rect 11220 11398 11246 11450
rect 10950 11396 11006 11398
rect 11030 11396 11086 11398
rect 11110 11396 11166 11398
rect 11190 11396 11246 11398
rect 10950 10362 11006 10364
rect 11030 10362 11086 10364
rect 11110 10362 11166 10364
rect 11190 10362 11246 10364
rect 10950 10310 10976 10362
rect 10976 10310 11006 10362
rect 11030 10310 11040 10362
rect 11040 10310 11086 10362
rect 11110 10310 11156 10362
rect 11156 10310 11166 10362
rect 11190 10310 11220 10362
rect 11220 10310 11246 10362
rect 10950 10308 11006 10310
rect 11030 10308 11086 10310
rect 11110 10308 11166 10310
rect 11190 10308 11246 10310
rect 10950 9274 11006 9276
rect 11030 9274 11086 9276
rect 11110 9274 11166 9276
rect 11190 9274 11246 9276
rect 10950 9222 10976 9274
rect 10976 9222 11006 9274
rect 11030 9222 11040 9274
rect 11040 9222 11086 9274
rect 11110 9222 11156 9274
rect 11156 9222 11166 9274
rect 11190 9222 11220 9274
rect 11220 9222 11246 9274
rect 10950 9220 11006 9222
rect 11030 9220 11086 9222
rect 11110 9220 11166 9222
rect 11190 9220 11246 9222
rect 10950 8186 11006 8188
rect 11030 8186 11086 8188
rect 11110 8186 11166 8188
rect 11190 8186 11246 8188
rect 10950 8134 10976 8186
rect 10976 8134 11006 8186
rect 11030 8134 11040 8186
rect 11040 8134 11086 8186
rect 11110 8134 11156 8186
rect 11156 8134 11166 8186
rect 11190 8134 11220 8186
rect 11220 8134 11246 8186
rect 10950 8132 11006 8134
rect 11030 8132 11086 8134
rect 11110 8132 11166 8134
rect 11190 8132 11246 8134
rect 10950 7098 11006 7100
rect 11030 7098 11086 7100
rect 11110 7098 11166 7100
rect 11190 7098 11246 7100
rect 10950 7046 10976 7098
rect 10976 7046 11006 7098
rect 11030 7046 11040 7098
rect 11040 7046 11086 7098
rect 11110 7046 11156 7098
rect 11156 7046 11166 7098
rect 11190 7046 11220 7098
rect 11220 7046 11246 7098
rect 10950 7044 11006 7046
rect 11030 7044 11086 7046
rect 11110 7044 11166 7046
rect 11190 7044 11246 7046
rect 10950 6010 11006 6012
rect 11030 6010 11086 6012
rect 11110 6010 11166 6012
rect 11190 6010 11246 6012
rect 10950 5958 10976 6010
rect 10976 5958 11006 6010
rect 11030 5958 11040 6010
rect 11040 5958 11086 6010
rect 11110 5958 11156 6010
rect 11156 5958 11166 6010
rect 11190 5958 11220 6010
rect 11220 5958 11246 6010
rect 10950 5956 11006 5958
rect 11030 5956 11086 5958
rect 11110 5956 11166 5958
rect 11190 5956 11246 5958
rect 12898 5364 12954 5400
rect 12898 5344 12900 5364
rect 12900 5344 12952 5364
rect 12952 5344 12954 5364
rect 11058 5208 11114 5264
rect 10950 4922 11006 4924
rect 11030 4922 11086 4924
rect 11110 4922 11166 4924
rect 11190 4922 11246 4924
rect 10950 4870 10976 4922
rect 10976 4870 11006 4922
rect 11030 4870 11040 4922
rect 11040 4870 11086 4922
rect 11110 4870 11156 4922
rect 11156 4870 11166 4922
rect 11190 4870 11220 4922
rect 11220 4870 11246 4922
rect 10950 4868 11006 4870
rect 11030 4868 11086 4870
rect 11110 4868 11166 4870
rect 11190 4868 11246 4870
rect 12622 5072 12678 5128
rect 10950 3834 11006 3836
rect 11030 3834 11086 3836
rect 11110 3834 11166 3836
rect 11190 3834 11246 3836
rect 10950 3782 10976 3834
rect 10976 3782 11006 3834
rect 11030 3782 11040 3834
rect 11040 3782 11086 3834
rect 11110 3782 11156 3834
rect 11156 3782 11166 3834
rect 11190 3782 11220 3834
rect 11220 3782 11246 3834
rect 10950 3780 11006 3782
rect 11030 3780 11086 3782
rect 11110 3780 11166 3782
rect 11190 3780 11246 3782
rect 10506 856 10562 912
rect 10950 2746 11006 2748
rect 11030 2746 11086 2748
rect 11110 2746 11166 2748
rect 11190 2746 11246 2748
rect 10950 2694 10976 2746
rect 10976 2694 11006 2746
rect 11030 2694 11040 2746
rect 11040 2694 11086 2746
rect 11110 2694 11156 2746
rect 11156 2694 11166 2746
rect 11190 2694 11220 2746
rect 11220 2694 11246 2746
rect 10950 2692 11006 2694
rect 11030 2692 11086 2694
rect 11110 2692 11166 2694
rect 11190 2692 11246 2694
rect 13449 17434 13505 17436
rect 13529 17434 13585 17436
rect 13609 17434 13665 17436
rect 13689 17434 13745 17436
rect 13449 17382 13475 17434
rect 13475 17382 13505 17434
rect 13529 17382 13539 17434
rect 13539 17382 13585 17434
rect 13609 17382 13655 17434
rect 13655 17382 13665 17434
rect 13689 17382 13719 17434
rect 13719 17382 13745 17434
rect 13449 17380 13505 17382
rect 13529 17380 13585 17382
rect 13609 17380 13665 17382
rect 13689 17380 13745 17382
rect 13449 16346 13505 16348
rect 13529 16346 13585 16348
rect 13609 16346 13665 16348
rect 13689 16346 13745 16348
rect 13449 16294 13475 16346
rect 13475 16294 13505 16346
rect 13529 16294 13539 16346
rect 13539 16294 13585 16346
rect 13609 16294 13655 16346
rect 13655 16294 13665 16346
rect 13689 16294 13719 16346
rect 13719 16294 13745 16346
rect 13449 16292 13505 16294
rect 13529 16292 13585 16294
rect 13609 16292 13665 16294
rect 13689 16292 13745 16294
rect 13449 15258 13505 15260
rect 13529 15258 13585 15260
rect 13609 15258 13665 15260
rect 13689 15258 13745 15260
rect 13449 15206 13475 15258
rect 13475 15206 13505 15258
rect 13529 15206 13539 15258
rect 13539 15206 13585 15258
rect 13609 15206 13655 15258
rect 13655 15206 13665 15258
rect 13689 15206 13719 15258
rect 13719 15206 13745 15258
rect 13449 15204 13505 15206
rect 13529 15204 13585 15206
rect 13609 15204 13665 15206
rect 13689 15204 13745 15206
rect 13449 14170 13505 14172
rect 13529 14170 13585 14172
rect 13609 14170 13665 14172
rect 13689 14170 13745 14172
rect 13449 14118 13475 14170
rect 13475 14118 13505 14170
rect 13529 14118 13539 14170
rect 13539 14118 13585 14170
rect 13609 14118 13655 14170
rect 13655 14118 13665 14170
rect 13689 14118 13719 14170
rect 13719 14118 13745 14170
rect 13449 14116 13505 14118
rect 13529 14116 13585 14118
rect 13609 14116 13665 14118
rect 13689 14116 13745 14118
rect 13449 13082 13505 13084
rect 13529 13082 13585 13084
rect 13609 13082 13665 13084
rect 13689 13082 13745 13084
rect 13449 13030 13475 13082
rect 13475 13030 13505 13082
rect 13529 13030 13539 13082
rect 13539 13030 13585 13082
rect 13609 13030 13655 13082
rect 13655 13030 13665 13082
rect 13689 13030 13719 13082
rect 13719 13030 13745 13082
rect 13449 13028 13505 13030
rect 13529 13028 13585 13030
rect 13609 13028 13665 13030
rect 13689 13028 13745 13030
rect 13726 12416 13782 12472
rect 13449 11994 13505 11996
rect 13529 11994 13585 11996
rect 13609 11994 13665 11996
rect 13689 11994 13745 11996
rect 13449 11942 13475 11994
rect 13475 11942 13505 11994
rect 13529 11942 13539 11994
rect 13539 11942 13585 11994
rect 13609 11942 13655 11994
rect 13655 11942 13665 11994
rect 13689 11942 13719 11994
rect 13719 11942 13745 11994
rect 13449 11940 13505 11942
rect 13529 11940 13585 11942
rect 13609 11940 13665 11942
rect 13689 11940 13745 11942
rect 13449 10906 13505 10908
rect 13529 10906 13585 10908
rect 13609 10906 13665 10908
rect 13689 10906 13745 10908
rect 13449 10854 13475 10906
rect 13475 10854 13505 10906
rect 13529 10854 13539 10906
rect 13539 10854 13585 10906
rect 13609 10854 13655 10906
rect 13655 10854 13665 10906
rect 13689 10854 13719 10906
rect 13719 10854 13745 10906
rect 13449 10852 13505 10854
rect 13529 10852 13585 10854
rect 13609 10852 13665 10854
rect 13689 10852 13745 10854
rect 13449 9818 13505 9820
rect 13529 9818 13585 9820
rect 13609 9818 13665 9820
rect 13689 9818 13745 9820
rect 13449 9766 13475 9818
rect 13475 9766 13505 9818
rect 13529 9766 13539 9818
rect 13539 9766 13585 9818
rect 13609 9766 13655 9818
rect 13655 9766 13665 9818
rect 13689 9766 13719 9818
rect 13719 9766 13745 9818
rect 13449 9764 13505 9766
rect 13529 9764 13585 9766
rect 13609 9764 13665 9766
rect 13689 9764 13745 9766
rect 13449 8730 13505 8732
rect 13529 8730 13585 8732
rect 13609 8730 13665 8732
rect 13689 8730 13745 8732
rect 13449 8678 13475 8730
rect 13475 8678 13505 8730
rect 13529 8678 13539 8730
rect 13539 8678 13585 8730
rect 13609 8678 13655 8730
rect 13655 8678 13665 8730
rect 13689 8678 13719 8730
rect 13719 8678 13745 8730
rect 13449 8676 13505 8678
rect 13529 8676 13585 8678
rect 13609 8676 13665 8678
rect 13689 8676 13745 8678
rect 13449 7642 13505 7644
rect 13529 7642 13585 7644
rect 13609 7642 13665 7644
rect 13689 7642 13745 7644
rect 13449 7590 13475 7642
rect 13475 7590 13505 7642
rect 13529 7590 13539 7642
rect 13539 7590 13585 7642
rect 13609 7590 13655 7642
rect 13655 7590 13665 7642
rect 13689 7590 13719 7642
rect 13719 7590 13745 7642
rect 13449 7588 13505 7590
rect 13529 7588 13585 7590
rect 13609 7588 13665 7590
rect 13689 7588 13745 7590
rect 13358 7384 13414 7440
rect 13449 6554 13505 6556
rect 13529 6554 13585 6556
rect 13609 6554 13665 6556
rect 13689 6554 13745 6556
rect 13449 6502 13475 6554
rect 13475 6502 13505 6554
rect 13529 6502 13539 6554
rect 13539 6502 13585 6554
rect 13609 6502 13655 6554
rect 13655 6502 13665 6554
rect 13689 6502 13719 6554
rect 13719 6502 13745 6554
rect 13449 6500 13505 6502
rect 13529 6500 13585 6502
rect 13609 6500 13665 6502
rect 13689 6500 13745 6502
rect 15474 17448 15530 17504
rect 13449 5466 13505 5468
rect 13529 5466 13585 5468
rect 13609 5466 13665 5468
rect 13689 5466 13745 5468
rect 13449 5414 13475 5466
rect 13475 5414 13505 5466
rect 13529 5414 13539 5466
rect 13539 5414 13585 5466
rect 13609 5414 13655 5466
rect 13655 5414 13665 5466
rect 13689 5414 13719 5466
rect 13719 5414 13745 5466
rect 13449 5412 13505 5414
rect 13529 5412 13585 5414
rect 13609 5412 13665 5414
rect 13689 5412 13745 5414
rect 13449 4378 13505 4380
rect 13529 4378 13585 4380
rect 13609 4378 13665 4380
rect 13689 4378 13745 4380
rect 13449 4326 13475 4378
rect 13475 4326 13505 4378
rect 13529 4326 13539 4378
rect 13539 4326 13585 4378
rect 13609 4326 13655 4378
rect 13655 4326 13665 4378
rect 13689 4326 13719 4378
rect 13719 4326 13745 4378
rect 13449 4324 13505 4326
rect 13529 4324 13585 4326
rect 13609 4324 13665 4326
rect 13689 4324 13745 4326
rect 13449 3290 13505 3292
rect 13529 3290 13585 3292
rect 13609 3290 13665 3292
rect 13689 3290 13745 3292
rect 13449 3238 13475 3290
rect 13475 3238 13505 3290
rect 13529 3238 13539 3290
rect 13539 3238 13585 3290
rect 13609 3238 13655 3290
rect 13655 3238 13665 3290
rect 13689 3238 13719 3290
rect 13719 3238 13745 3290
rect 13449 3236 13505 3238
rect 13529 3236 13585 3238
rect 13609 3236 13665 3238
rect 13689 3236 13745 3238
rect 13449 2202 13505 2204
rect 13529 2202 13585 2204
rect 13609 2202 13665 2204
rect 13689 2202 13745 2204
rect 13449 2150 13475 2202
rect 13475 2150 13505 2202
rect 13529 2150 13539 2202
rect 13539 2150 13585 2202
rect 13609 2150 13655 2202
rect 13655 2150 13665 2202
rect 13689 2150 13719 2202
rect 13719 2150 13745 2202
rect 13449 2148 13505 2150
rect 13529 2148 13585 2150
rect 13609 2148 13665 2150
rect 13689 2148 13745 2150
rect 14462 2488 14518 2544
<< metal3 >>
rect 10225 19138 10291 19141
rect 10358 19138 10364 19140
rect 10225 19136 10364 19138
rect 10225 19080 10230 19136
rect 10286 19080 10364 19136
rect 10225 19078 10364 19080
rect 10225 19075 10291 19078
rect 10358 19076 10364 19078
rect 10428 19076 10434 19140
rect 0 18322 800 18352
rect 4061 18322 4127 18325
rect 0 18320 4127 18322
rect 0 18264 4066 18320
rect 4122 18264 4127 18320
rect 0 18262 4127 18264
rect 0 18232 800 18262
rect 4061 18259 4127 18262
rect 15469 17506 15535 17509
rect 16400 17506 17200 17536
rect 15469 17504 17200 17506
rect 15469 17448 15474 17504
rect 15530 17448 17200 17504
rect 15469 17446 17200 17448
rect 15469 17443 15535 17446
rect 3442 17440 3762 17441
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3762 17440
rect 3442 17375 3762 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 13437 17440 13757 17441
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 16400 17416 17200 17446
rect 13437 17375 13757 17376
rect 5941 16896 6261 16897
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 16831 6261 16832
rect 10938 16896 11258 16897
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11258 16896
rect 10938 16831 11258 16832
rect 3442 16352 3762 16353
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3762 16352
rect 3442 16287 3762 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 13437 16352 13757 16353
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 16287 13757 16288
rect 5941 15808 6261 15809
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 15743 6261 15744
rect 10938 15808 11258 15809
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11258 15808
rect 10938 15743 11258 15744
rect 3442 15264 3762 15265
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3762 15264
rect 3442 15199 3762 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 13437 15264 13757 15265
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 15199 13757 15200
rect 0 15058 800 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 800 14998
rect 2773 14995 2839 14998
rect 5941 14720 6261 14721
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 14655 6261 14656
rect 10938 14720 11258 14721
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11258 14720
rect 10938 14655 11258 14656
rect 3442 14176 3762 14177
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3762 14176
rect 3442 14111 3762 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 13437 14176 13757 14177
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 14111 13757 14112
rect 5941 13632 6261 13633
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 13567 6261 13568
rect 10938 13632 11258 13633
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11258 13632
rect 10938 13567 11258 13568
rect 3442 13088 3762 13089
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3762 13088
rect 3442 13023 3762 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 13437 13088 13757 13089
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 13023 13757 13024
rect 5941 12544 6261 12545
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 12479 6261 12480
rect 10938 12544 11258 12545
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11258 12544
rect 10938 12479 11258 12480
rect 13721 12474 13787 12477
rect 16400 12474 17200 12504
rect 13721 12472 17200 12474
rect 13721 12416 13726 12472
rect 13782 12416 17200 12472
rect 13721 12414 17200 12416
rect 13721 12411 13787 12414
rect 16400 12384 17200 12414
rect 3442 12000 3762 12001
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3762 12000
rect 3442 11935 3762 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 13437 12000 13757 12001
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 11935 13757 11936
rect 0 11658 800 11688
rect 3325 11658 3391 11661
rect 0 11656 3391 11658
rect 0 11600 3330 11656
rect 3386 11600 3391 11656
rect 0 11598 3391 11600
rect 0 11568 800 11598
rect 3325 11595 3391 11598
rect 5941 11456 6261 11457
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 11391 6261 11392
rect 10938 11456 11258 11457
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11258 11456
rect 10938 11391 11258 11392
rect 3442 10912 3762 10913
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3762 10912
rect 3442 10847 3762 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 13437 10912 13757 10913
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 10847 13757 10848
rect 5941 10368 6261 10369
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 10303 6261 10304
rect 10938 10368 11258 10369
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11258 10368
rect 10938 10303 11258 10304
rect 10358 9964 10364 10028
rect 10428 10026 10434 10028
rect 10501 10026 10567 10029
rect 10428 10024 10567 10026
rect 10428 9968 10506 10024
rect 10562 9968 10567 10024
rect 10428 9966 10567 9968
rect 10428 9964 10434 9966
rect 10501 9963 10567 9966
rect 3442 9824 3762 9825
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3762 9824
rect 3442 9759 3762 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 13437 9824 13757 9825
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 9759 13757 9760
rect 9489 9618 9555 9621
rect 9262 9616 9555 9618
rect 9262 9560 9494 9616
rect 9550 9560 9555 9616
rect 9262 9558 9555 9560
rect 9262 9346 9322 9558
rect 9489 9555 9555 9558
rect 10225 9618 10291 9621
rect 10358 9618 10364 9620
rect 10225 9616 10364 9618
rect 10225 9560 10230 9616
rect 10286 9560 10364 9616
rect 10225 9558 10364 9560
rect 10225 9555 10291 9558
rect 10358 9556 10364 9558
rect 10428 9556 10434 9620
rect 9438 9420 9444 9484
rect 9508 9482 9514 9484
rect 9581 9482 9647 9485
rect 9508 9480 9647 9482
rect 9508 9424 9586 9480
rect 9642 9424 9647 9480
rect 9508 9422 9647 9424
rect 9508 9420 9514 9422
rect 9581 9419 9647 9422
rect 9581 9346 9647 9349
rect 9262 9344 9647 9346
rect 9262 9288 9586 9344
rect 9642 9288 9647 9344
rect 9262 9286 9647 9288
rect 9581 9283 9647 9286
rect 5941 9280 6261 9281
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 9215 6261 9216
rect 10938 9280 11258 9281
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11258 9280
rect 10938 9215 11258 9216
rect 3442 8736 3762 8737
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3762 8736
rect 3442 8671 3762 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 13437 8736 13757 8737
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 8671 13757 8672
rect 0 8394 800 8424
rect 1485 8394 1551 8397
rect 0 8392 1551 8394
rect 0 8336 1490 8392
rect 1546 8336 1551 8392
rect 0 8334 1551 8336
rect 0 8304 800 8334
rect 1485 8331 1551 8334
rect 5941 8192 6261 8193
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 8127 6261 8128
rect 10938 8192 11258 8193
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11258 8192
rect 10938 8127 11258 8128
rect 3442 7648 3762 7649
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3762 7648
rect 3442 7583 3762 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 13437 7648 13757 7649
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 7583 13757 7584
rect 13353 7442 13419 7445
rect 16400 7442 17200 7472
rect 13353 7440 17200 7442
rect 13353 7384 13358 7440
rect 13414 7384 17200 7440
rect 13353 7382 17200 7384
rect 13353 7379 13419 7382
rect 16400 7352 17200 7382
rect 5941 7104 6261 7105
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 7039 6261 7040
rect 10938 7104 11258 7105
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11258 7104
rect 10938 7039 11258 7040
rect 3442 6560 3762 6561
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3762 6560
rect 3442 6495 3762 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 13437 6560 13757 6561
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 6495 13757 6496
rect 5941 6016 6261 6017
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 5951 6261 5952
rect 10938 6016 11258 6017
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11258 6016
rect 10938 5951 11258 5952
rect 3442 5472 3762 5473
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3762 5472
rect 3442 5407 3762 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 13437 5472 13757 5473
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 5407 13757 5408
rect 9397 5402 9463 5405
rect 12893 5402 12959 5405
rect 9397 5400 12959 5402
rect 9397 5344 9402 5400
rect 9458 5344 12898 5400
rect 12954 5344 12959 5400
rect 9397 5342 12959 5344
rect 9397 5339 9463 5342
rect 12893 5339 12959 5342
rect 6821 5266 6887 5269
rect 11053 5266 11119 5269
rect 6821 5264 11119 5266
rect 6821 5208 6826 5264
rect 6882 5208 11058 5264
rect 11114 5208 11119 5264
rect 6821 5206 11119 5208
rect 6821 5203 6887 5206
rect 11053 5203 11119 5206
rect 8201 5130 8267 5133
rect 12617 5130 12683 5133
rect 8201 5128 12683 5130
rect 8201 5072 8206 5128
rect 8262 5072 12622 5128
rect 12678 5072 12683 5128
rect 8201 5070 12683 5072
rect 8201 5067 8267 5070
rect 12617 5067 12683 5070
rect 0 4994 800 5024
rect 2957 4994 3023 4997
rect 0 4992 3023 4994
rect 0 4936 2962 4992
rect 3018 4936 3023 4992
rect 0 4934 3023 4936
rect 0 4904 800 4934
rect 2957 4931 3023 4934
rect 5941 4928 6261 4929
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 4863 6261 4864
rect 10938 4928 11258 4929
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11258 4928
rect 10938 4863 11258 4864
rect 3442 4384 3762 4385
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3762 4384
rect 3442 4319 3762 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 13437 4384 13757 4385
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 4319 13757 4320
rect 5941 3840 6261 3841
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 3775 6261 3776
rect 10938 3840 11258 3841
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11258 3840
rect 10938 3775 11258 3776
rect 3442 3296 3762 3297
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3762 3296
rect 3442 3231 3762 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 13437 3296 13757 3297
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 3231 13757 3232
rect 5941 2752 6261 2753
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2687 6261 2688
rect 10938 2752 11258 2753
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11258 2752
rect 10938 2687 11258 2688
rect 14457 2546 14523 2549
rect 16400 2546 17200 2576
rect 14457 2544 17200 2546
rect 14457 2488 14462 2544
rect 14518 2488 17200 2544
rect 14457 2486 17200 2488
rect 14457 2483 14523 2486
rect 16400 2456 17200 2486
rect 3442 2208 3762 2209
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3762 2208
rect 3442 2143 3762 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 13437 2208 13757 2209
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2143 13757 2144
rect 0 1730 800 1760
rect 1577 1730 1643 1733
rect 0 1728 1643 1730
rect 0 1672 1582 1728
rect 1638 1672 1643 1728
rect 0 1670 1643 1672
rect 0 1640 800 1670
rect 1577 1667 1643 1670
rect 5349 914 5415 917
rect 9121 914 9187 917
rect 5349 912 9187 914
rect 5349 856 5354 912
rect 5410 856 9126 912
rect 9182 856 9187 912
rect 5349 854 9187 856
rect 5349 851 5415 854
rect 9121 851 9187 854
rect 9438 852 9444 916
rect 9508 914 9514 916
rect 9581 914 9647 917
rect 9508 912 9647 914
rect 9508 856 9586 912
rect 9642 856 9647 912
rect 9508 854 9647 856
rect 9508 852 9514 854
rect 9581 851 9647 854
rect 10358 852 10364 916
rect 10428 914 10434 916
rect 10501 914 10567 917
rect 10428 912 10567 914
rect 10428 856 10506 912
rect 10562 856 10567 912
rect 10428 854 10567 856
rect 10428 852 10434 854
rect 10501 851 10567 854
<< via3 >>
rect 10364 19076 10428 19140
rect 3450 17436 3514 17440
rect 3450 17380 3454 17436
rect 3454 17380 3510 17436
rect 3510 17380 3514 17436
rect 3450 17376 3514 17380
rect 3530 17436 3594 17440
rect 3530 17380 3534 17436
rect 3534 17380 3590 17436
rect 3590 17380 3594 17436
rect 3530 17376 3594 17380
rect 3610 17436 3674 17440
rect 3610 17380 3614 17436
rect 3614 17380 3670 17436
rect 3670 17380 3674 17436
rect 3610 17376 3674 17380
rect 3690 17436 3754 17440
rect 3690 17380 3694 17436
rect 3694 17380 3750 17436
rect 3750 17380 3754 17436
rect 3690 17376 3754 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 13445 17436 13509 17440
rect 13445 17380 13449 17436
rect 13449 17380 13505 17436
rect 13505 17380 13509 17436
rect 13445 17376 13509 17380
rect 13525 17436 13589 17440
rect 13525 17380 13529 17436
rect 13529 17380 13585 17436
rect 13585 17380 13589 17436
rect 13525 17376 13589 17380
rect 13605 17436 13669 17440
rect 13605 17380 13609 17436
rect 13609 17380 13665 17436
rect 13665 17380 13669 17436
rect 13605 17376 13669 17380
rect 13685 17436 13749 17440
rect 13685 17380 13689 17436
rect 13689 17380 13745 17436
rect 13745 17380 13749 17436
rect 13685 17376 13749 17380
rect 5949 16892 6013 16896
rect 5949 16836 5953 16892
rect 5953 16836 6009 16892
rect 6009 16836 6013 16892
rect 5949 16832 6013 16836
rect 6029 16892 6093 16896
rect 6029 16836 6033 16892
rect 6033 16836 6089 16892
rect 6089 16836 6093 16892
rect 6029 16832 6093 16836
rect 6109 16892 6173 16896
rect 6109 16836 6113 16892
rect 6113 16836 6169 16892
rect 6169 16836 6173 16892
rect 6109 16832 6173 16836
rect 6189 16892 6253 16896
rect 6189 16836 6193 16892
rect 6193 16836 6249 16892
rect 6249 16836 6253 16892
rect 6189 16832 6253 16836
rect 10946 16892 11010 16896
rect 10946 16836 10950 16892
rect 10950 16836 11006 16892
rect 11006 16836 11010 16892
rect 10946 16832 11010 16836
rect 11026 16892 11090 16896
rect 11026 16836 11030 16892
rect 11030 16836 11086 16892
rect 11086 16836 11090 16892
rect 11026 16832 11090 16836
rect 11106 16892 11170 16896
rect 11106 16836 11110 16892
rect 11110 16836 11166 16892
rect 11166 16836 11170 16892
rect 11106 16832 11170 16836
rect 11186 16892 11250 16896
rect 11186 16836 11190 16892
rect 11190 16836 11246 16892
rect 11246 16836 11250 16892
rect 11186 16832 11250 16836
rect 3450 16348 3514 16352
rect 3450 16292 3454 16348
rect 3454 16292 3510 16348
rect 3510 16292 3514 16348
rect 3450 16288 3514 16292
rect 3530 16348 3594 16352
rect 3530 16292 3534 16348
rect 3534 16292 3590 16348
rect 3590 16292 3594 16348
rect 3530 16288 3594 16292
rect 3610 16348 3674 16352
rect 3610 16292 3614 16348
rect 3614 16292 3670 16348
rect 3670 16292 3674 16348
rect 3610 16288 3674 16292
rect 3690 16348 3754 16352
rect 3690 16292 3694 16348
rect 3694 16292 3750 16348
rect 3750 16292 3754 16348
rect 3690 16288 3754 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 13445 16348 13509 16352
rect 13445 16292 13449 16348
rect 13449 16292 13505 16348
rect 13505 16292 13509 16348
rect 13445 16288 13509 16292
rect 13525 16348 13589 16352
rect 13525 16292 13529 16348
rect 13529 16292 13585 16348
rect 13585 16292 13589 16348
rect 13525 16288 13589 16292
rect 13605 16348 13669 16352
rect 13605 16292 13609 16348
rect 13609 16292 13665 16348
rect 13665 16292 13669 16348
rect 13605 16288 13669 16292
rect 13685 16348 13749 16352
rect 13685 16292 13689 16348
rect 13689 16292 13745 16348
rect 13745 16292 13749 16348
rect 13685 16288 13749 16292
rect 5949 15804 6013 15808
rect 5949 15748 5953 15804
rect 5953 15748 6009 15804
rect 6009 15748 6013 15804
rect 5949 15744 6013 15748
rect 6029 15804 6093 15808
rect 6029 15748 6033 15804
rect 6033 15748 6089 15804
rect 6089 15748 6093 15804
rect 6029 15744 6093 15748
rect 6109 15804 6173 15808
rect 6109 15748 6113 15804
rect 6113 15748 6169 15804
rect 6169 15748 6173 15804
rect 6109 15744 6173 15748
rect 6189 15804 6253 15808
rect 6189 15748 6193 15804
rect 6193 15748 6249 15804
rect 6249 15748 6253 15804
rect 6189 15744 6253 15748
rect 10946 15804 11010 15808
rect 10946 15748 10950 15804
rect 10950 15748 11006 15804
rect 11006 15748 11010 15804
rect 10946 15744 11010 15748
rect 11026 15804 11090 15808
rect 11026 15748 11030 15804
rect 11030 15748 11086 15804
rect 11086 15748 11090 15804
rect 11026 15744 11090 15748
rect 11106 15804 11170 15808
rect 11106 15748 11110 15804
rect 11110 15748 11166 15804
rect 11166 15748 11170 15804
rect 11106 15744 11170 15748
rect 11186 15804 11250 15808
rect 11186 15748 11190 15804
rect 11190 15748 11246 15804
rect 11246 15748 11250 15804
rect 11186 15744 11250 15748
rect 3450 15260 3514 15264
rect 3450 15204 3454 15260
rect 3454 15204 3510 15260
rect 3510 15204 3514 15260
rect 3450 15200 3514 15204
rect 3530 15260 3594 15264
rect 3530 15204 3534 15260
rect 3534 15204 3590 15260
rect 3590 15204 3594 15260
rect 3530 15200 3594 15204
rect 3610 15260 3674 15264
rect 3610 15204 3614 15260
rect 3614 15204 3670 15260
rect 3670 15204 3674 15260
rect 3610 15200 3674 15204
rect 3690 15260 3754 15264
rect 3690 15204 3694 15260
rect 3694 15204 3750 15260
rect 3750 15204 3754 15260
rect 3690 15200 3754 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 13445 15260 13509 15264
rect 13445 15204 13449 15260
rect 13449 15204 13505 15260
rect 13505 15204 13509 15260
rect 13445 15200 13509 15204
rect 13525 15260 13589 15264
rect 13525 15204 13529 15260
rect 13529 15204 13585 15260
rect 13585 15204 13589 15260
rect 13525 15200 13589 15204
rect 13605 15260 13669 15264
rect 13605 15204 13609 15260
rect 13609 15204 13665 15260
rect 13665 15204 13669 15260
rect 13605 15200 13669 15204
rect 13685 15260 13749 15264
rect 13685 15204 13689 15260
rect 13689 15204 13745 15260
rect 13745 15204 13749 15260
rect 13685 15200 13749 15204
rect 5949 14716 6013 14720
rect 5949 14660 5953 14716
rect 5953 14660 6009 14716
rect 6009 14660 6013 14716
rect 5949 14656 6013 14660
rect 6029 14716 6093 14720
rect 6029 14660 6033 14716
rect 6033 14660 6089 14716
rect 6089 14660 6093 14716
rect 6029 14656 6093 14660
rect 6109 14716 6173 14720
rect 6109 14660 6113 14716
rect 6113 14660 6169 14716
rect 6169 14660 6173 14716
rect 6109 14656 6173 14660
rect 6189 14716 6253 14720
rect 6189 14660 6193 14716
rect 6193 14660 6249 14716
rect 6249 14660 6253 14716
rect 6189 14656 6253 14660
rect 10946 14716 11010 14720
rect 10946 14660 10950 14716
rect 10950 14660 11006 14716
rect 11006 14660 11010 14716
rect 10946 14656 11010 14660
rect 11026 14716 11090 14720
rect 11026 14660 11030 14716
rect 11030 14660 11086 14716
rect 11086 14660 11090 14716
rect 11026 14656 11090 14660
rect 11106 14716 11170 14720
rect 11106 14660 11110 14716
rect 11110 14660 11166 14716
rect 11166 14660 11170 14716
rect 11106 14656 11170 14660
rect 11186 14716 11250 14720
rect 11186 14660 11190 14716
rect 11190 14660 11246 14716
rect 11246 14660 11250 14716
rect 11186 14656 11250 14660
rect 3450 14172 3514 14176
rect 3450 14116 3454 14172
rect 3454 14116 3510 14172
rect 3510 14116 3514 14172
rect 3450 14112 3514 14116
rect 3530 14172 3594 14176
rect 3530 14116 3534 14172
rect 3534 14116 3590 14172
rect 3590 14116 3594 14172
rect 3530 14112 3594 14116
rect 3610 14172 3674 14176
rect 3610 14116 3614 14172
rect 3614 14116 3670 14172
rect 3670 14116 3674 14172
rect 3610 14112 3674 14116
rect 3690 14172 3754 14176
rect 3690 14116 3694 14172
rect 3694 14116 3750 14172
rect 3750 14116 3754 14172
rect 3690 14112 3754 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 13445 14172 13509 14176
rect 13445 14116 13449 14172
rect 13449 14116 13505 14172
rect 13505 14116 13509 14172
rect 13445 14112 13509 14116
rect 13525 14172 13589 14176
rect 13525 14116 13529 14172
rect 13529 14116 13585 14172
rect 13585 14116 13589 14172
rect 13525 14112 13589 14116
rect 13605 14172 13669 14176
rect 13605 14116 13609 14172
rect 13609 14116 13665 14172
rect 13665 14116 13669 14172
rect 13605 14112 13669 14116
rect 13685 14172 13749 14176
rect 13685 14116 13689 14172
rect 13689 14116 13745 14172
rect 13745 14116 13749 14172
rect 13685 14112 13749 14116
rect 5949 13628 6013 13632
rect 5949 13572 5953 13628
rect 5953 13572 6009 13628
rect 6009 13572 6013 13628
rect 5949 13568 6013 13572
rect 6029 13628 6093 13632
rect 6029 13572 6033 13628
rect 6033 13572 6089 13628
rect 6089 13572 6093 13628
rect 6029 13568 6093 13572
rect 6109 13628 6173 13632
rect 6109 13572 6113 13628
rect 6113 13572 6169 13628
rect 6169 13572 6173 13628
rect 6109 13568 6173 13572
rect 6189 13628 6253 13632
rect 6189 13572 6193 13628
rect 6193 13572 6249 13628
rect 6249 13572 6253 13628
rect 6189 13568 6253 13572
rect 10946 13628 11010 13632
rect 10946 13572 10950 13628
rect 10950 13572 11006 13628
rect 11006 13572 11010 13628
rect 10946 13568 11010 13572
rect 11026 13628 11090 13632
rect 11026 13572 11030 13628
rect 11030 13572 11086 13628
rect 11086 13572 11090 13628
rect 11026 13568 11090 13572
rect 11106 13628 11170 13632
rect 11106 13572 11110 13628
rect 11110 13572 11166 13628
rect 11166 13572 11170 13628
rect 11106 13568 11170 13572
rect 11186 13628 11250 13632
rect 11186 13572 11190 13628
rect 11190 13572 11246 13628
rect 11246 13572 11250 13628
rect 11186 13568 11250 13572
rect 3450 13084 3514 13088
rect 3450 13028 3454 13084
rect 3454 13028 3510 13084
rect 3510 13028 3514 13084
rect 3450 13024 3514 13028
rect 3530 13084 3594 13088
rect 3530 13028 3534 13084
rect 3534 13028 3590 13084
rect 3590 13028 3594 13084
rect 3530 13024 3594 13028
rect 3610 13084 3674 13088
rect 3610 13028 3614 13084
rect 3614 13028 3670 13084
rect 3670 13028 3674 13084
rect 3610 13024 3674 13028
rect 3690 13084 3754 13088
rect 3690 13028 3694 13084
rect 3694 13028 3750 13084
rect 3750 13028 3754 13084
rect 3690 13024 3754 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 13445 13084 13509 13088
rect 13445 13028 13449 13084
rect 13449 13028 13505 13084
rect 13505 13028 13509 13084
rect 13445 13024 13509 13028
rect 13525 13084 13589 13088
rect 13525 13028 13529 13084
rect 13529 13028 13585 13084
rect 13585 13028 13589 13084
rect 13525 13024 13589 13028
rect 13605 13084 13669 13088
rect 13605 13028 13609 13084
rect 13609 13028 13665 13084
rect 13665 13028 13669 13084
rect 13605 13024 13669 13028
rect 13685 13084 13749 13088
rect 13685 13028 13689 13084
rect 13689 13028 13745 13084
rect 13745 13028 13749 13084
rect 13685 13024 13749 13028
rect 5949 12540 6013 12544
rect 5949 12484 5953 12540
rect 5953 12484 6009 12540
rect 6009 12484 6013 12540
rect 5949 12480 6013 12484
rect 6029 12540 6093 12544
rect 6029 12484 6033 12540
rect 6033 12484 6089 12540
rect 6089 12484 6093 12540
rect 6029 12480 6093 12484
rect 6109 12540 6173 12544
rect 6109 12484 6113 12540
rect 6113 12484 6169 12540
rect 6169 12484 6173 12540
rect 6109 12480 6173 12484
rect 6189 12540 6253 12544
rect 6189 12484 6193 12540
rect 6193 12484 6249 12540
rect 6249 12484 6253 12540
rect 6189 12480 6253 12484
rect 10946 12540 11010 12544
rect 10946 12484 10950 12540
rect 10950 12484 11006 12540
rect 11006 12484 11010 12540
rect 10946 12480 11010 12484
rect 11026 12540 11090 12544
rect 11026 12484 11030 12540
rect 11030 12484 11086 12540
rect 11086 12484 11090 12540
rect 11026 12480 11090 12484
rect 11106 12540 11170 12544
rect 11106 12484 11110 12540
rect 11110 12484 11166 12540
rect 11166 12484 11170 12540
rect 11106 12480 11170 12484
rect 11186 12540 11250 12544
rect 11186 12484 11190 12540
rect 11190 12484 11246 12540
rect 11246 12484 11250 12540
rect 11186 12480 11250 12484
rect 3450 11996 3514 12000
rect 3450 11940 3454 11996
rect 3454 11940 3510 11996
rect 3510 11940 3514 11996
rect 3450 11936 3514 11940
rect 3530 11996 3594 12000
rect 3530 11940 3534 11996
rect 3534 11940 3590 11996
rect 3590 11940 3594 11996
rect 3530 11936 3594 11940
rect 3610 11996 3674 12000
rect 3610 11940 3614 11996
rect 3614 11940 3670 11996
rect 3670 11940 3674 11996
rect 3610 11936 3674 11940
rect 3690 11996 3754 12000
rect 3690 11940 3694 11996
rect 3694 11940 3750 11996
rect 3750 11940 3754 11996
rect 3690 11936 3754 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 13445 11996 13509 12000
rect 13445 11940 13449 11996
rect 13449 11940 13505 11996
rect 13505 11940 13509 11996
rect 13445 11936 13509 11940
rect 13525 11996 13589 12000
rect 13525 11940 13529 11996
rect 13529 11940 13585 11996
rect 13585 11940 13589 11996
rect 13525 11936 13589 11940
rect 13605 11996 13669 12000
rect 13605 11940 13609 11996
rect 13609 11940 13665 11996
rect 13665 11940 13669 11996
rect 13605 11936 13669 11940
rect 13685 11996 13749 12000
rect 13685 11940 13689 11996
rect 13689 11940 13745 11996
rect 13745 11940 13749 11996
rect 13685 11936 13749 11940
rect 5949 11452 6013 11456
rect 5949 11396 5953 11452
rect 5953 11396 6009 11452
rect 6009 11396 6013 11452
rect 5949 11392 6013 11396
rect 6029 11452 6093 11456
rect 6029 11396 6033 11452
rect 6033 11396 6089 11452
rect 6089 11396 6093 11452
rect 6029 11392 6093 11396
rect 6109 11452 6173 11456
rect 6109 11396 6113 11452
rect 6113 11396 6169 11452
rect 6169 11396 6173 11452
rect 6109 11392 6173 11396
rect 6189 11452 6253 11456
rect 6189 11396 6193 11452
rect 6193 11396 6249 11452
rect 6249 11396 6253 11452
rect 6189 11392 6253 11396
rect 10946 11452 11010 11456
rect 10946 11396 10950 11452
rect 10950 11396 11006 11452
rect 11006 11396 11010 11452
rect 10946 11392 11010 11396
rect 11026 11452 11090 11456
rect 11026 11396 11030 11452
rect 11030 11396 11086 11452
rect 11086 11396 11090 11452
rect 11026 11392 11090 11396
rect 11106 11452 11170 11456
rect 11106 11396 11110 11452
rect 11110 11396 11166 11452
rect 11166 11396 11170 11452
rect 11106 11392 11170 11396
rect 11186 11452 11250 11456
rect 11186 11396 11190 11452
rect 11190 11396 11246 11452
rect 11246 11396 11250 11452
rect 11186 11392 11250 11396
rect 3450 10908 3514 10912
rect 3450 10852 3454 10908
rect 3454 10852 3510 10908
rect 3510 10852 3514 10908
rect 3450 10848 3514 10852
rect 3530 10908 3594 10912
rect 3530 10852 3534 10908
rect 3534 10852 3590 10908
rect 3590 10852 3594 10908
rect 3530 10848 3594 10852
rect 3610 10908 3674 10912
rect 3610 10852 3614 10908
rect 3614 10852 3670 10908
rect 3670 10852 3674 10908
rect 3610 10848 3674 10852
rect 3690 10908 3754 10912
rect 3690 10852 3694 10908
rect 3694 10852 3750 10908
rect 3750 10852 3754 10908
rect 3690 10848 3754 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 13445 10908 13509 10912
rect 13445 10852 13449 10908
rect 13449 10852 13505 10908
rect 13505 10852 13509 10908
rect 13445 10848 13509 10852
rect 13525 10908 13589 10912
rect 13525 10852 13529 10908
rect 13529 10852 13585 10908
rect 13585 10852 13589 10908
rect 13525 10848 13589 10852
rect 13605 10908 13669 10912
rect 13605 10852 13609 10908
rect 13609 10852 13665 10908
rect 13665 10852 13669 10908
rect 13605 10848 13669 10852
rect 13685 10908 13749 10912
rect 13685 10852 13689 10908
rect 13689 10852 13745 10908
rect 13745 10852 13749 10908
rect 13685 10848 13749 10852
rect 5949 10364 6013 10368
rect 5949 10308 5953 10364
rect 5953 10308 6009 10364
rect 6009 10308 6013 10364
rect 5949 10304 6013 10308
rect 6029 10364 6093 10368
rect 6029 10308 6033 10364
rect 6033 10308 6089 10364
rect 6089 10308 6093 10364
rect 6029 10304 6093 10308
rect 6109 10364 6173 10368
rect 6109 10308 6113 10364
rect 6113 10308 6169 10364
rect 6169 10308 6173 10364
rect 6109 10304 6173 10308
rect 6189 10364 6253 10368
rect 6189 10308 6193 10364
rect 6193 10308 6249 10364
rect 6249 10308 6253 10364
rect 6189 10304 6253 10308
rect 10946 10364 11010 10368
rect 10946 10308 10950 10364
rect 10950 10308 11006 10364
rect 11006 10308 11010 10364
rect 10946 10304 11010 10308
rect 11026 10364 11090 10368
rect 11026 10308 11030 10364
rect 11030 10308 11086 10364
rect 11086 10308 11090 10364
rect 11026 10304 11090 10308
rect 11106 10364 11170 10368
rect 11106 10308 11110 10364
rect 11110 10308 11166 10364
rect 11166 10308 11170 10364
rect 11106 10304 11170 10308
rect 11186 10364 11250 10368
rect 11186 10308 11190 10364
rect 11190 10308 11246 10364
rect 11246 10308 11250 10364
rect 11186 10304 11250 10308
rect 10364 9964 10428 10028
rect 3450 9820 3514 9824
rect 3450 9764 3454 9820
rect 3454 9764 3510 9820
rect 3510 9764 3514 9820
rect 3450 9760 3514 9764
rect 3530 9820 3594 9824
rect 3530 9764 3534 9820
rect 3534 9764 3590 9820
rect 3590 9764 3594 9820
rect 3530 9760 3594 9764
rect 3610 9820 3674 9824
rect 3610 9764 3614 9820
rect 3614 9764 3670 9820
rect 3670 9764 3674 9820
rect 3610 9760 3674 9764
rect 3690 9820 3754 9824
rect 3690 9764 3694 9820
rect 3694 9764 3750 9820
rect 3750 9764 3754 9820
rect 3690 9760 3754 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 13445 9820 13509 9824
rect 13445 9764 13449 9820
rect 13449 9764 13505 9820
rect 13505 9764 13509 9820
rect 13445 9760 13509 9764
rect 13525 9820 13589 9824
rect 13525 9764 13529 9820
rect 13529 9764 13585 9820
rect 13585 9764 13589 9820
rect 13525 9760 13589 9764
rect 13605 9820 13669 9824
rect 13605 9764 13609 9820
rect 13609 9764 13665 9820
rect 13665 9764 13669 9820
rect 13605 9760 13669 9764
rect 13685 9820 13749 9824
rect 13685 9764 13689 9820
rect 13689 9764 13745 9820
rect 13745 9764 13749 9820
rect 13685 9760 13749 9764
rect 10364 9556 10428 9620
rect 9444 9420 9508 9484
rect 5949 9276 6013 9280
rect 5949 9220 5953 9276
rect 5953 9220 6009 9276
rect 6009 9220 6013 9276
rect 5949 9216 6013 9220
rect 6029 9276 6093 9280
rect 6029 9220 6033 9276
rect 6033 9220 6089 9276
rect 6089 9220 6093 9276
rect 6029 9216 6093 9220
rect 6109 9276 6173 9280
rect 6109 9220 6113 9276
rect 6113 9220 6169 9276
rect 6169 9220 6173 9276
rect 6109 9216 6173 9220
rect 6189 9276 6253 9280
rect 6189 9220 6193 9276
rect 6193 9220 6249 9276
rect 6249 9220 6253 9276
rect 6189 9216 6253 9220
rect 10946 9276 11010 9280
rect 10946 9220 10950 9276
rect 10950 9220 11006 9276
rect 11006 9220 11010 9276
rect 10946 9216 11010 9220
rect 11026 9276 11090 9280
rect 11026 9220 11030 9276
rect 11030 9220 11086 9276
rect 11086 9220 11090 9276
rect 11026 9216 11090 9220
rect 11106 9276 11170 9280
rect 11106 9220 11110 9276
rect 11110 9220 11166 9276
rect 11166 9220 11170 9276
rect 11106 9216 11170 9220
rect 11186 9276 11250 9280
rect 11186 9220 11190 9276
rect 11190 9220 11246 9276
rect 11246 9220 11250 9276
rect 11186 9216 11250 9220
rect 3450 8732 3514 8736
rect 3450 8676 3454 8732
rect 3454 8676 3510 8732
rect 3510 8676 3514 8732
rect 3450 8672 3514 8676
rect 3530 8732 3594 8736
rect 3530 8676 3534 8732
rect 3534 8676 3590 8732
rect 3590 8676 3594 8732
rect 3530 8672 3594 8676
rect 3610 8732 3674 8736
rect 3610 8676 3614 8732
rect 3614 8676 3670 8732
rect 3670 8676 3674 8732
rect 3610 8672 3674 8676
rect 3690 8732 3754 8736
rect 3690 8676 3694 8732
rect 3694 8676 3750 8732
rect 3750 8676 3754 8732
rect 3690 8672 3754 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 13445 8732 13509 8736
rect 13445 8676 13449 8732
rect 13449 8676 13505 8732
rect 13505 8676 13509 8732
rect 13445 8672 13509 8676
rect 13525 8732 13589 8736
rect 13525 8676 13529 8732
rect 13529 8676 13585 8732
rect 13585 8676 13589 8732
rect 13525 8672 13589 8676
rect 13605 8732 13669 8736
rect 13605 8676 13609 8732
rect 13609 8676 13665 8732
rect 13665 8676 13669 8732
rect 13605 8672 13669 8676
rect 13685 8732 13749 8736
rect 13685 8676 13689 8732
rect 13689 8676 13745 8732
rect 13745 8676 13749 8732
rect 13685 8672 13749 8676
rect 5949 8188 6013 8192
rect 5949 8132 5953 8188
rect 5953 8132 6009 8188
rect 6009 8132 6013 8188
rect 5949 8128 6013 8132
rect 6029 8188 6093 8192
rect 6029 8132 6033 8188
rect 6033 8132 6089 8188
rect 6089 8132 6093 8188
rect 6029 8128 6093 8132
rect 6109 8188 6173 8192
rect 6109 8132 6113 8188
rect 6113 8132 6169 8188
rect 6169 8132 6173 8188
rect 6109 8128 6173 8132
rect 6189 8188 6253 8192
rect 6189 8132 6193 8188
rect 6193 8132 6249 8188
rect 6249 8132 6253 8188
rect 6189 8128 6253 8132
rect 10946 8188 11010 8192
rect 10946 8132 10950 8188
rect 10950 8132 11006 8188
rect 11006 8132 11010 8188
rect 10946 8128 11010 8132
rect 11026 8188 11090 8192
rect 11026 8132 11030 8188
rect 11030 8132 11086 8188
rect 11086 8132 11090 8188
rect 11026 8128 11090 8132
rect 11106 8188 11170 8192
rect 11106 8132 11110 8188
rect 11110 8132 11166 8188
rect 11166 8132 11170 8188
rect 11106 8128 11170 8132
rect 11186 8188 11250 8192
rect 11186 8132 11190 8188
rect 11190 8132 11246 8188
rect 11246 8132 11250 8188
rect 11186 8128 11250 8132
rect 3450 7644 3514 7648
rect 3450 7588 3454 7644
rect 3454 7588 3510 7644
rect 3510 7588 3514 7644
rect 3450 7584 3514 7588
rect 3530 7644 3594 7648
rect 3530 7588 3534 7644
rect 3534 7588 3590 7644
rect 3590 7588 3594 7644
rect 3530 7584 3594 7588
rect 3610 7644 3674 7648
rect 3610 7588 3614 7644
rect 3614 7588 3670 7644
rect 3670 7588 3674 7644
rect 3610 7584 3674 7588
rect 3690 7644 3754 7648
rect 3690 7588 3694 7644
rect 3694 7588 3750 7644
rect 3750 7588 3754 7644
rect 3690 7584 3754 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 13445 7644 13509 7648
rect 13445 7588 13449 7644
rect 13449 7588 13505 7644
rect 13505 7588 13509 7644
rect 13445 7584 13509 7588
rect 13525 7644 13589 7648
rect 13525 7588 13529 7644
rect 13529 7588 13585 7644
rect 13585 7588 13589 7644
rect 13525 7584 13589 7588
rect 13605 7644 13669 7648
rect 13605 7588 13609 7644
rect 13609 7588 13665 7644
rect 13665 7588 13669 7644
rect 13605 7584 13669 7588
rect 13685 7644 13749 7648
rect 13685 7588 13689 7644
rect 13689 7588 13745 7644
rect 13745 7588 13749 7644
rect 13685 7584 13749 7588
rect 5949 7100 6013 7104
rect 5949 7044 5953 7100
rect 5953 7044 6009 7100
rect 6009 7044 6013 7100
rect 5949 7040 6013 7044
rect 6029 7100 6093 7104
rect 6029 7044 6033 7100
rect 6033 7044 6089 7100
rect 6089 7044 6093 7100
rect 6029 7040 6093 7044
rect 6109 7100 6173 7104
rect 6109 7044 6113 7100
rect 6113 7044 6169 7100
rect 6169 7044 6173 7100
rect 6109 7040 6173 7044
rect 6189 7100 6253 7104
rect 6189 7044 6193 7100
rect 6193 7044 6249 7100
rect 6249 7044 6253 7100
rect 6189 7040 6253 7044
rect 10946 7100 11010 7104
rect 10946 7044 10950 7100
rect 10950 7044 11006 7100
rect 11006 7044 11010 7100
rect 10946 7040 11010 7044
rect 11026 7100 11090 7104
rect 11026 7044 11030 7100
rect 11030 7044 11086 7100
rect 11086 7044 11090 7100
rect 11026 7040 11090 7044
rect 11106 7100 11170 7104
rect 11106 7044 11110 7100
rect 11110 7044 11166 7100
rect 11166 7044 11170 7100
rect 11106 7040 11170 7044
rect 11186 7100 11250 7104
rect 11186 7044 11190 7100
rect 11190 7044 11246 7100
rect 11246 7044 11250 7100
rect 11186 7040 11250 7044
rect 3450 6556 3514 6560
rect 3450 6500 3454 6556
rect 3454 6500 3510 6556
rect 3510 6500 3514 6556
rect 3450 6496 3514 6500
rect 3530 6556 3594 6560
rect 3530 6500 3534 6556
rect 3534 6500 3590 6556
rect 3590 6500 3594 6556
rect 3530 6496 3594 6500
rect 3610 6556 3674 6560
rect 3610 6500 3614 6556
rect 3614 6500 3670 6556
rect 3670 6500 3674 6556
rect 3610 6496 3674 6500
rect 3690 6556 3754 6560
rect 3690 6500 3694 6556
rect 3694 6500 3750 6556
rect 3750 6500 3754 6556
rect 3690 6496 3754 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 13445 6556 13509 6560
rect 13445 6500 13449 6556
rect 13449 6500 13505 6556
rect 13505 6500 13509 6556
rect 13445 6496 13509 6500
rect 13525 6556 13589 6560
rect 13525 6500 13529 6556
rect 13529 6500 13585 6556
rect 13585 6500 13589 6556
rect 13525 6496 13589 6500
rect 13605 6556 13669 6560
rect 13605 6500 13609 6556
rect 13609 6500 13665 6556
rect 13665 6500 13669 6556
rect 13605 6496 13669 6500
rect 13685 6556 13749 6560
rect 13685 6500 13689 6556
rect 13689 6500 13745 6556
rect 13745 6500 13749 6556
rect 13685 6496 13749 6500
rect 5949 6012 6013 6016
rect 5949 5956 5953 6012
rect 5953 5956 6009 6012
rect 6009 5956 6013 6012
rect 5949 5952 6013 5956
rect 6029 6012 6093 6016
rect 6029 5956 6033 6012
rect 6033 5956 6089 6012
rect 6089 5956 6093 6012
rect 6029 5952 6093 5956
rect 6109 6012 6173 6016
rect 6109 5956 6113 6012
rect 6113 5956 6169 6012
rect 6169 5956 6173 6012
rect 6109 5952 6173 5956
rect 6189 6012 6253 6016
rect 6189 5956 6193 6012
rect 6193 5956 6249 6012
rect 6249 5956 6253 6012
rect 6189 5952 6253 5956
rect 10946 6012 11010 6016
rect 10946 5956 10950 6012
rect 10950 5956 11006 6012
rect 11006 5956 11010 6012
rect 10946 5952 11010 5956
rect 11026 6012 11090 6016
rect 11026 5956 11030 6012
rect 11030 5956 11086 6012
rect 11086 5956 11090 6012
rect 11026 5952 11090 5956
rect 11106 6012 11170 6016
rect 11106 5956 11110 6012
rect 11110 5956 11166 6012
rect 11166 5956 11170 6012
rect 11106 5952 11170 5956
rect 11186 6012 11250 6016
rect 11186 5956 11190 6012
rect 11190 5956 11246 6012
rect 11246 5956 11250 6012
rect 11186 5952 11250 5956
rect 3450 5468 3514 5472
rect 3450 5412 3454 5468
rect 3454 5412 3510 5468
rect 3510 5412 3514 5468
rect 3450 5408 3514 5412
rect 3530 5468 3594 5472
rect 3530 5412 3534 5468
rect 3534 5412 3590 5468
rect 3590 5412 3594 5468
rect 3530 5408 3594 5412
rect 3610 5468 3674 5472
rect 3610 5412 3614 5468
rect 3614 5412 3670 5468
rect 3670 5412 3674 5468
rect 3610 5408 3674 5412
rect 3690 5468 3754 5472
rect 3690 5412 3694 5468
rect 3694 5412 3750 5468
rect 3750 5412 3754 5468
rect 3690 5408 3754 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 13445 5468 13509 5472
rect 13445 5412 13449 5468
rect 13449 5412 13505 5468
rect 13505 5412 13509 5468
rect 13445 5408 13509 5412
rect 13525 5468 13589 5472
rect 13525 5412 13529 5468
rect 13529 5412 13585 5468
rect 13585 5412 13589 5468
rect 13525 5408 13589 5412
rect 13605 5468 13669 5472
rect 13605 5412 13609 5468
rect 13609 5412 13665 5468
rect 13665 5412 13669 5468
rect 13605 5408 13669 5412
rect 13685 5468 13749 5472
rect 13685 5412 13689 5468
rect 13689 5412 13745 5468
rect 13745 5412 13749 5468
rect 13685 5408 13749 5412
rect 5949 4924 6013 4928
rect 5949 4868 5953 4924
rect 5953 4868 6009 4924
rect 6009 4868 6013 4924
rect 5949 4864 6013 4868
rect 6029 4924 6093 4928
rect 6029 4868 6033 4924
rect 6033 4868 6089 4924
rect 6089 4868 6093 4924
rect 6029 4864 6093 4868
rect 6109 4924 6173 4928
rect 6109 4868 6113 4924
rect 6113 4868 6169 4924
rect 6169 4868 6173 4924
rect 6109 4864 6173 4868
rect 6189 4924 6253 4928
rect 6189 4868 6193 4924
rect 6193 4868 6249 4924
rect 6249 4868 6253 4924
rect 6189 4864 6253 4868
rect 10946 4924 11010 4928
rect 10946 4868 10950 4924
rect 10950 4868 11006 4924
rect 11006 4868 11010 4924
rect 10946 4864 11010 4868
rect 11026 4924 11090 4928
rect 11026 4868 11030 4924
rect 11030 4868 11086 4924
rect 11086 4868 11090 4924
rect 11026 4864 11090 4868
rect 11106 4924 11170 4928
rect 11106 4868 11110 4924
rect 11110 4868 11166 4924
rect 11166 4868 11170 4924
rect 11106 4864 11170 4868
rect 11186 4924 11250 4928
rect 11186 4868 11190 4924
rect 11190 4868 11246 4924
rect 11246 4868 11250 4924
rect 11186 4864 11250 4868
rect 3450 4380 3514 4384
rect 3450 4324 3454 4380
rect 3454 4324 3510 4380
rect 3510 4324 3514 4380
rect 3450 4320 3514 4324
rect 3530 4380 3594 4384
rect 3530 4324 3534 4380
rect 3534 4324 3590 4380
rect 3590 4324 3594 4380
rect 3530 4320 3594 4324
rect 3610 4380 3674 4384
rect 3610 4324 3614 4380
rect 3614 4324 3670 4380
rect 3670 4324 3674 4380
rect 3610 4320 3674 4324
rect 3690 4380 3754 4384
rect 3690 4324 3694 4380
rect 3694 4324 3750 4380
rect 3750 4324 3754 4380
rect 3690 4320 3754 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 13445 4380 13509 4384
rect 13445 4324 13449 4380
rect 13449 4324 13505 4380
rect 13505 4324 13509 4380
rect 13445 4320 13509 4324
rect 13525 4380 13589 4384
rect 13525 4324 13529 4380
rect 13529 4324 13585 4380
rect 13585 4324 13589 4380
rect 13525 4320 13589 4324
rect 13605 4380 13669 4384
rect 13605 4324 13609 4380
rect 13609 4324 13665 4380
rect 13665 4324 13669 4380
rect 13605 4320 13669 4324
rect 13685 4380 13749 4384
rect 13685 4324 13689 4380
rect 13689 4324 13745 4380
rect 13745 4324 13749 4380
rect 13685 4320 13749 4324
rect 5949 3836 6013 3840
rect 5949 3780 5953 3836
rect 5953 3780 6009 3836
rect 6009 3780 6013 3836
rect 5949 3776 6013 3780
rect 6029 3836 6093 3840
rect 6029 3780 6033 3836
rect 6033 3780 6089 3836
rect 6089 3780 6093 3836
rect 6029 3776 6093 3780
rect 6109 3836 6173 3840
rect 6109 3780 6113 3836
rect 6113 3780 6169 3836
rect 6169 3780 6173 3836
rect 6109 3776 6173 3780
rect 6189 3836 6253 3840
rect 6189 3780 6193 3836
rect 6193 3780 6249 3836
rect 6249 3780 6253 3836
rect 6189 3776 6253 3780
rect 10946 3836 11010 3840
rect 10946 3780 10950 3836
rect 10950 3780 11006 3836
rect 11006 3780 11010 3836
rect 10946 3776 11010 3780
rect 11026 3836 11090 3840
rect 11026 3780 11030 3836
rect 11030 3780 11086 3836
rect 11086 3780 11090 3836
rect 11026 3776 11090 3780
rect 11106 3836 11170 3840
rect 11106 3780 11110 3836
rect 11110 3780 11166 3836
rect 11166 3780 11170 3836
rect 11106 3776 11170 3780
rect 11186 3836 11250 3840
rect 11186 3780 11190 3836
rect 11190 3780 11246 3836
rect 11246 3780 11250 3836
rect 11186 3776 11250 3780
rect 3450 3292 3514 3296
rect 3450 3236 3454 3292
rect 3454 3236 3510 3292
rect 3510 3236 3514 3292
rect 3450 3232 3514 3236
rect 3530 3292 3594 3296
rect 3530 3236 3534 3292
rect 3534 3236 3590 3292
rect 3590 3236 3594 3292
rect 3530 3232 3594 3236
rect 3610 3292 3674 3296
rect 3610 3236 3614 3292
rect 3614 3236 3670 3292
rect 3670 3236 3674 3292
rect 3610 3232 3674 3236
rect 3690 3292 3754 3296
rect 3690 3236 3694 3292
rect 3694 3236 3750 3292
rect 3750 3236 3754 3292
rect 3690 3232 3754 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 13445 3292 13509 3296
rect 13445 3236 13449 3292
rect 13449 3236 13505 3292
rect 13505 3236 13509 3292
rect 13445 3232 13509 3236
rect 13525 3292 13589 3296
rect 13525 3236 13529 3292
rect 13529 3236 13585 3292
rect 13585 3236 13589 3292
rect 13525 3232 13589 3236
rect 13605 3292 13669 3296
rect 13605 3236 13609 3292
rect 13609 3236 13665 3292
rect 13665 3236 13669 3292
rect 13605 3232 13669 3236
rect 13685 3292 13749 3296
rect 13685 3236 13689 3292
rect 13689 3236 13745 3292
rect 13745 3236 13749 3292
rect 13685 3232 13749 3236
rect 5949 2748 6013 2752
rect 5949 2692 5953 2748
rect 5953 2692 6009 2748
rect 6009 2692 6013 2748
rect 5949 2688 6013 2692
rect 6029 2748 6093 2752
rect 6029 2692 6033 2748
rect 6033 2692 6089 2748
rect 6089 2692 6093 2748
rect 6029 2688 6093 2692
rect 6109 2748 6173 2752
rect 6109 2692 6113 2748
rect 6113 2692 6169 2748
rect 6169 2692 6173 2748
rect 6109 2688 6173 2692
rect 6189 2748 6253 2752
rect 6189 2692 6193 2748
rect 6193 2692 6249 2748
rect 6249 2692 6253 2748
rect 6189 2688 6253 2692
rect 10946 2748 11010 2752
rect 10946 2692 10950 2748
rect 10950 2692 11006 2748
rect 11006 2692 11010 2748
rect 10946 2688 11010 2692
rect 11026 2748 11090 2752
rect 11026 2692 11030 2748
rect 11030 2692 11086 2748
rect 11086 2692 11090 2748
rect 11026 2688 11090 2692
rect 11106 2748 11170 2752
rect 11106 2692 11110 2748
rect 11110 2692 11166 2748
rect 11166 2692 11170 2748
rect 11106 2688 11170 2692
rect 11186 2748 11250 2752
rect 11186 2692 11190 2748
rect 11190 2692 11246 2748
rect 11246 2692 11250 2748
rect 11186 2688 11250 2692
rect 3450 2204 3514 2208
rect 3450 2148 3454 2204
rect 3454 2148 3510 2204
rect 3510 2148 3514 2204
rect 3450 2144 3514 2148
rect 3530 2204 3594 2208
rect 3530 2148 3534 2204
rect 3534 2148 3590 2204
rect 3590 2148 3594 2204
rect 3530 2144 3594 2148
rect 3610 2204 3674 2208
rect 3610 2148 3614 2204
rect 3614 2148 3670 2204
rect 3670 2148 3674 2204
rect 3610 2144 3674 2148
rect 3690 2204 3754 2208
rect 3690 2148 3694 2204
rect 3694 2148 3750 2204
rect 3750 2148 3754 2204
rect 3690 2144 3754 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 13445 2204 13509 2208
rect 13445 2148 13449 2204
rect 13449 2148 13505 2204
rect 13505 2148 13509 2204
rect 13445 2144 13509 2148
rect 13525 2204 13589 2208
rect 13525 2148 13529 2204
rect 13529 2148 13585 2204
rect 13585 2148 13589 2204
rect 13525 2144 13589 2148
rect 13605 2204 13669 2208
rect 13605 2148 13609 2204
rect 13609 2148 13665 2204
rect 13665 2148 13669 2204
rect 13605 2144 13669 2148
rect 13685 2204 13749 2208
rect 13685 2148 13689 2204
rect 13689 2148 13745 2204
rect 13745 2148 13749 2204
rect 13685 2144 13749 2148
rect 9444 852 9508 916
rect 10364 852 10428 916
<< metal4 >>
rect 10363 19140 10429 19141
rect 10363 19076 10364 19140
rect 10428 19076 10429 19140
rect 10363 19075 10429 19076
rect 3442 17440 3763 17456
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3763 17440
rect 3442 16352 3763 17376
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3763 16352
rect 3442 15264 3763 16288
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3763 15264
rect 3442 14176 3763 15200
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3763 14176
rect 3442 13088 3763 14112
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3763 13088
rect 3442 12000 3763 13024
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3763 12000
rect 3442 10912 3763 11936
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3763 10912
rect 3442 9824 3763 10848
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3763 9824
rect 3442 8736 3763 9760
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3763 8736
rect 3442 7648 3763 8672
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3763 7648
rect 3442 6560 3763 7584
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3763 6560
rect 3442 5472 3763 6496
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3763 5472
rect 3442 4384 3763 5408
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3763 4384
rect 3442 3296 3763 4320
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3763 3296
rect 3442 2208 3763 3232
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3763 2208
rect 3442 2128 3763 2144
rect 5941 16896 6261 17456
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 15808 6261 16832
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 14720 6261 15744
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 13632 6261 14656
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 12544 6261 13568
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 11456 6261 12480
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 10368 6261 11392
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 9280 6261 10304
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 8192 6261 9216
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 7104 6261 8128
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 6016 6261 7040
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 4928 6261 5952
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 3840 6261 4864
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 2752 6261 3776
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2128 6261 2688
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 10366 10029 10426 19075
rect 10938 16896 11259 17456
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11259 16896
rect 10938 15808 11259 16832
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11259 15808
rect 10938 14720 11259 15744
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11259 14720
rect 10938 13632 11259 14656
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11259 13632
rect 10938 12544 11259 13568
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11259 12544
rect 10938 11456 11259 12480
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11259 11456
rect 10938 10368 11259 11392
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11259 10368
rect 10363 10028 10429 10029
rect 10363 9964 10364 10028
rect 10428 9964 10429 10028
rect 10363 9963 10429 9964
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 10363 9620 10429 9621
rect 10363 9556 10364 9620
rect 10428 9556 10429 9620
rect 10363 9555 10429 9556
rect 9443 9484 9509 9485
rect 9443 9420 9444 9484
rect 9508 9420 9509 9484
rect 9443 9419 9509 9420
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 9446 917 9506 9419
rect 10366 917 10426 9555
rect 10938 9280 11259 10304
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11259 9280
rect 10938 8192 11259 9216
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11259 8192
rect 10938 7104 11259 8128
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11259 7104
rect 10938 6016 11259 7040
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11259 6016
rect 10938 4928 11259 5952
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11259 4928
rect 10938 3840 11259 4864
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11259 3840
rect 10938 2752 11259 3776
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11259 2752
rect 10938 2128 11259 2688
rect 13437 17440 13757 17456
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 16352 13757 17376
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 15264 13757 16288
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 14176 13757 15200
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 13088 13757 14112
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 12000 13757 13024
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 10912 13757 11936
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 9824 13757 10848
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 8736 13757 9760
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 7648 13757 8672
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 6560 13757 7584
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 5472 13757 6496
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 4384 13757 5408
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 3296 13757 4320
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 13437 2208 13757 3232
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2128 13757 2144
rect 9443 916 9509 917
rect 9443 852 9444 916
rect 9508 852 9509 916
rect 9443 851 9509 852
rect 10363 916 10429 917
rect 10363 852 10364 916
rect 10428 852 10429 916
rect 10363 851 10429 852
use sky130_fd_sc_hd__decap_12  FILLER_1_15 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608910539
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608910539
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1608910539
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608910539
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1608910539
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1608910539
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1608910539
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1608910539
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608910539
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608910539
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608910539
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608910539
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608910539
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608910539
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1608910539
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1608910539
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1608910539
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15640 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608910539
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608910539
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608910539
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1608910539
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1608910539
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1608910539
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1608910539
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1608910539
transform 1 0 6716 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1608910539
transform 1 0 6440 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_46
timestamp 1608910539
transform 1 0 5336 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_65
timestamp 1608910539
transform 1 0 7084 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1608910539
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1608910539
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1608910539
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1608910539
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_76
timestamp 1608910539
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1608910539
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1608910539
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_80
timestamp 1608910539
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1608910539
transform 1 0 8648 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1608910539
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1608910539
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _36_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_95
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1608910539
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1608910539
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1608910539
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1608910539
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp 1608910539
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1608910539
transform 1 0 12236 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_116
timestamp 1608910539
transform 1 0 11776 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_113
timestamp 1608910539
transform 1 0 11500 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_107
timestamp 1608910539
transform 1 0 10948 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608910539
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1608910539
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1608910539
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1608910539
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1608910539
transform 1 0 15640 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_39
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1608910539
transform 1 0 4784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_50
timestamp 1608910539
transform 1 0 5704 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__02__A
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608910539
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608910539
transform 1 0 5152 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1608910539
transform 1 0 6164 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1608910539
transform 1 0 5796 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1608910539
transform 1 0 8648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1608910539
transform 1 0 8280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1608910539
transform 1 0 7912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1608910539
transform 1 0 7544 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1608910539
transform 1 0 7176 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp 1608910539
transform 1 0 9936 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_91
timestamp 1608910539
transform 1 0 9476 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_86
timestamp 1608910539
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1608910539
transform 1 0 10396 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1608910539
transform 1 0 10028 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1608910539
transform 1 0 9568 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1608910539
transform 1 0 9108 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608910539
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_114
timestamp 1608910539
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_105
timestamp 1608910539
transform 1 0 10764 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1608910539
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608910539
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1608910539
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1608910539
transform 1 0 10856 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1608910539
transform 1 0 14076 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608910539
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1608910539
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1608910539
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608910539
transform 1 0 13156 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1608910539
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_153
timestamp 1608910539
transform 1 0 15180 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1608910539
transform 1 0 4784 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1608910539
transform 1 0 4416 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_50
timestamp 1608910539
transform 1 0 5704 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1608910539
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1608910539
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1608910539
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_58
timestamp 1608910539
transform 1 0 6440 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1608910539
transform 1 0 6532 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1608910539
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_65
timestamp 1608910539
transform 1 0 7084 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_63
timestamp 1608910539
transform 1 0 6900 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1608910539
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1608910539
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1608910539
transform 1 0 6900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1608910539
transform 1 0 7728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1608910539
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1608910539
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1608910539
transform 1 0 8096 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1608910539
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1608910539
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1608910539
transform 1 0 8188 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1608910539
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1608910539
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1608910539
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1608910539
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1608910539
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608910539
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608910539
transform 1 0 10028 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1608910539
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_111
timestamp 1608910539
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1608910539
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1608910539
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1608910539
transform 1 0 10764 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608910539
transform 1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1608910539
transform 1 0 11960 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608910539
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608910539
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608910539
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1608910539
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608910539
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1608910539
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1608910539
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1608910539
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1608910539
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608910539
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608910539
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1608910539
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608910539
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1608910539
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1608910539
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1608910539
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1608910539
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1608910539
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1608910539
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_30
timestamp 1608910539
transform 1 0 3864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_23
timestamp 1608910539
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3312 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1608910539
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1608910539
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1608910539
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1608910539
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1608910539
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1608910539
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1608910539
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1608910539
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608910539
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608910539
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608910539
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608910539
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1608910539
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1608910539
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1608910539
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1608910539
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1608910539
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1608910539
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608910539
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608910539
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608910539
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608910539
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1608910539
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1608910539
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1608910539
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1608910539
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1608910539
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1608910539
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_56
timestamp 1608910539
transform 1 0 6256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608910539
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_117
timestamp 1608910539
transform 1 0 11868 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1608910539
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_137
timestamp 1608910539
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 13524 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1608910539
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1608910539
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_16
timestamp 1608910539
transform 1 0 2576 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_17
timestamp 1608910539
transform 1 0 2668 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_5
timestamp 1608910539
transform 1 0 1564 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1608910539
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_41
timestamp 1608910539
transform 1 0 4876 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_29
timestamp 1608910539
transform 1 0 3772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_56
timestamp 1608910539
transform 1 0 6256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608910539
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1608910539
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8096 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7360 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1608910539
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1608910539
transform 1 0 9936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8924 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_118
timestamp 1608910539
transform 1 0 11960 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_106
timestamp 1608910539
transform 1 0 10856 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608910539
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_108
timestamp 1608910539
transform 1 0 11040 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_142
timestamp 1608910539
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_130
timestamp 1608910539
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1608910539
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1608910539
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1608910539
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1608910539
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1608910539
transform 1 0 2484 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_41
timestamp 1608910539
transform 1 0 4876 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_22
timestamp 1608910539
transform 1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1608910539
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1608910539
transform 1 0 3680 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_15_53
timestamp 1608910539
transform 1 0 5980 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7636 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1608910539
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _01_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 10764 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1608910539
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1608910539
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608910539
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608910539
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_56
timestamp 1608910539
transform 1 0 6256 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6624 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_69
timestamp 1608910539
transform 1 0 7452 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7820 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_100
timestamp 1608910539
transform 1 0 10304 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1608910539
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_124
timestamp 1608910539
transform 1 0 12512 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_112
timestamp 1608910539
transform 1 0 11408 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_136
timestamp 1608910539
transform 1 0 13616 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1608910539
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608910539
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1608910539
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608910539
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1608910539
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1608910539
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608910539
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7360 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_96
timestamp 1608910539
transform 1 0 9936 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_84
timestamp 1608910539
transform 1 0 8832 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608910539
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_108
timestamp 1608910539
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1608910539
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1608910539
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608910539
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608910539
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1608910539
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_44
timestamp 1608910539
transform 1 0 5152 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6072 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_18_74
timestamp 1608910539
transform 1 0 7912 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_86
timestamp 1608910539
transform 1 0 9016 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1608910539
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1608910539
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1608910539
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1608910539
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1608910539
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1608910539
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1608910539
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_40
timestamp 1608910539
transform 1 0 4784 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1608910539
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1608910539
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608910539
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608910539
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1608910539
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1608910539
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608910539
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608910539
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1608910539
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp 1608910539
transform 1 0 14076 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1608910539
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1608910539
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1608910539
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608910539
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_27
timestamp 1608910539
transform 1 0 3588 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4324 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608910539
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1608910539
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1608910539
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1608910539
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1608910539
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1608910539
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608910539
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_56
timestamp 1608910539
transform 1 0 6256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_73
timestamp 1608910539
transform 1 0 7820 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_64
timestamp 1608910539
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1608910539
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1608910539
transform 1 0 7268 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1608910539
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1608910539
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1608910539
transform 1 0 8924 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1608910539
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1608910539
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1608910539
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_135
timestamp 1608910539
transform 1 0 13524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1608910539
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1608910539
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608910539
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_36
timestamp 1608910539
transform 1 0 4416 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp 1608910539
transform 1 0 3588 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608910539
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608910539
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608910539
transform 1 0 4508 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608910539
transform 1 0 3864 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608910539
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_52
timestamp 1608910539
transform 1 0 5888 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_43
timestamp 1608910539
transform 1 0 5060 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__03__A
timestamp 1608910539
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1608910539
transform 1 0 5336 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1608910539
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1608910539
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1608910539
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1608910539
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1608910539
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1608910539
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608910539
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1608910539
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1608910539
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1608910539
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1608910539
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1608910539
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1608910539
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1608910539
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1608910539
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1608910539
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1608910539
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1608910539
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1608910539
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1608910539
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1608910539
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1608910539
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1608910539
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1608910539
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1608910539
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1608910539
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608910539
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1608910539
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1608910539
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608910539
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1608910539
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1608910539
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1608910539
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1608910539
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_75
timestamp 1608910539
transform 1 0 8004 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_63
timestamp 1608910539
transform 1 0 6900 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1608910539
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1608910539
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1608910539
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_87
timestamp 1608910539
transform 1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1608910539
transform 1 0 12604 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_118
timestamp 1608910539
transform 1 0 11960 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1608910539
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1608910539
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1608910539
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1608910539
transform 1 0 13708 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1608910539
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1608910539
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_156
timestamp 1608910539
transform 1 0 15456 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_149
timestamp 1608910539
transform 1 0 14812 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1608910539
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 16400 12384 17200 12504 6 ccff_tail
port 2 nsew signal tristate
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[0]
port 3 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_in[10]
port 4 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[11]
port 5 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_in[12]
port 6 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_in[13]
port 7 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_in[14]
port 8 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_in[15]
port 9 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[16]
port 10 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_in[17]
port 11 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[18]
port 12 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_in[19]
port 13 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[1]
port 14 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[2]
port 15 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[3]
port 16 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[4]
port 17 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[5]
port 18 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[6]
port 19 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[7]
port 20 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[8]
port 21 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[9]
port 22 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 23 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_out[10]
port 24 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[11]
port 25 nsew signal tristate
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_out[12]
port 26 nsew signal tristate
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_out[13]
port 27 nsew signal tristate
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[14]
port 28 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[15]
port 29 nsew signal tristate
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_out[16]
port 30 nsew signal tristate
rlabel metal2 s 7470 0 7526 800 6 chany_bottom_out[17]
port 31 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_out[18]
port 32 nsew signal tristate
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_out[19]
port 33 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 34 nsew signal tristate
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 35 nsew signal tristate
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_out[3]
port 36 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 37 nsew signal tristate
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[5]
port 38 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[6]
port 39 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[7]
port 40 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_out[8]
port 41 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_out[9]
port 42 nsew signal tristate
rlabel metal2 s 8942 19200 8998 20000 6 chany_top_in[0]
port 43 nsew signal input
rlabel metal2 s 13174 19200 13230 20000 6 chany_top_in[10]
port 44 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[11]
port 45 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[12]
port 46 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[13]
port 47 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 chany_top_in[14]
port 48 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[15]
port 49 nsew signal input
rlabel metal2 s 15658 19200 15714 20000 6 chany_top_in[16]
port 50 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[17]
port 51 nsew signal input
rlabel metal2 s 16486 19200 16542 20000 6 chany_top_in[18]
port 52 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 53 nsew signal input
rlabel metal2 s 9402 19200 9458 20000 6 chany_top_in[1]
port 54 nsew signal input
rlabel metal2 s 9770 19200 9826 20000 6 chany_top_in[2]
port 55 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[3]
port 56 nsew signal input
rlabel metal2 s 10690 19200 10746 20000 6 chany_top_in[4]
port 57 nsew signal input
rlabel metal2 s 11058 19200 11114 20000 6 chany_top_in[5]
port 58 nsew signal input
rlabel metal2 s 11518 19200 11574 20000 6 chany_top_in[6]
port 59 nsew signal input
rlabel metal2 s 11886 19200 11942 20000 6 chany_top_in[7]
port 60 nsew signal input
rlabel metal2 s 12346 19200 12402 20000 6 chany_top_in[8]
port 61 nsew signal input
rlabel metal2 s 12714 19200 12770 20000 6 chany_top_in[9]
port 62 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 63 nsew signal tristate
rlabel metal2 s 4802 19200 4858 20000 6 chany_top_out[10]
port 64 nsew signal tristate
rlabel metal2 s 5170 19200 5226 20000 6 chany_top_out[11]
port 65 nsew signal tristate
rlabel metal2 s 5630 19200 5686 20000 6 chany_top_out[12]
port 66 nsew signal tristate
rlabel metal2 s 5998 19200 6054 20000 6 chany_top_out[13]
port 67 nsew signal tristate
rlabel metal2 s 6458 19200 6514 20000 6 chany_top_out[14]
port 68 nsew signal tristate
rlabel metal2 s 6826 19200 6882 20000 6 chany_top_out[15]
port 69 nsew signal tristate
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[16]
port 70 nsew signal tristate
rlabel metal2 s 7746 19200 7802 20000 6 chany_top_out[17]
port 71 nsew signal tristate
rlabel metal2 s 8114 19200 8170 20000 6 chany_top_out[18]
port 72 nsew signal tristate
rlabel metal2 s 8574 19200 8630 20000 6 chany_top_out[19]
port 73 nsew signal tristate
rlabel metal2 s 1030 19200 1086 20000 6 chany_top_out[1]
port 74 nsew signal tristate
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 75 nsew signal tristate
rlabel metal2 s 1858 19200 1914 20000 6 chany_top_out[3]
port 76 nsew signal tristate
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 77 nsew signal tristate
rlabel metal2 s 2686 19200 2742 20000 6 chany_top_out[5]
port 78 nsew signal tristate
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 79 nsew signal tristate
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[7]
port 80 nsew signal tristate
rlabel metal2 s 3974 19200 4030 20000 6 chany_top_out[8]
port 81 nsew signal tristate
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[9]
port 82 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 83 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 84 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 85 nsew signal tristate
rlabel metal3 s 0 4904 800 5024 6 left_grid_pin_0_
port 86 nsew signal tristate
rlabel metal3 s 16400 7352 17200 7472 6 prog_clk_0_E_in
port 87 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 right_width_0_height_0__pin_0_
port 88 nsew signal input
rlabel metal3 s 16400 2456 17200 2576 6 right_width_0_height_0__pin_1_lower
port 89 nsew signal tristate
rlabel metal3 s 16400 17416 17200 17536 6 right_width_0_height_0__pin_1_upper
port 90 nsew signal tristate
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 91 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 92 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 94 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 95 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
