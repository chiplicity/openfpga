magic
tech sky130A
magscale 1 2
timestamp 1606227864
<< locali >>
rect 8309 18683 8343 18853
rect 13921 18071 13955 18173
rect 7389 17595 7423 17697
rect 7481 17595 7515 17765
rect 14381 12767 14415 12937
rect 9965 10455 9999 10557
rect 6469 7803 6503 8041
<< viali >>
rect 1961 20009 1995 20043
rect 4537 20009 4571 20043
rect 5365 20009 5399 20043
rect 5825 20009 5859 20043
rect 9137 20009 9171 20043
rect 13185 20009 13219 20043
rect 15669 20009 15703 20043
rect 16773 20009 16807 20043
rect 17325 20009 17359 20043
rect 18521 20009 18555 20043
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 3525 19873 3559 19907
rect 4445 19873 4479 19907
rect 5733 19873 5767 19907
rect 9045 19873 9079 19907
rect 11060 19873 11094 19907
rect 13001 19873 13035 19907
rect 13829 19873 13863 19907
rect 14565 19873 14599 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 16589 19873 16623 19907
rect 17141 19873 17175 19907
rect 18337 19873 18371 19907
rect 4721 19805 4755 19839
rect 6009 19805 6043 19839
rect 9321 19805 9355 19839
rect 10793 19805 10827 19839
rect 14105 19805 14139 19839
rect 14841 19805 14875 19839
rect 2513 19737 2547 19771
rect 16221 19737 16255 19771
rect 4077 19669 4111 19703
rect 8677 19669 8711 19703
rect 12173 19669 12207 19703
rect 6469 19465 6503 19499
rect 14657 19465 14691 19499
rect 2329 19329 2363 19363
rect 14197 19329 14231 19363
rect 15209 19329 15243 19363
rect 1593 19261 1627 19295
rect 2145 19261 2179 19295
rect 3065 19261 3099 19295
rect 5089 19261 5123 19295
rect 6837 19261 6871 19295
rect 9229 19261 9263 19295
rect 11529 19261 11563 19295
rect 12909 19261 12943 19295
rect 14105 19261 14139 19295
rect 16129 19261 16163 19295
rect 16865 19261 16899 19295
rect 17417 19261 17451 19295
rect 18061 19261 18095 19295
rect 18613 19261 18647 19295
rect 19165 19261 19199 19295
rect 3332 19193 3366 19227
rect 5356 19193 5390 19227
rect 7082 19193 7116 19227
rect 9496 19193 9530 19227
rect 15025 19193 15059 19227
rect 16405 19193 16439 19227
rect 1777 19125 1811 19159
rect 4445 19125 4479 19159
rect 8217 19125 8251 19159
rect 8769 19125 8803 19159
rect 10609 19125 10643 19159
rect 11713 19125 11747 19159
rect 13093 19125 13127 19159
rect 13645 19125 13679 19159
rect 14013 19125 14047 19159
rect 15117 19125 15151 19159
rect 17049 19125 17083 19159
rect 17601 19125 17635 19159
rect 18245 19125 18279 19159
rect 18797 19125 18831 19159
rect 19349 19125 19383 19159
rect 2789 18921 2823 18955
rect 3249 18921 3283 18955
rect 4077 18921 4111 18955
rect 4537 18921 4571 18955
rect 8769 18921 8803 18955
rect 8861 18921 8895 18955
rect 2329 18853 2363 18887
rect 7941 18853 7975 18887
rect 8309 18853 8343 18887
rect 9934 18853 9968 18887
rect 12081 18853 12115 18887
rect 12817 18853 12851 18887
rect 15761 18853 15795 18887
rect 17325 18853 17359 18887
rect 18061 18853 18095 18887
rect 18797 18853 18831 18887
rect 2053 18785 2087 18819
rect 3157 18785 3191 18819
rect 4445 18785 4479 18819
rect 5457 18785 5491 18819
rect 6101 18785 6135 18819
rect 7665 18785 7699 18819
rect 3341 18717 3375 18751
rect 4629 18717 4663 18751
rect 5549 18717 5583 18751
rect 5733 18717 5767 18751
rect 9689 18785 9723 18819
rect 11805 18785 11839 18819
rect 12541 18785 12575 18819
rect 13820 18785 13854 18819
rect 15485 18785 15519 18819
rect 16313 18785 16347 18819
rect 16589 18785 16623 18819
rect 17049 18785 17083 18819
rect 17785 18785 17819 18819
rect 18521 18785 18555 18819
rect 9045 18717 9079 18751
rect 13553 18717 13587 18751
rect 8309 18649 8343 18683
rect 8401 18649 8435 18683
rect 5089 18581 5123 18615
rect 11069 18581 11103 18615
rect 14933 18581 14967 18615
rect 14289 18377 14323 18411
rect 6469 18309 6503 18343
rect 2145 18241 2179 18275
rect 7389 18241 7423 18275
rect 9505 18241 9539 18275
rect 9689 18241 9723 18275
rect 15209 18241 15243 18275
rect 15669 18241 15703 18275
rect 16589 18241 16623 18275
rect 18245 18241 18279 18275
rect 1409 18173 1443 18207
rect 1961 18173 1995 18207
rect 2697 18173 2731 18207
rect 2964 18173 2998 18207
rect 5089 18173 5123 18207
rect 7656 18173 7690 18207
rect 10333 18173 10367 18207
rect 12449 18173 12483 18207
rect 13921 18173 13955 18207
rect 14105 18173 14139 18207
rect 15025 18173 15059 18207
rect 16313 18173 16347 18207
rect 18061 18173 18095 18207
rect 5356 18105 5390 18139
rect 10600 18105 10634 18139
rect 12716 18105 12750 18139
rect 15117 18105 15151 18139
rect 1593 18037 1627 18071
rect 4077 18037 4111 18071
rect 8769 18037 8803 18071
rect 9045 18037 9079 18071
rect 9413 18037 9447 18071
rect 11713 18037 11747 18071
rect 13829 18037 13863 18071
rect 13921 18037 13955 18071
rect 14657 18037 14691 18071
rect 1961 17833 1995 17867
rect 2513 17833 2547 17867
rect 3065 17833 3099 17867
rect 3433 17833 3467 17867
rect 5641 17833 5675 17867
rect 6101 17833 6135 17867
rect 8033 17833 8067 17867
rect 10425 17833 10459 17867
rect 12449 17833 12483 17867
rect 14197 17833 14231 17867
rect 14565 17833 14599 17867
rect 14657 17833 14691 17867
rect 15301 17833 15335 17867
rect 15669 17833 15703 17867
rect 7481 17765 7515 17799
rect 17202 17765 17236 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2881 17697 2915 17731
rect 6009 17697 6043 17731
rect 6837 17697 6871 17731
rect 7113 17697 7147 17731
rect 7389 17697 7423 17731
rect 6193 17629 6227 17663
rect 7389 17561 7423 17595
rect 7941 17697 7975 17731
rect 8861 17697 8895 17731
rect 10333 17697 10367 17731
rect 12817 17697 12851 17731
rect 8217 17629 8251 17663
rect 9045 17629 9079 17663
rect 10609 17629 10643 17663
rect 10977 17629 11011 17663
rect 12909 17629 12943 17663
rect 13001 17629 13035 17663
rect 14749 17629 14783 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 16957 17629 16991 17663
rect 7481 17561 7515 17595
rect 7573 17561 7607 17595
rect 9965 17493 9999 17527
rect 18337 17493 18371 17527
rect 6193 17289 6227 17323
rect 7665 17289 7699 17323
rect 9965 17289 9999 17323
rect 16497 17289 16531 17323
rect 19073 17289 19107 17323
rect 18061 17221 18095 17255
rect 2329 17153 2363 17187
rect 7941 17153 7975 17187
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 12541 17153 12575 17187
rect 17141 17153 17175 17187
rect 18613 17153 18647 17187
rect 19533 17153 19567 17187
rect 19625 17153 19659 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 2789 17085 2823 17119
rect 3056 17085 3090 17119
rect 4813 17085 4847 17119
rect 7849 17085 7883 17119
rect 8769 17085 8803 17119
rect 10333 17085 10367 17119
rect 12081 17085 12115 17119
rect 14381 17085 14415 17119
rect 14648 17085 14682 17119
rect 18429 17085 18463 17119
rect 5080 17017 5114 17051
rect 9045 17017 9079 17051
rect 12808 17017 12842 17051
rect 16037 17017 16071 17051
rect 16865 17017 16899 17051
rect 17509 17017 17543 17051
rect 19441 17017 19475 17051
rect 1685 16949 1719 16983
rect 4169 16949 4203 16983
rect 11897 16949 11931 16983
rect 13921 16949 13955 16983
rect 15761 16949 15795 16983
rect 16957 16949 16991 16983
rect 18521 16949 18555 16983
rect 1777 16745 1811 16779
rect 4537 16745 4571 16779
rect 4997 16745 5031 16779
rect 5549 16745 5583 16779
rect 6009 16745 6043 16779
rect 11161 16745 11195 16779
rect 12357 16745 12391 16779
rect 17325 16745 17359 16779
rect 4905 16677 4939 16711
rect 6561 16677 6595 16711
rect 7564 16677 7598 16711
rect 18052 16677 18086 16711
rect 1593 16609 1627 16643
rect 2145 16609 2179 16643
rect 5917 16609 5951 16643
rect 7297 16609 7331 16643
rect 9781 16609 9815 16643
rect 10048 16609 10082 16643
rect 12725 16609 12759 16643
rect 15945 16609 15979 16643
rect 16212 16609 16246 16643
rect 17785 16609 17819 16643
rect 2329 16541 2363 16575
rect 5181 16541 5215 16575
rect 6101 16541 6135 16575
rect 12817 16541 12851 16575
rect 13001 16541 13035 16575
rect 8677 16405 8711 16439
rect 19165 16405 19199 16439
rect 1593 16201 1627 16235
rect 2881 16201 2915 16235
rect 6009 16201 6043 16235
rect 10793 16201 10827 16235
rect 13829 16201 13863 16235
rect 15301 16201 15335 16235
rect 15577 16201 15611 16235
rect 2145 16065 2179 16099
rect 4077 16065 4111 16099
rect 11529 16065 11563 16099
rect 11621 16065 11655 16099
rect 14657 16065 14691 16099
rect 16221 16065 16255 16099
rect 1409 15997 1443 16031
rect 1961 15997 1995 16031
rect 2697 15997 2731 16031
rect 3801 15997 3835 16031
rect 4629 15997 4663 16031
rect 6837 15997 6871 16031
rect 9413 15997 9447 16031
rect 9680 15997 9714 16031
rect 12449 15997 12483 16031
rect 15485 15997 15519 16031
rect 4896 15929 4930 15963
rect 7104 15929 7138 15963
rect 11437 15929 11471 15963
rect 12694 15929 12728 15963
rect 14565 15929 14599 15963
rect 16037 15929 16071 15963
rect 3433 15861 3467 15895
rect 3893 15861 3927 15895
rect 6285 15861 6319 15895
rect 8217 15861 8251 15895
rect 8953 15861 8987 15895
rect 11069 15861 11103 15895
rect 14105 15861 14139 15895
rect 14473 15861 14507 15895
rect 15945 15861 15979 15895
rect 1961 15657 1995 15691
rect 6561 15657 6595 15691
rect 6929 15657 6963 15691
rect 7021 15657 7055 15691
rect 7573 15657 7607 15691
rect 8033 15657 8067 15691
rect 9689 15657 9723 15691
rect 10057 15657 10091 15691
rect 10149 15657 10183 15691
rect 11437 15657 11471 15691
rect 12449 15657 12483 15691
rect 12817 15657 12851 15691
rect 17141 15657 17175 15691
rect 2596 15589 2630 15623
rect 7941 15589 7975 15623
rect 13728 15589 13762 15623
rect 18328 15589 18362 15623
rect 1777 15521 1811 15555
rect 5549 15521 5583 15555
rect 11805 15521 11839 15555
rect 13461 15521 13495 15555
rect 15761 15521 15795 15555
rect 16028 15521 16062 15555
rect 2329 15453 2363 15487
rect 4077 15453 4111 15487
rect 4905 15453 4939 15487
rect 7205 15453 7239 15487
rect 8217 15453 8251 15487
rect 10333 15453 10367 15487
rect 11897 15453 11931 15487
rect 12081 15453 12115 15487
rect 12909 15453 12943 15487
rect 13093 15453 13127 15487
rect 18061 15453 18095 15487
rect 3709 15317 3743 15351
rect 5365 15317 5399 15351
rect 14841 15317 14875 15351
rect 19441 15317 19475 15351
rect 2605 15113 2639 15147
rect 6101 15113 6135 15147
rect 7021 15113 7055 15147
rect 9873 15113 9907 15147
rect 13737 15113 13771 15147
rect 15945 15113 15979 15147
rect 10977 15045 11011 15079
rect 13093 15045 13127 15079
rect 2145 14977 2179 15011
rect 3065 14977 3099 15011
rect 3249 14977 3283 15011
rect 8493 14977 8527 15011
rect 11437 14977 11471 15011
rect 11529 14977 11563 15011
rect 12449 14977 12483 15011
rect 14197 14977 14231 15011
rect 14381 14977 14415 15011
rect 16497 14977 16531 15011
rect 18705 14977 18739 15011
rect 1858 14909 1892 14943
rect 2973 14909 3007 14943
rect 4721 14909 4755 14943
rect 7205 14909 7239 14943
rect 11345 14909 11379 14943
rect 13277 14909 13311 14943
rect 18521 14909 18555 14943
rect 4988 14841 5022 14875
rect 8760 14841 8794 14875
rect 16313 14841 16347 14875
rect 16957 14841 16991 14875
rect 18889 14841 18923 14875
rect 14105 14773 14139 14807
rect 16405 14773 16439 14807
rect 18061 14773 18095 14807
rect 18429 14773 18463 14807
rect 1593 14569 1627 14603
rect 5733 14569 5767 14603
rect 9045 14569 9079 14603
rect 14473 14569 14507 14603
rect 16865 14569 16899 14603
rect 2237 14501 2271 14535
rect 6552 14501 6586 14535
rect 10784 14501 10818 14535
rect 17509 14501 17543 14535
rect 18236 14501 18270 14535
rect 1409 14433 1443 14467
rect 1961 14433 1995 14467
rect 4353 14433 4387 14467
rect 4620 14433 4654 14467
rect 8953 14433 8987 14467
rect 12357 14433 12391 14467
rect 13093 14433 13127 14467
rect 13360 14433 13394 14467
rect 15485 14433 15519 14467
rect 15752 14433 15786 14467
rect 6285 14365 6319 14399
rect 8125 14365 8159 14399
rect 9137 14365 9171 14399
rect 10517 14365 10551 14399
rect 12541 14365 12575 14399
rect 17969 14365 18003 14399
rect 7665 14229 7699 14263
rect 8585 14229 8619 14263
rect 11897 14229 11931 14263
rect 19349 14229 19383 14263
rect 4537 14025 4571 14059
rect 9321 14025 9355 14059
rect 12633 14025 12667 14059
rect 15025 14025 15059 14059
rect 17417 14025 17451 14059
rect 18061 14025 18095 14059
rect 5549 13957 5583 13991
rect 6837 13957 6871 13991
rect 12081 13957 12115 13991
rect 1869 13889 1903 13923
rect 2421 13889 2455 13923
rect 4997 13889 5031 13923
rect 5181 13889 5215 13923
rect 6101 13889 6135 13923
rect 7481 13889 7515 13923
rect 7941 13889 7975 13923
rect 10517 13889 10551 13923
rect 11437 13889 11471 13923
rect 11529 13889 11563 13923
rect 13277 13889 13311 13923
rect 15485 13889 15519 13923
rect 15669 13889 15703 13923
rect 18521 13889 18555 13923
rect 18705 13889 18739 13923
rect 1685 13821 1719 13855
rect 2688 13821 2722 13855
rect 6009 13821 6043 13855
rect 7297 13821 7331 13855
rect 8208 13821 8242 13855
rect 10241 13821 10275 13855
rect 12265 13821 12299 13855
rect 16037 13821 16071 13855
rect 4905 13753 4939 13787
rect 7205 13753 7239 13787
rect 16304 13753 16338 13787
rect 18429 13753 18463 13787
rect 3801 13685 3835 13719
rect 5917 13685 5951 13719
rect 10977 13685 11011 13719
rect 11345 13685 11379 13719
rect 13001 13685 13035 13719
rect 13093 13685 13127 13719
rect 15393 13685 15427 13719
rect 1593 13481 1627 13515
rect 2697 13481 2731 13515
rect 3157 13481 3191 13515
rect 4077 13481 4111 13515
rect 4537 13481 4571 13515
rect 5273 13481 5307 13515
rect 5733 13481 5767 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 8493 13481 8527 13515
rect 13921 13481 13955 13515
rect 14565 13481 14599 13515
rect 14657 13481 14691 13515
rect 15761 13481 15795 13515
rect 4445 13413 4479 13447
rect 6552 13413 6586 13447
rect 17960 13413 17994 13447
rect 1409 13345 1443 13379
rect 1961 13345 1995 13379
rect 3065 13345 3099 13379
rect 5641 13345 5675 13379
rect 10149 13345 10183 13379
rect 12808 13345 12842 13379
rect 16129 13345 16163 13379
rect 16773 13345 16807 13379
rect 17693 13345 17727 13379
rect 2145 13277 2179 13311
rect 3341 13277 3375 13311
rect 4629 13277 4663 13311
rect 5917 13277 5951 13311
rect 6285 13277 6319 13311
rect 8677 13277 8711 13311
rect 9689 13277 9723 13311
rect 12541 13277 12575 13311
rect 14841 13277 14875 13311
rect 16221 13277 16255 13311
rect 16405 13277 16439 13311
rect 7665 13141 7699 13175
rect 11437 13141 11471 13175
rect 14197 13141 14231 13175
rect 19073 13141 19107 13175
rect 2513 12937 2547 12971
rect 7573 12937 7607 12971
rect 10701 12937 10735 12971
rect 11529 12937 11563 12971
rect 12449 12937 12483 12971
rect 14381 12937 14415 12971
rect 16681 12937 16715 12971
rect 16957 12937 16991 12971
rect 18061 12937 18095 12971
rect 1961 12869 1995 12903
rect 4629 12869 4663 12903
rect 10609 12869 10643 12903
rect 6193 12801 6227 12835
rect 11161 12801 11195 12835
rect 11345 12801 11379 12835
rect 12081 12801 12115 12835
rect 13001 12801 13035 12835
rect 14105 12801 14139 12835
rect 15301 12801 15335 12835
rect 17509 12801 17543 12835
rect 18705 12801 18739 12835
rect 1777 12733 1811 12767
rect 2329 12733 2363 12767
rect 3249 12733 3283 12767
rect 7757 12733 7791 12767
rect 9229 12733 9263 12767
rect 9496 12733 9530 12767
rect 13921 12733 13955 12767
rect 14381 12733 14415 12767
rect 14657 12733 14691 12767
rect 15568 12733 15602 12767
rect 17417 12733 17451 12767
rect 3516 12665 3550 12699
rect 11069 12665 11103 12699
rect 11989 12665 12023 12699
rect 12817 12665 12851 12699
rect 18429 12665 18463 12699
rect 11897 12597 11931 12631
rect 12909 12597 12943 12631
rect 13461 12597 13495 12631
rect 13829 12597 13863 12631
rect 14473 12597 14507 12631
rect 17325 12597 17359 12631
rect 18521 12597 18555 12631
rect 3525 12393 3559 12427
rect 5641 12393 5675 12427
rect 9137 12393 9171 12427
rect 10057 12393 10091 12427
rect 13645 12393 13679 12427
rect 14933 12393 14967 12427
rect 16681 12393 16715 12427
rect 17601 12393 17635 12427
rect 2329 12325 2363 12359
rect 3065 12325 3099 12359
rect 6184 12325 6218 12359
rect 10149 12325 10183 12359
rect 12256 12325 12290 12359
rect 15568 12325 15602 12359
rect 17969 12325 18003 12359
rect 2053 12257 2087 12291
rect 2789 12257 2823 12291
rect 4528 12257 4562 12291
rect 8013 12257 8047 12291
rect 11989 12257 12023 12291
rect 14013 12257 14047 12291
rect 15117 12257 15151 12291
rect 15301 12257 15335 12291
rect 18061 12257 18095 12291
rect 4261 12189 4295 12223
rect 5917 12189 5951 12223
rect 7757 12189 7791 12223
rect 10333 12189 10367 12223
rect 14105 12189 14139 12223
rect 14197 12189 14231 12223
rect 18245 12189 18279 12223
rect 9689 12121 9723 12155
rect 7297 12053 7331 12087
rect 13369 12053 13403 12087
rect 1593 11849 1627 11883
rect 2881 11849 2915 11883
rect 5181 11849 5215 11883
rect 12449 11849 12483 11883
rect 16957 11849 16991 11883
rect 19993 11849 20027 11883
rect 6377 11713 6411 11747
rect 7389 11713 7423 11747
rect 9781 11713 9815 11747
rect 13093 11713 13127 11747
rect 13461 11713 13495 11747
rect 17601 11713 17635 11747
rect 1409 11645 1443 11679
rect 1961 11645 1995 11679
rect 2237 11645 2271 11679
rect 2697 11645 2731 11679
rect 3801 11645 3835 11679
rect 4068 11645 4102 11679
rect 7205 11645 7239 11679
rect 10048 11645 10082 11679
rect 14381 11645 14415 11679
rect 17417 11645 17451 11679
rect 18613 11645 18647 11679
rect 6101 11577 6135 11611
rect 6193 11577 6227 11611
rect 7656 11577 7690 11611
rect 14626 11577 14660 11611
rect 17325 11577 17359 11611
rect 18061 11577 18095 11611
rect 18880 11577 18914 11611
rect 5733 11509 5767 11543
rect 7021 11509 7055 11543
rect 8769 11509 8803 11543
rect 11161 11509 11195 11543
rect 12817 11509 12851 11543
rect 12909 11509 12943 11543
rect 15761 11509 15795 11543
rect 16037 11509 16071 11543
rect 4537 11305 4571 11339
rect 4905 11305 4939 11339
rect 5549 11305 5583 11339
rect 6837 11305 6871 11339
rect 7297 11305 7331 11339
rect 7849 11305 7883 11339
rect 10241 11305 10275 11339
rect 12633 11305 12667 11339
rect 13277 11305 13311 11339
rect 15761 11305 15795 11339
rect 16313 11305 16347 11339
rect 16681 11305 16715 11339
rect 18705 11305 18739 11339
rect 4997 11237 5031 11271
rect 17592 11237 17626 11271
rect 2421 11169 2455 11203
rect 5917 11169 5951 11203
rect 7205 11169 7239 11203
rect 8217 11169 8251 11203
rect 8309 11169 8343 11203
rect 9781 11169 9815 11203
rect 10609 11169 10643 11203
rect 11621 11169 11655 11203
rect 11713 11169 11747 11203
rect 13645 11169 13679 11203
rect 15669 11169 15703 11203
rect 17325 11169 17359 11203
rect 2513 11101 2547 11135
rect 2605 11101 2639 11135
rect 5089 11101 5123 11135
rect 6009 11101 6043 11135
rect 6193 11101 6227 11135
rect 7481 11101 7515 11135
rect 8401 11101 8435 11135
rect 10701 11101 10735 11135
rect 10793 11101 10827 11135
rect 11805 11101 11839 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 13829 11101 13863 11135
rect 15853 11101 15887 11135
rect 16773 11101 16807 11135
rect 16865 11101 16899 11135
rect 11253 11033 11287 11067
rect 12265 11033 12299 11067
rect 15301 11033 15335 11067
rect 2053 10965 2087 10999
rect 2513 10761 2547 10795
rect 7481 10761 7515 10795
rect 11437 10761 11471 10795
rect 14749 10761 14783 10795
rect 16313 10761 16347 10795
rect 19441 10761 19475 10795
rect 1961 10625 1995 10659
rect 3157 10625 3191 10659
rect 4077 10625 4111 10659
rect 5273 10625 5307 10659
rect 8033 10625 8067 10659
rect 12909 10625 12943 10659
rect 13369 10625 13403 10659
rect 15485 10625 15519 10659
rect 15669 10625 15703 10659
rect 16865 10625 16899 10659
rect 1777 10557 1811 10591
rect 3985 10557 4019 10591
rect 5917 10557 5951 10591
rect 9137 10557 9171 10591
rect 9965 10557 9999 10591
rect 10057 10557 10091 10591
rect 10324 10557 10358 10591
rect 12817 10557 12851 10591
rect 18061 10557 18095 10591
rect 18328 10557 18362 10591
rect 2881 10489 2915 10523
rect 7849 10489 7883 10523
rect 8493 10489 8527 10523
rect 13636 10489 13670 10523
rect 16773 10489 16807 10523
rect 2973 10421 3007 10455
rect 3525 10421 3559 10455
rect 3893 10421 3927 10455
rect 5733 10421 5767 10455
rect 7941 10421 7975 10455
rect 8953 10421 8987 10455
rect 9965 10421 9999 10455
rect 12633 10421 12667 10455
rect 15025 10421 15059 10455
rect 15393 10421 15427 10455
rect 16681 10421 16715 10455
rect 5457 10217 5491 10251
rect 7757 10217 7791 10251
rect 12449 10217 12483 10251
rect 14105 10217 14139 10251
rect 1860 10149 1894 10183
rect 4344 10149 4378 10183
rect 12970 10149 13004 10183
rect 16304 10149 16338 10183
rect 1593 10081 1627 10115
rect 4077 10081 4111 10115
rect 6377 10081 6411 10115
rect 6644 10081 6678 10115
rect 8401 10081 8435 10115
rect 8493 10081 8527 10115
rect 11069 10081 11103 10115
rect 11336 10081 11370 10115
rect 3249 10013 3283 10047
rect 8677 10013 8711 10047
rect 12725 10013 12759 10047
rect 16037 10013 16071 10047
rect 17417 9945 17451 9979
rect 2973 9877 3007 9911
rect 8033 9877 8067 9911
rect 3525 9673 3559 9707
rect 16773 9673 16807 9707
rect 1961 9605 1995 9639
rect 6469 9605 6503 9639
rect 9965 9605 9999 9639
rect 10241 9605 10275 9639
rect 12449 9605 12483 9639
rect 3157 9537 3191 9571
rect 4077 9537 4111 9571
rect 5089 9537 5123 9571
rect 7389 9537 7423 9571
rect 10793 9537 10827 9571
rect 13001 9537 13035 9571
rect 15393 9537 15427 9571
rect 17049 9537 17083 9571
rect 1777 9469 1811 9503
rect 7297 9469 7331 9503
rect 8585 9469 8619 9503
rect 8852 9469 8886 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 15660 9469 15694 9503
rect 2881 9401 2915 9435
rect 3985 9401 4019 9435
rect 5356 9401 5390 9435
rect 10701 9401 10735 9435
rect 2513 9333 2547 9367
rect 2973 9333 3007 9367
rect 3893 9333 3927 9367
rect 6837 9333 6871 9367
rect 7205 9333 7239 9367
rect 10609 9333 10643 9367
rect 1961 9129 1995 9163
rect 2973 9129 3007 9163
rect 6101 9129 6135 9163
rect 8401 9129 8435 9163
rect 2881 9061 2915 9095
rect 1777 8993 1811 9027
rect 6469 8993 6503 9027
rect 7113 8993 7147 9027
rect 8769 8993 8803 9027
rect 3157 8925 3191 8959
rect 6561 8925 6595 8959
rect 6745 8925 6779 8959
rect 8861 8925 8895 8959
rect 9045 8925 9079 8959
rect 2513 8857 2547 8891
rect 9229 8585 9263 8619
rect 3801 8517 3835 8551
rect 1777 8449 1811 8483
rect 4353 8449 4387 8483
rect 5641 8449 5675 8483
rect 7481 8449 7515 8483
rect 2044 8381 2078 8415
rect 5457 8381 5491 8415
rect 7849 8381 7883 8415
rect 8105 8381 8139 8415
rect 4169 8313 4203 8347
rect 7205 8313 7239 8347
rect 7297 8313 7331 8347
rect 3157 8245 3191 8279
rect 4261 8245 4295 8279
rect 6837 8245 6871 8279
rect 4077 8041 4111 8075
rect 4537 8041 4571 8075
rect 5457 8041 5491 8075
rect 6469 8041 6503 8075
rect 7941 8041 7975 8075
rect 8309 8041 8343 8075
rect 8861 8041 8895 8075
rect 19073 8041 19107 8075
rect 2136 7973 2170 8007
rect 5549 7973 5583 8007
rect 1869 7905 1903 7939
rect 4445 7905 4479 7939
rect 4629 7837 4663 7871
rect 5641 7837 5675 7871
rect 6828 7973 6862 8007
rect 8769 7905 8803 7939
rect 18889 7905 18923 7939
rect 6561 7837 6595 7871
rect 8953 7837 8987 7871
rect 4997 7769 5031 7803
rect 6469 7769 6503 7803
rect 3249 7701 3283 7735
rect 5089 7701 5123 7735
rect 8401 7701 8435 7735
rect 4261 7497 4295 7531
rect 19533 7497 19567 7531
rect 2513 7361 2547 7395
rect 7665 7361 7699 7395
rect 8677 7361 8711 7395
rect 2881 7293 2915 7327
rect 4537 7293 4571 7327
rect 4793 7293 4827 7327
rect 7389 7293 7423 7327
rect 8493 7293 8527 7327
rect 19355 7293 19389 7327
rect 2237 7225 2271 7259
rect 3148 7225 3182 7259
rect 7481 7225 7515 7259
rect 1869 7157 1903 7191
rect 2329 7157 2363 7191
rect 5917 7157 5951 7191
rect 6285 7157 6319 7191
rect 7021 7157 7055 7191
rect 8033 7157 8067 7191
rect 8401 7157 8435 7191
rect 2973 6953 3007 6987
rect 7757 6953 7791 6987
rect 5908 6885 5942 6919
rect 7665 6885 7699 6919
rect 1869 6817 1903 6851
rect 3341 6817 3375 6851
rect 4077 6817 4111 6851
rect 5641 6817 5675 6851
rect 19717 6817 19751 6851
rect 20269 6817 20303 6851
rect 2053 6749 2087 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 7849 6749 7883 6783
rect 7021 6681 7055 6715
rect 7297 6681 7331 6715
rect 19901 6681 19935 6715
rect 20453 6681 20487 6715
rect 7113 6409 7147 6443
rect 20729 6409 20763 6443
rect 7665 6273 7699 6307
rect 7481 6205 7515 6239
rect 20551 6205 20585 6239
rect 7573 6069 7607 6103
rect 20729 5321 20763 5355
rect 20545 5117 20579 5151
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2774 20040 2780 20052
rect 1995 20012 2780 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 5353 20043 5411 20049
rect 5353 20040 5365 20043
rect 4571 20012 5365 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 5353 20009 5365 20012
rect 5399 20009 5411 20043
rect 5353 20003 5411 20009
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 5813 20043 5871 20049
rect 5813 20040 5825 20043
rect 5776 20012 5825 20040
rect 5776 20000 5782 20012
rect 5813 20009 5825 20012
rect 5859 20009 5871 20043
rect 5813 20003 5871 20009
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9490 20040 9496 20052
rect 9171 20012 9496 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9490 20000 9496 20012
rect 9548 20000 9554 20052
rect 13173 20043 13231 20049
rect 13173 20009 13185 20043
rect 13219 20040 13231 20043
rect 13630 20040 13636 20052
rect 13219 20012 13636 20040
rect 13219 20009 13231 20012
rect 13173 20003 13231 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15252 20012 15669 20040
rect 15252 20000 15258 20012
rect 15657 20009 15669 20012
rect 15703 20009 15715 20043
rect 15657 20003 15715 20009
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 16632 20012 16773 20040
rect 16632 20000 16638 20012
rect 16761 20009 16773 20012
rect 16807 20009 16819 20043
rect 16761 20003 16819 20009
rect 17313 20043 17371 20049
rect 17313 20009 17325 20043
rect 17359 20040 17371 20043
rect 17402 20040 17408 20052
rect 17359 20012 17408 20040
rect 17359 20009 17371 20012
rect 17313 20003 17371 20009
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18380 20012 18521 20040
rect 18380 20000 18386 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 3513 19907 3571 19913
rect 3513 19873 3525 19907
rect 3559 19904 3571 19907
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3559 19876 4445 19904
rect 3559 19873 3571 19876
rect 3513 19867 3571 19873
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19904 5779 19907
rect 6362 19904 6368 19916
rect 5767 19876 6368 19904
rect 5767 19873 5779 19876
rect 5721 19867 5779 19873
rect 6362 19864 6368 19876
rect 6420 19904 6426 19916
rect 9033 19907 9091 19913
rect 9033 19904 9045 19907
rect 6420 19876 9045 19904
rect 6420 19864 6426 19876
rect 9033 19873 9045 19876
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 11048 19907 11106 19913
rect 11048 19873 11060 19907
rect 11094 19904 11106 19907
rect 11606 19904 11612 19916
rect 11094 19876 11612 19904
rect 11094 19873 11106 19876
rect 11048 19867 11106 19873
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 12989 19907 13047 19913
rect 12989 19904 13001 19907
rect 12860 19876 13001 19904
rect 12860 19864 12866 19876
rect 12989 19873 13001 19876
rect 13035 19873 13047 19907
rect 13814 19904 13820 19916
rect 13775 19876 13820 19904
rect 12989 19867 13047 19873
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 14553 19907 14611 19913
rect 14553 19904 14565 19907
rect 13924 19876 14565 19904
rect 4706 19836 4712 19848
rect 4667 19808 4712 19836
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 5997 19839 6055 19845
rect 5997 19805 6009 19839
rect 6043 19836 6055 19839
rect 6454 19836 6460 19848
rect 6043 19808 6460 19836
rect 6043 19805 6055 19808
rect 5997 19799 6055 19805
rect 6454 19796 6460 19808
rect 6512 19796 6518 19848
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 2866 19768 2872 19780
rect 2547 19740 2872 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 2958 19660 2964 19712
rect 3016 19700 3022 19712
rect 4065 19703 4123 19709
rect 4065 19700 4077 19703
rect 3016 19672 4077 19700
rect 3016 19660 3022 19672
rect 4065 19669 4077 19672
rect 4111 19669 4123 19703
rect 4065 19663 4123 19669
rect 8665 19703 8723 19709
rect 8665 19669 8677 19703
rect 8711 19700 8723 19703
rect 8846 19700 8852 19712
rect 8711 19672 8852 19700
rect 8711 19669 8723 19672
rect 8665 19663 8723 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9324 19700 9352 19799
rect 10318 19796 10324 19848
rect 10376 19836 10382 19848
rect 10781 19839 10839 19845
rect 10781 19836 10793 19839
rect 10376 19808 10793 19836
rect 10376 19796 10382 19808
rect 10781 19805 10793 19808
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 13354 19796 13360 19848
rect 13412 19836 13418 19848
rect 13924 19836 13952 19876
rect 14553 19873 14565 19876
rect 14599 19873 14611 19907
rect 14553 19867 14611 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15252 19876 15485 19904
rect 15252 19864 15258 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19873 16083 19907
rect 16574 19904 16580 19916
rect 16535 19876 16580 19904
rect 16025 19867 16083 19873
rect 14090 19836 14096 19848
rect 13412 19808 13952 19836
rect 14051 19808 14096 19836
rect 13412 19796 13418 19808
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14829 19839 14887 19845
rect 14829 19805 14841 19839
rect 14875 19836 14887 19839
rect 16040 19836 16068 19867
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16666 19864 16672 19916
rect 16724 19904 16730 19916
rect 17129 19907 17187 19913
rect 17129 19904 17141 19907
rect 16724 19876 17141 19904
rect 16724 19864 16730 19876
rect 17129 19873 17141 19876
rect 17175 19873 17187 19907
rect 17129 19867 17187 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18782 19904 18788 19916
rect 18371 19876 18788 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 14875 19808 16068 19836
rect 14875 19805 14887 19808
rect 14829 19799 14887 19805
rect 15562 19728 15568 19780
rect 15620 19768 15626 19780
rect 16209 19771 16267 19777
rect 16209 19768 16221 19771
rect 15620 19740 16221 19768
rect 15620 19728 15626 19740
rect 16209 19737 16221 19740
rect 16255 19737 16267 19771
rect 16209 19731 16267 19737
rect 9858 19700 9864 19712
rect 9324 19672 9864 19700
rect 9858 19660 9864 19672
rect 9916 19700 9922 19712
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 9916 19672 12173 19700
rect 9916 19660 9922 19672
rect 12161 19669 12173 19672
rect 12207 19669 12219 19703
rect 12161 19663 12219 19669
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 2498 19456 2504 19508
rect 2556 19496 2562 19508
rect 6454 19496 6460 19508
rect 2556 19468 6316 19496
rect 6415 19468 6460 19496
rect 2556 19456 2562 19468
rect 6288 19428 6316 19468
rect 6454 19456 6460 19468
rect 6512 19456 6518 19508
rect 7190 19496 7196 19508
rect 6564 19468 7196 19496
rect 6564 19428 6592 19468
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 14645 19499 14703 19505
rect 14645 19496 14657 19499
rect 13872 19468 14657 19496
rect 13872 19456 13878 19468
rect 14645 19465 14657 19468
rect 14691 19465 14703 19499
rect 14645 19459 14703 19465
rect 6288 19400 6592 19428
rect 13740 19400 14320 19428
rect 1762 19320 1768 19372
rect 1820 19360 1826 19372
rect 2317 19363 2375 19369
rect 2317 19360 2329 19363
rect 1820 19332 2329 19360
rect 1820 19320 1826 19332
rect 2317 19329 2329 19332
rect 2363 19329 2375 19363
rect 2317 19323 2375 19329
rect 1578 19292 1584 19304
rect 1539 19264 1584 19292
rect 1578 19252 1584 19264
rect 1636 19252 1642 19304
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 2958 19292 2964 19304
rect 2179 19264 2964 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 3053 19295 3111 19301
rect 3053 19261 3065 19295
rect 3099 19261 3111 19295
rect 3053 19255 3111 19261
rect 198 19184 204 19236
rect 256 19224 262 19236
rect 2406 19224 2412 19236
rect 256 19196 2412 19224
rect 256 19184 262 19196
rect 2406 19184 2412 19196
rect 2464 19184 2470 19236
rect 3068 19224 3096 19255
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3200 19264 5028 19292
rect 3200 19252 3206 19264
rect 3320 19227 3378 19233
rect 3068 19196 3188 19224
rect 1670 19116 1676 19168
rect 1728 19156 1734 19168
rect 1765 19159 1823 19165
rect 1765 19156 1777 19159
rect 1728 19128 1777 19156
rect 1728 19116 1734 19128
rect 1765 19125 1777 19128
rect 1811 19125 1823 19159
rect 3160 19156 3188 19196
rect 3320 19193 3332 19227
rect 3366 19224 3378 19227
rect 5000 19224 5028 19264
rect 5074 19252 5080 19304
rect 5132 19292 5138 19304
rect 6730 19292 6736 19304
rect 5132 19264 5177 19292
rect 5276 19264 6736 19292
rect 5132 19252 5138 19264
rect 5276 19224 5304 19264
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7374 19292 7380 19304
rect 6871 19264 7380 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7374 19252 7380 19264
rect 7432 19292 7438 19304
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 7432 19264 9229 19292
rect 7432 19252 7438 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 10502 19292 10508 19304
rect 9217 19255 9275 19261
rect 9324 19264 10508 19292
rect 3366 19196 4752 19224
rect 5000 19196 5304 19224
rect 5344 19227 5402 19233
rect 3366 19193 3378 19196
rect 3320 19187 3378 19193
rect 4724 19168 4752 19196
rect 5344 19193 5356 19227
rect 5390 19224 5402 19227
rect 5718 19224 5724 19236
rect 5390 19196 5724 19224
rect 5390 19193 5402 19196
rect 5344 19187 5402 19193
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 6454 19184 6460 19236
rect 6512 19224 6518 19236
rect 7070 19227 7128 19233
rect 7070 19224 7082 19227
rect 6512 19196 7082 19224
rect 6512 19184 6518 19196
rect 7070 19193 7082 19196
rect 7116 19193 7128 19227
rect 7070 19187 7128 19193
rect 7190 19184 7196 19236
rect 7248 19224 7254 19236
rect 9324 19224 9352 19264
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11112 19264 11529 19292
rect 11112 19252 11118 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 12618 19252 12624 19304
rect 12676 19292 12682 19304
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12676 19264 12909 19292
rect 12676 19252 12682 19264
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 13740 19292 13768 19400
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14185 19363 14243 19369
rect 14185 19360 14197 19363
rect 13872 19332 14197 19360
rect 13872 19320 13878 19332
rect 14185 19329 14197 19332
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 12897 19255 12955 19261
rect 13004 19264 13768 19292
rect 9490 19233 9496 19236
rect 9484 19224 9496 19233
rect 7248 19196 9352 19224
rect 9451 19196 9496 19224
rect 7248 19184 7254 19196
rect 9484 19187 9496 19196
rect 9490 19184 9496 19187
rect 9548 19184 9554 19236
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 13004 19224 13032 19264
rect 13906 19252 13912 19304
rect 13964 19292 13970 19304
rect 14093 19295 14151 19301
rect 14093 19292 14105 19295
rect 13964 19264 14105 19292
rect 13964 19252 13970 19264
rect 14093 19261 14105 19264
rect 14139 19261 14151 19295
rect 14292 19292 14320 19400
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 15197 19363 15255 19369
rect 15197 19360 15209 19363
rect 15068 19332 15209 19360
rect 15068 19320 15074 19332
rect 15197 19329 15209 19332
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 15746 19292 15752 19304
rect 14292 19264 15752 19292
rect 14093 19255 14151 19261
rect 15746 19252 15752 19264
rect 15804 19252 15810 19304
rect 16114 19292 16120 19304
rect 16075 19264 16120 19292
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16850 19292 16856 19304
rect 16811 19264 16856 19292
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17405 19295 17463 19301
rect 17405 19261 17417 19295
rect 17451 19261 17463 19295
rect 17405 19255 17463 19261
rect 15013 19227 15071 19233
rect 15013 19224 15025 19227
rect 9640 19196 13032 19224
rect 13648 19196 15025 19224
rect 9640 19184 9646 19196
rect 3694 19156 3700 19168
rect 3160 19128 3700 19156
rect 1765 19119 1823 19125
rect 3694 19116 3700 19128
rect 3752 19116 3758 19168
rect 3786 19116 3792 19168
rect 3844 19156 3850 19168
rect 4433 19159 4491 19165
rect 4433 19156 4445 19159
rect 3844 19128 4445 19156
rect 3844 19116 3850 19128
rect 4433 19125 4445 19128
rect 4479 19125 4491 19159
rect 4433 19119 4491 19125
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 8205 19159 8263 19165
rect 8205 19156 8217 19159
rect 4764 19128 8217 19156
rect 4764 19116 4770 19128
rect 8205 19125 8217 19128
rect 8251 19125 8263 19159
rect 8754 19156 8760 19168
rect 8715 19128 8760 19156
rect 8205 19119 8263 19125
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 10597 19159 10655 19165
rect 10597 19156 10609 19159
rect 9732 19128 10609 19156
rect 9732 19116 9738 19128
rect 10597 19125 10609 19128
rect 10643 19125 10655 19159
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 10597 19119 10655 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 12342 19156 12348 19168
rect 11848 19128 12348 19156
rect 11848 19116 11854 19128
rect 12342 19116 12348 19128
rect 12400 19116 12406 19168
rect 13081 19159 13139 19165
rect 13081 19125 13093 19159
rect 13127 19156 13139 19159
rect 13170 19156 13176 19168
rect 13127 19128 13176 19156
rect 13127 19125 13139 19128
rect 13081 19119 13139 19125
rect 13170 19116 13176 19128
rect 13228 19116 13234 19168
rect 13648 19165 13676 19196
rect 15013 19193 15025 19196
rect 15059 19193 15071 19227
rect 15013 19187 15071 19193
rect 16393 19227 16451 19233
rect 16393 19193 16405 19227
rect 16439 19224 16451 19227
rect 17420 19224 17448 19255
rect 17954 19252 17960 19304
rect 18012 19292 18018 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 18012 19264 18061 19292
rect 18012 19252 18018 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18598 19292 18604 19304
rect 18559 19264 18604 19292
rect 18049 19255 18107 19261
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 19153 19295 19211 19301
rect 19153 19292 19165 19295
rect 18800 19264 19165 19292
rect 16439 19196 17448 19224
rect 16439 19193 16451 19196
rect 16393 19187 16451 19193
rect 18138 19184 18144 19236
rect 18196 19224 18202 19236
rect 18800 19224 18828 19264
rect 19153 19261 19165 19264
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 18196 19196 18828 19224
rect 18196 19184 18202 19196
rect 18874 19184 18880 19236
rect 18932 19224 18938 19236
rect 18932 19196 19380 19224
rect 18932 19184 18938 19196
rect 13633 19159 13691 19165
rect 13633 19125 13645 19159
rect 13679 19125 13691 19159
rect 13998 19156 14004 19168
rect 13959 19128 14004 19156
rect 13633 19119 13691 19125
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 15105 19159 15163 19165
rect 15105 19156 15117 19159
rect 14332 19128 15117 19156
rect 14332 19116 14338 19128
rect 15105 19125 15117 19128
rect 15151 19125 15163 19159
rect 15105 19119 15163 19125
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 17037 19159 17095 19165
rect 17037 19156 17049 19159
rect 16080 19128 17049 19156
rect 16080 19116 16086 19128
rect 17037 19125 17049 19128
rect 17083 19125 17095 19159
rect 17037 19119 17095 19125
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17589 19159 17647 19165
rect 17589 19156 17601 19159
rect 17184 19128 17601 19156
rect 17184 19116 17190 19128
rect 17589 19125 17601 19128
rect 17635 19125 17647 19159
rect 17589 19119 17647 19125
rect 17862 19116 17868 19168
rect 17920 19156 17926 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 17920 19128 18245 19156
rect 17920 19116 17926 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 18785 19159 18843 19165
rect 18785 19125 18797 19159
rect 18831 19156 18843 19159
rect 19242 19156 19248 19168
rect 18831 19128 19248 19156
rect 18831 19125 18843 19128
rect 18785 19119 18843 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 19352 19165 19380 19196
rect 19337 19159 19395 19165
rect 19337 19125 19349 19159
rect 19383 19125 19395 19159
rect 19337 19119 19395 19125
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2777 18955 2835 18961
rect 2777 18952 2789 18955
rect 2056 18924 2789 18952
rect 2056 18825 2084 18924
rect 2777 18921 2789 18924
rect 2823 18921 2835 18955
rect 2777 18915 2835 18921
rect 3237 18955 3295 18961
rect 3237 18921 3249 18955
rect 3283 18952 3295 18955
rect 4065 18955 4123 18961
rect 4065 18952 4077 18955
rect 3283 18924 4077 18952
rect 3283 18921 3295 18924
rect 3237 18915 3295 18921
rect 4065 18921 4077 18924
rect 4111 18921 4123 18955
rect 4065 18915 4123 18921
rect 4525 18955 4583 18961
rect 4525 18921 4537 18955
rect 4571 18952 4583 18955
rect 5258 18952 5264 18964
rect 4571 18924 5264 18952
rect 4571 18921 4583 18924
rect 4525 18915 4583 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 8754 18952 8760 18964
rect 6788 18924 8616 18952
rect 8715 18924 8760 18952
rect 6788 18912 6794 18924
rect 2314 18884 2320 18896
rect 2275 18856 2320 18884
rect 2314 18844 2320 18856
rect 2372 18844 2378 18896
rect 7929 18887 7987 18893
rect 7929 18884 7941 18887
rect 2967 18856 7941 18884
rect 2041 18819 2099 18825
rect 2041 18785 2053 18819
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 2406 18776 2412 18828
rect 2464 18816 2470 18828
rect 2967 18816 2995 18856
rect 7929 18853 7941 18856
rect 7975 18853 7987 18887
rect 7929 18847 7987 18853
rect 8297 18887 8355 18893
rect 8297 18853 8309 18887
rect 8343 18884 8355 18887
rect 8588 18884 8616 18924
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 8904 18924 8949 18952
rect 9784 18924 11652 18952
rect 8904 18912 8910 18924
rect 9784 18884 9812 18924
rect 8343 18856 8524 18884
rect 8588 18856 9812 18884
rect 8343 18853 8355 18856
rect 8297 18847 8355 18853
rect 3142 18816 3148 18828
rect 2464 18788 2995 18816
rect 3103 18788 3148 18816
rect 2464 18776 2470 18788
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 4246 18776 4252 18828
rect 4304 18816 4310 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 4304 18788 4445 18816
rect 4304 18776 4310 18788
rect 4433 18785 4445 18788
rect 4479 18816 4491 18819
rect 5445 18819 5503 18825
rect 4479 18788 5396 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 2682 18748 2688 18760
rect 1544 18720 2688 18748
rect 1544 18708 1550 18720
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 3326 18748 3332 18760
rect 3287 18720 3332 18748
rect 3326 18708 3332 18720
rect 3384 18708 3390 18760
rect 3786 18708 3792 18760
rect 3844 18748 3850 18760
rect 4617 18751 4675 18757
rect 4617 18748 4629 18751
rect 3844 18720 4629 18748
rect 3844 18708 3850 18720
rect 4617 18717 4629 18720
rect 4663 18717 4675 18751
rect 4617 18711 4675 18717
rect 5166 18640 5172 18692
rect 5224 18640 5230 18692
rect 5368 18680 5396 18788
rect 5445 18785 5457 18819
rect 5491 18816 5503 18819
rect 6089 18819 6147 18825
rect 6089 18816 6101 18819
rect 5491 18788 6101 18816
rect 5491 18785 5503 18788
rect 5445 18779 5503 18785
rect 6089 18785 6101 18788
rect 6135 18785 6147 18819
rect 6089 18779 6147 18785
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18816 7711 18819
rect 8496 18816 8524 18856
rect 9858 18844 9864 18896
rect 9916 18893 9922 18896
rect 9916 18887 9980 18893
rect 9916 18853 9934 18887
rect 9968 18853 9980 18887
rect 11624 18884 11652 18924
rect 11698 18912 11704 18964
rect 11756 18952 11762 18964
rect 14550 18952 14556 18964
rect 11756 18924 14556 18952
rect 11756 18912 11762 18924
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 18598 18952 18604 18964
rect 17328 18924 18604 18952
rect 11974 18884 11980 18896
rect 11624 18856 11980 18884
rect 9916 18847 9980 18853
rect 9916 18844 9922 18847
rect 11974 18844 11980 18856
rect 12032 18844 12038 18896
rect 12069 18887 12127 18893
rect 12069 18853 12081 18887
rect 12115 18884 12127 18887
rect 12802 18884 12808 18896
rect 12115 18856 12664 18884
rect 12763 18856 12808 18884
rect 12115 18853 12127 18856
rect 12069 18847 12127 18853
rect 9398 18816 9404 18828
rect 7699 18788 8432 18816
rect 8496 18788 9404 18816
rect 7699 18785 7711 18788
rect 7653 18779 7711 18785
rect 5534 18748 5540 18760
rect 5495 18720 5540 18748
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 5718 18748 5724 18760
rect 5631 18720 5724 18748
rect 5718 18708 5724 18720
rect 5776 18748 5782 18760
rect 6454 18748 6460 18760
rect 5776 18720 6460 18748
rect 5776 18708 5782 18720
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 8404 18689 8432 18788
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9640 18788 9689 18816
rect 9640 18776 9646 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 11793 18819 11851 18825
rect 9677 18779 9735 18785
rect 9784 18788 11100 18816
rect 9033 18751 9091 18757
rect 9033 18717 9045 18751
rect 9079 18717 9091 18751
rect 9033 18711 9091 18717
rect 8297 18683 8355 18689
rect 8297 18680 8309 18683
rect 5368 18652 8309 18680
rect 8297 18649 8309 18652
rect 8343 18649 8355 18683
rect 8297 18643 8355 18649
rect 8389 18683 8447 18689
rect 8389 18649 8401 18683
rect 8435 18649 8447 18683
rect 8389 18643 8447 18649
rect 5077 18615 5135 18621
rect 5077 18581 5089 18615
rect 5123 18612 5135 18615
rect 5184 18612 5212 18640
rect 5123 18584 5212 18612
rect 9048 18612 9076 18711
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 9784 18748 9812 18788
rect 9180 18720 9812 18748
rect 9180 18708 9186 18720
rect 11072 18680 11100 18788
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 12158 18816 12164 18828
rect 11839 18788 12164 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12158 18776 12164 18788
rect 12216 18776 12222 18828
rect 12526 18816 12532 18828
rect 12487 18788 12532 18816
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 12636 18816 12664 18856
rect 12802 18844 12808 18856
rect 12860 18844 12866 18896
rect 15194 18884 15200 18896
rect 12912 18856 15200 18884
rect 12912 18816 12940 18856
rect 15194 18844 15200 18856
rect 15252 18844 15258 18896
rect 15749 18887 15807 18893
rect 15749 18853 15761 18887
rect 15795 18884 15807 18887
rect 16850 18884 16856 18896
rect 15795 18856 16856 18884
rect 15795 18853 15807 18856
rect 15749 18847 15807 18853
rect 16850 18844 16856 18856
rect 16908 18844 16914 18896
rect 17328 18893 17356 18924
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 17313 18887 17371 18893
rect 17313 18853 17325 18887
rect 17359 18853 17371 18887
rect 17313 18847 17371 18853
rect 18049 18887 18107 18893
rect 18049 18853 18061 18887
rect 18095 18884 18107 18887
rect 18138 18884 18144 18896
rect 18095 18856 18144 18884
rect 18095 18853 18107 18856
rect 18049 18847 18107 18853
rect 18138 18844 18144 18856
rect 18196 18844 18202 18896
rect 18782 18884 18788 18896
rect 18743 18856 18788 18884
rect 18782 18844 18788 18856
rect 18840 18844 18846 18896
rect 13814 18825 13820 18828
rect 13808 18816 13820 18825
rect 12636 18788 12940 18816
rect 13775 18788 13820 18816
rect 13808 18779 13820 18788
rect 13814 18776 13820 18779
rect 13872 18776 13878 18828
rect 15473 18819 15531 18825
rect 15473 18785 15485 18819
rect 15519 18816 15531 18819
rect 15562 18816 15568 18828
rect 15519 18788 15568 18816
rect 15519 18785 15531 18788
rect 15473 18779 15531 18785
rect 15562 18776 15568 18788
rect 15620 18776 15626 18828
rect 16298 18816 16304 18828
rect 16259 18788 16304 18816
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 16577 18819 16635 18825
rect 16577 18785 16589 18819
rect 16623 18816 16635 18819
rect 16666 18816 16672 18828
rect 16623 18788 16672 18816
rect 16623 18785 16635 18788
rect 16577 18779 16635 18785
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 17037 18819 17095 18825
rect 17037 18785 17049 18819
rect 17083 18785 17095 18819
rect 17037 18779 17095 18785
rect 17773 18819 17831 18825
rect 17773 18785 17785 18819
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 18509 18819 18567 18825
rect 18509 18785 18521 18819
rect 18555 18816 18567 18819
rect 18555 18788 18828 18816
rect 18555 18785 18567 18788
rect 18509 18779 18567 18785
rect 11146 18708 11152 18760
rect 11204 18748 11210 18760
rect 12066 18748 12072 18760
rect 11204 18720 12072 18748
rect 11204 18708 11210 18720
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 13541 18751 13599 18757
rect 13541 18748 13553 18751
rect 12492 18720 13553 18748
rect 12492 18708 12498 18720
rect 13541 18717 13553 18720
rect 13587 18717 13599 18751
rect 13541 18711 13599 18717
rect 16390 18708 16396 18760
rect 16448 18748 16454 18760
rect 17052 18748 17080 18779
rect 16448 18720 17080 18748
rect 16448 18708 16454 18720
rect 11882 18680 11888 18692
rect 11072 18652 11888 18680
rect 11882 18640 11888 18652
rect 11940 18640 11946 18692
rect 15654 18680 15660 18692
rect 14844 18652 15660 18680
rect 9490 18612 9496 18624
rect 9048 18584 9496 18612
rect 5123 18581 5135 18584
rect 5077 18575 5135 18581
rect 9490 18572 9496 18584
rect 9548 18612 9554 18624
rect 11057 18615 11115 18621
rect 11057 18612 11069 18615
rect 9548 18584 11069 18612
rect 9548 18572 9554 18584
rect 11057 18581 11069 18584
rect 11103 18581 11115 18615
rect 11057 18575 11115 18581
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 14844 18612 14872 18652
rect 15654 18640 15660 18652
rect 15712 18640 15718 18692
rect 17788 18680 17816 18779
rect 18800 18760 18828 18788
rect 18782 18708 18788 18760
rect 18840 18708 18846 18760
rect 18506 18680 18512 18692
rect 17788 18652 18512 18680
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 11204 18584 14872 18612
rect 14921 18615 14979 18621
rect 11204 18572 11210 18584
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15010 18612 15016 18624
rect 14967 18584 15016 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 3602 18368 3608 18420
rect 3660 18408 3666 18420
rect 3660 18380 11376 18408
rect 3660 18368 3666 18380
rect 2406 18340 2412 18352
rect 1504 18312 2412 18340
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 1504 18204 1532 18312
rect 2406 18300 2412 18312
rect 2464 18300 2470 18352
rect 3694 18300 3700 18352
rect 3752 18340 3758 18352
rect 4706 18340 4712 18352
rect 3752 18312 4712 18340
rect 3752 18300 3758 18312
rect 4706 18300 4712 18312
rect 4764 18300 4770 18352
rect 6454 18340 6460 18352
rect 6415 18312 6460 18340
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 1578 18232 1584 18284
rect 1636 18272 1642 18284
rect 2133 18275 2191 18281
rect 2133 18272 2145 18275
rect 1636 18244 2145 18272
rect 1636 18232 1642 18244
rect 2133 18241 2145 18244
rect 2179 18241 2191 18275
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 2133 18235 2191 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9493 18275 9551 18281
rect 9493 18272 9505 18275
rect 9088 18244 9505 18272
rect 9088 18232 9094 18244
rect 9493 18241 9505 18244
rect 9539 18241 9551 18275
rect 9674 18272 9680 18284
rect 9635 18244 9680 18272
rect 9493 18235 9551 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 1443 18176 1532 18204
rect 1949 18207 2007 18213
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1949 18173 1961 18207
rect 1995 18204 2007 18207
rect 2314 18204 2320 18216
rect 1995 18176 2320 18204
rect 1995 18173 2007 18176
rect 1949 18167 2007 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2685 18207 2743 18213
rect 2685 18173 2697 18207
rect 2731 18173 2743 18207
rect 2685 18167 2743 18173
rect 2952 18207 3010 18213
rect 2952 18173 2964 18207
rect 2998 18204 3010 18207
rect 3786 18204 3792 18216
rect 2998 18176 3792 18204
rect 2998 18173 3010 18176
rect 2952 18167 3010 18173
rect 1118 18096 1124 18148
rect 1176 18136 1182 18148
rect 2700 18136 2728 18167
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 4706 18164 4712 18216
rect 4764 18204 4770 18216
rect 5074 18204 5080 18216
rect 4764 18176 5080 18204
rect 4764 18164 4770 18176
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 7644 18207 7702 18213
rect 7644 18173 7656 18207
rect 7690 18204 7702 18207
rect 9692 18204 9720 18232
rect 7690 18176 9720 18204
rect 7690 18173 7702 18176
rect 7644 18167 7702 18173
rect 9766 18164 9772 18216
rect 9824 18204 9830 18216
rect 10318 18204 10324 18216
rect 9824 18176 10324 18204
rect 9824 18164 9830 18176
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 11146 18204 11152 18216
rect 10428 18176 11152 18204
rect 3510 18136 3516 18148
rect 1176 18108 1716 18136
rect 2700 18108 3516 18136
rect 1176 18096 1182 18108
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 1688 18068 1716 18108
rect 3510 18096 3516 18108
rect 3568 18096 3574 18148
rect 5344 18139 5402 18145
rect 3620 18108 4200 18136
rect 3620 18068 3648 18108
rect 4062 18068 4068 18080
rect 1688 18040 3648 18068
rect 4023 18040 4068 18068
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4172 18068 4200 18108
rect 5344 18105 5356 18139
rect 5390 18136 5402 18139
rect 5902 18136 5908 18148
rect 5390 18108 5908 18136
rect 5390 18105 5402 18108
rect 5344 18099 5402 18105
rect 5902 18096 5908 18108
rect 5960 18096 5966 18148
rect 10428 18136 10456 18176
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 10594 18145 10600 18148
rect 10588 18136 10600 18145
rect 6012 18108 10456 18136
rect 10555 18108 10600 18136
rect 6012 18068 6040 18108
rect 10588 18099 10600 18108
rect 10594 18096 10600 18099
rect 10652 18096 10658 18148
rect 11348 18136 11376 18380
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 14240 18380 14289 18408
rect 14240 18368 14246 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 13998 18300 14004 18352
rect 14056 18340 14062 18352
rect 14056 18312 15700 18340
rect 14056 18300 14062 18312
rect 15194 18272 15200 18284
rect 14200 18244 15200 18272
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 12434 18204 12440 18216
rect 12308 18176 12440 18204
rect 12308 18164 12314 18176
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 12492 18176 12537 18204
rect 12636 18176 13921 18204
rect 12492 18164 12498 18176
rect 12636 18136 12664 18176
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 14090 18204 14096 18216
rect 14051 18176 14096 18204
rect 13909 18167 13967 18173
rect 14090 18164 14096 18176
rect 14148 18164 14154 18216
rect 11348 18108 12664 18136
rect 12704 18139 12762 18145
rect 12704 18105 12716 18139
rect 12750 18136 12762 18139
rect 12986 18136 12992 18148
rect 12750 18108 12992 18136
rect 12750 18105 12762 18108
rect 12704 18099 12762 18105
rect 12986 18096 12992 18108
rect 13044 18136 13050 18148
rect 14200 18136 14228 18244
rect 15194 18232 15200 18244
rect 15252 18232 15258 18284
rect 15672 18281 15700 18312
rect 17770 18300 17776 18352
rect 17828 18340 17834 18352
rect 22462 18340 22468 18352
rect 17828 18312 22468 18340
rect 17828 18300 17834 18312
rect 22462 18300 22468 18312
rect 22520 18300 22526 18352
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18241 15715 18275
rect 16574 18272 16580 18284
rect 16535 18244 16580 18272
rect 15657 18235 15715 18241
rect 16574 18232 16580 18244
rect 16632 18232 16638 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 18012 18244 18245 18272
rect 18012 18232 18018 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 14366 18164 14372 18216
rect 14424 18204 14430 18216
rect 15013 18207 15071 18213
rect 15013 18204 15025 18207
rect 14424 18176 15025 18204
rect 14424 18164 14430 18176
rect 15013 18173 15025 18176
rect 15059 18173 15071 18207
rect 15013 18167 15071 18173
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16301 18207 16359 18213
rect 16301 18204 16313 18207
rect 15896 18176 16313 18204
rect 15896 18164 15902 18176
rect 16301 18173 16313 18176
rect 16347 18173 16359 18207
rect 16301 18167 16359 18173
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 19058 18204 19064 18216
rect 18095 18176 19064 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 15102 18136 15108 18148
rect 13044 18108 14228 18136
rect 14384 18108 15108 18136
rect 13044 18096 13050 18108
rect 4172 18040 6040 18068
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 7558 18068 7564 18080
rect 6328 18040 7564 18068
rect 6328 18028 6334 18040
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 8754 18068 8760 18080
rect 8715 18040 8760 18068
rect 8754 18028 8760 18040
rect 8812 18028 8818 18080
rect 9030 18068 9036 18080
rect 8991 18040 9036 18068
rect 9030 18028 9036 18040
rect 9088 18028 9094 18080
rect 9398 18068 9404 18080
rect 9359 18040 9404 18068
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 11146 18068 11152 18080
rect 10468 18040 11152 18068
rect 10468 18028 10474 18040
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 11698 18068 11704 18080
rect 11659 18040 11704 18068
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 13814 18068 13820 18080
rect 13775 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 14384 18068 14412 18108
rect 15102 18096 15108 18108
rect 15160 18096 15166 18148
rect 19518 18096 19524 18148
rect 19576 18136 19582 18148
rect 20162 18136 20168 18148
rect 19576 18108 20168 18136
rect 19576 18096 19582 18108
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 22002 18136 22008 18148
rect 20864 18108 22008 18136
rect 20864 18096 20870 18108
rect 22002 18096 22008 18108
rect 22060 18096 22066 18148
rect 13955 18040 14412 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 14550 18028 14556 18080
rect 14608 18068 14614 18080
rect 14645 18071 14703 18077
rect 14645 18068 14657 18071
rect 14608 18040 14657 18068
rect 14608 18028 14614 18040
rect 14645 18037 14657 18040
rect 14691 18037 14703 18071
rect 14645 18031 14703 18037
rect 19886 18028 19892 18080
rect 19944 18068 19950 18080
rect 20622 18068 20628 18080
rect 19944 18040 20628 18068
rect 19944 18028 19950 18040
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 21542 18068 21548 18080
rect 20956 18040 21548 18068
rect 20956 18028 20962 18040
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2501 17867 2559 17873
rect 2501 17833 2513 17867
rect 2547 17864 2559 17867
rect 2774 17864 2780 17876
rect 2547 17836 2780 17864
rect 2547 17833 2559 17836
rect 2501 17827 2559 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 3050 17864 3056 17876
rect 3011 17836 3056 17864
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3142 17824 3148 17876
rect 3200 17864 3206 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3200 17836 3433 17864
rect 3200 17824 3206 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 3421 17827 3479 17833
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5592 17836 5641 17864
rect 5592 17824 5598 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 6089 17867 6147 17873
rect 6089 17833 6101 17867
rect 6135 17864 6147 17867
rect 6178 17864 6184 17876
rect 6135 17836 6184 17864
rect 6135 17833 6147 17836
rect 6089 17827 6147 17833
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 8021 17867 8079 17873
rect 6748 17836 7972 17864
rect 2332 17768 4936 17796
rect 1762 17728 1768 17740
rect 1723 17700 1768 17728
rect 1762 17688 1768 17700
rect 1820 17688 1826 17740
rect 2332 17737 2360 17768
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 2317 17691 2375 17697
rect 2406 17688 2412 17740
rect 2464 17728 2470 17740
rect 2869 17731 2927 17737
rect 2869 17728 2881 17731
rect 2464 17700 2881 17728
rect 2464 17688 2470 17700
rect 2869 17697 2881 17700
rect 2915 17697 2927 17731
rect 2869 17691 2927 17697
rect 3326 17688 3332 17740
rect 3384 17728 3390 17740
rect 4062 17728 4068 17740
rect 3384 17700 4068 17728
rect 3384 17688 3390 17700
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4908 17592 4936 17768
rect 5997 17731 6055 17737
rect 5997 17697 6009 17731
rect 6043 17728 6055 17731
rect 6748 17728 6776 17836
rect 7469 17799 7527 17805
rect 7469 17796 7481 17799
rect 6840 17768 7481 17796
rect 6840 17737 6868 17768
rect 7469 17765 7481 17768
rect 7515 17765 7527 17799
rect 7944 17796 7972 17836
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 9030 17864 9036 17876
rect 8067 17836 9036 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 9950 17824 9956 17876
rect 10008 17864 10014 17876
rect 10413 17867 10471 17873
rect 10413 17864 10425 17867
rect 10008 17836 10425 17864
rect 10008 17824 10014 17836
rect 10413 17833 10425 17836
rect 10459 17833 10471 17867
rect 10413 17827 10471 17833
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 13906 17864 13912 17876
rect 12483 17836 13912 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 14274 17864 14280 17876
rect 14231 17836 14280 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14550 17864 14556 17876
rect 14511 17836 14556 17864
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 14645 17867 14703 17873
rect 14645 17833 14657 17867
rect 14691 17864 14703 17867
rect 15289 17867 15347 17873
rect 15289 17864 15301 17867
rect 14691 17836 15301 17864
rect 14691 17833 14703 17836
rect 14645 17827 14703 17833
rect 15289 17833 15301 17836
rect 15335 17833 15347 17867
rect 15654 17864 15660 17876
rect 15615 17836 15660 17864
rect 15289 17827 15347 17833
rect 15654 17824 15660 17836
rect 15712 17864 15718 17876
rect 16022 17864 16028 17876
rect 15712 17836 16028 17864
rect 15712 17824 15718 17836
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 9398 17796 9404 17808
rect 7944 17768 9404 17796
rect 7469 17759 7527 17765
rect 9398 17756 9404 17768
rect 9456 17756 9462 17808
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 12250 17796 12256 17808
rect 9824 17768 12256 17796
rect 9824 17756 9830 17768
rect 12250 17756 12256 17768
rect 12308 17756 12314 17808
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 15252 17768 15792 17796
rect 15252 17756 15258 17768
rect 6043 17700 6776 17728
rect 6825 17731 6883 17737
rect 6043 17697 6055 17700
rect 5997 17691 6055 17697
rect 6825 17697 6837 17731
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7147 17700 7389 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7926 17728 7932 17740
rect 7887 17700 7932 17728
rect 7377 17691 7435 17697
rect 7926 17688 7932 17700
rect 7984 17688 7990 17740
rect 8849 17731 8907 17737
rect 8849 17697 8861 17731
rect 8895 17728 8907 17731
rect 9950 17728 9956 17740
rect 8895 17700 9956 17728
rect 8895 17697 8907 17700
rect 8849 17691 8907 17697
rect 9950 17688 9956 17700
rect 10008 17688 10014 17740
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17697 10379 17731
rect 12802 17728 12808 17740
rect 12763 17700 12808 17728
rect 10321 17691 10379 17697
rect 5902 17620 5908 17672
rect 5960 17660 5966 17672
rect 6181 17663 6239 17669
rect 6181 17660 6193 17663
rect 5960 17632 6193 17660
rect 5960 17620 5966 17632
rect 6181 17629 6193 17632
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17660 8263 17663
rect 8294 17660 8300 17672
rect 8251 17632 8300 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 8294 17620 8300 17632
rect 8352 17660 8358 17672
rect 8754 17660 8760 17672
rect 8352 17632 8760 17660
rect 8352 17620 8358 17632
rect 8754 17620 8760 17632
rect 8812 17620 8818 17672
rect 9033 17663 9091 17669
rect 9033 17629 9045 17663
rect 9079 17629 9091 17663
rect 9033 17623 9091 17629
rect 7377 17595 7435 17601
rect 7377 17592 7389 17595
rect 4908 17564 7389 17592
rect 7377 17561 7389 17564
rect 7423 17561 7435 17595
rect 7377 17555 7435 17561
rect 7469 17595 7527 17601
rect 7469 17561 7481 17595
rect 7515 17592 7527 17595
rect 7561 17595 7619 17601
rect 7561 17592 7573 17595
rect 7515 17564 7573 17592
rect 7515 17561 7527 17564
rect 7469 17555 7527 17561
rect 7561 17561 7573 17564
rect 7607 17561 7619 17595
rect 7561 17555 7619 17561
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 9048 17524 9076 17623
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 10336 17660 10364 17691
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 15764 17728 15792 17768
rect 17126 17756 17132 17808
rect 17184 17805 17190 17808
rect 17184 17799 17248 17805
rect 17184 17765 17202 17799
rect 17236 17765 17248 17799
rect 17184 17759 17248 17765
rect 17184 17756 17190 17759
rect 17770 17728 17776 17740
rect 15764 17700 15884 17728
rect 10594 17660 10600 17672
rect 9456 17632 10364 17660
rect 10555 17632 10600 17660
rect 9456 17620 9462 17632
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10962 17660 10968 17672
rect 10923 17632 10968 17660
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17629 12955 17663
rect 12897 17623 12955 17629
rect 12912 17592 12940 17623
rect 12986 17620 12992 17672
rect 13044 17660 13050 17672
rect 13044 17632 13089 17660
rect 13044 17620 13050 17632
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 13872 17632 14749 17660
rect 13872 17620 13878 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 15654 17620 15660 17672
rect 15712 17660 15718 17672
rect 15856 17669 15884 17700
rect 15948 17700 17776 17728
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15712 17632 15761 17660
rect 15712 17620 15718 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15948 17592 15976 17700
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 16945 17663 17003 17669
rect 16945 17660 16957 17663
rect 16540 17632 16957 17660
rect 16540 17620 16546 17632
rect 16945 17629 16957 17632
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 12912 17564 15976 17592
rect 5868 17496 9076 17524
rect 9953 17527 10011 17533
rect 5868 17484 5874 17496
rect 9953 17493 9965 17527
rect 9999 17524 10011 17527
rect 10410 17524 10416 17536
rect 9999 17496 10416 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 18325 17527 18383 17533
rect 18325 17493 18337 17527
rect 18371 17524 18383 17527
rect 18598 17524 18604 17536
rect 18371 17496 18604 17524
rect 18371 17493 18383 17496
rect 18325 17487 18383 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 5810 17320 5816 17332
rect 1504 17292 5816 17320
rect 1504 17125 1532 17292
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 5960 17292 6193 17320
rect 5960 17280 5966 17292
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7653 17323 7711 17329
rect 7653 17320 7665 17323
rect 7432 17292 7665 17320
rect 7432 17280 7438 17292
rect 7653 17289 7665 17292
rect 7699 17289 7711 17323
rect 9950 17320 9956 17332
rect 9911 17292 9956 17320
rect 7653 17283 7711 17289
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 13538 17320 13544 17332
rect 12768 17292 13544 17320
rect 12768 17280 12774 17292
rect 13538 17280 13544 17292
rect 13596 17280 13602 17332
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 14424 17292 15424 17320
rect 14424 17280 14430 17292
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2406 17184 2412 17196
rect 2363 17156 2412 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 7926 17184 7932 17196
rect 7887 17156 7932 17184
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 10410 17184 10416 17196
rect 10371 17156 10416 17184
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 11698 17184 11704 17196
rect 10643 17156 11704 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 12492 17156 12541 17184
rect 12492 17144 12498 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 2038 17116 2044 17128
rect 1999 17088 2044 17116
rect 1489 17079 1547 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 3044 17119 3102 17125
rect 3044 17085 3056 17119
rect 3090 17116 3102 17119
rect 3326 17116 3332 17128
rect 3090 17088 3332 17116
rect 3090 17085 3102 17088
rect 3044 17079 3102 17085
rect 2792 17048 2820 17079
rect 3326 17076 3332 17088
rect 3384 17076 3390 17128
rect 4706 17076 4712 17128
rect 4764 17116 4770 17128
rect 4801 17119 4859 17125
rect 4801 17116 4813 17119
rect 4764 17088 4813 17116
rect 4764 17076 4770 17088
rect 4801 17085 4813 17088
rect 4847 17085 4859 17119
rect 4801 17079 4859 17085
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7064 17088 7849 17116
rect 7064 17076 7070 17088
rect 7837 17085 7849 17088
rect 7883 17085 7895 17119
rect 7837 17079 7895 17085
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17116 8815 17119
rect 9674 17116 9680 17128
rect 8803 17088 9680 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 10321 17119 10379 17125
rect 10321 17085 10333 17119
rect 10367 17116 10379 17119
rect 10962 17116 10968 17128
rect 10367 17088 10968 17116
rect 10367 17085 10379 17088
rect 10321 17079 10379 17085
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 12069 17119 12127 17125
rect 12069 17085 12081 17119
rect 12115 17116 12127 17119
rect 13262 17116 13268 17128
rect 12115 17088 13268 17116
rect 12115 17085 12127 17088
rect 12069 17079 12127 17085
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 14636 17119 14694 17125
rect 14636 17085 14648 17119
rect 14682 17116 14694 17119
rect 15010 17116 15016 17128
rect 14682 17088 15016 17116
rect 14682 17085 14694 17088
rect 14636 17079 14694 17085
rect 4724 17048 4752 17076
rect 2792 17020 4752 17048
rect 5068 17051 5126 17057
rect 5068 17017 5080 17051
rect 5114 17048 5126 17051
rect 5258 17048 5264 17060
rect 5114 17020 5264 17048
rect 5114 17017 5126 17020
rect 5068 17011 5126 17017
rect 5258 17008 5264 17020
rect 5316 17008 5322 17060
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 9033 17051 9091 17057
rect 9033 17048 9045 17051
rect 6972 17020 9045 17048
rect 6972 17008 6978 17020
rect 9033 17017 9045 17020
rect 9079 17017 9091 17051
rect 9033 17011 9091 17017
rect 12796 17051 12854 17057
rect 12796 17017 12808 17051
rect 12842 17048 12854 17051
rect 13078 17048 13084 17060
rect 12842 17020 13084 17048
rect 12842 17017 12854 17020
rect 12796 17011 12854 17017
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 14384 17048 14412 17079
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15396 17116 15424 17292
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 16485 17323 16543 17329
rect 16485 17320 16497 17323
rect 16356 17292 16497 17320
rect 16356 17280 16362 17292
rect 16485 17289 16497 17292
rect 16531 17289 16543 17323
rect 19058 17320 19064 17332
rect 19019 17292 19064 17320
rect 16485 17283 16543 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 18049 17255 18107 17261
rect 18049 17221 18061 17255
rect 18095 17252 18107 17255
rect 18095 17224 19564 17252
rect 18095 17221 18107 17224
rect 18049 17215 18107 17221
rect 17126 17184 17132 17196
rect 17087 17156 17132 17184
rect 17126 17144 17132 17156
rect 17184 17144 17190 17196
rect 18598 17184 18604 17196
rect 18559 17156 18604 17184
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 19536 17193 19564 17224
rect 19521 17187 19579 17193
rect 19521 17153 19533 17187
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 18417 17119 18475 17125
rect 15396 17088 16988 17116
rect 15470 17048 15476 17060
rect 14384 17020 15476 17048
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 16025 17051 16083 17057
rect 16025 17017 16037 17051
rect 16071 17048 16083 17051
rect 16853 17051 16911 17057
rect 16853 17048 16865 17051
rect 16071 17020 16865 17048
rect 16071 17017 16083 17020
rect 16025 17011 16083 17017
rect 16853 17017 16865 17020
rect 16899 17017 16911 17051
rect 16960 17048 16988 17088
rect 18417 17085 18429 17119
rect 18463 17116 18475 17119
rect 18966 17116 18972 17128
rect 18463 17088 18972 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 18966 17076 18972 17088
rect 19024 17076 19030 17128
rect 19150 17076 19156 17128
rect 19208 17116 19214 17128
rect 19628 17116 19656 17147
rect 19208 17088 19656 17116
rect 19208 17076 19214 17088
rect 17497 17051 17555 17057
rect 16960 17020 17080 17048
rect 16853 17011 16911 17017
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 4157 16983 4215 16989
rect 4157 16980 4169 16983
rect 4120 16952 4169 16980
rect 4120 16940 4126 16952
rect 4157 16949 4169 16952
rect 4203 16949 4215 16983
rect 4157 16943 4215 16949
rect 11885 16983 11943 16989
rect 11885 16949 11897 16983
rect 11931 16980 11943 16983
rect 12434 16980 12440 16992
rect 11931 16952 12440 16980
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 12434 16940 12440 16952
rect 12492 16980 12498 16992
rect 12894 16980 12900 16992
rect 12492 16952 12900 16980
rect 12492 16940 12498 16952
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 12986 16940 12992 16992
rect 13044 16980 13050 16992
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13044 16952 13921 16980
rect 13044 16940 13050 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 13909 16943 13967 16949
rect 14550 16940 14556 16992
rect 14608 16980 14614 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 14608 16952 15761 16980
rect 14608 16940 14614 16952
rect 15749 16949 15761 16952
rect 15795 16949 15807 16983
rect 16942 16980 16948 16992
rect 16903 16952 16948 16980
rect 15749 16943 15807 16949
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17052 16980 17080 17020
rect 17497 17017 17509 17051
rect 17543 17048 17555 17051
rect 19429 17051 19487 17057
rect 19429 17048 19441 17051
rect 17543 17020 19441 17048
rect 17543 17017 17555 17020
rect 17497 17011 17555 17017
rect 19429 17017 19441 17020
rect 19475 17017 19487 17051
rect 19429 17011 19487 17017
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 17052 16952 18521 16980
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1765 16779 1823 16785
rect 1765 16745 1777 16779
rect 1811 16745 1823 16779
rect 1765 16739 1823 16745
rect 1780 16708 1808 16739
rect 2038 16736 2044 16788
rect 2096 16776 2102 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 2096 16748 4537 16776
rect 2096 16736 2102 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 4985 16779 5043 16785
rect 4985 16745 4997 16779
rect 5031 16776 5043 16779
rect 5537 16779 5595 16785
rect 5537 16776 5549 16779
rect 5031 16748 5549 16776
rect 5031 16745 5043 16748
rect 4985 16739 5043 16745
rect 5537 16745 5549 16748
rect 5583 16745 5595 16779
rect 5537 16739 5595 16745
rect 5997 16779 6055 16785
rect 5997 16745 6009 16779
rect 6043 16776 6055 16779
rect 6638 16776 6644 16788
rect 6043 16748 6644 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6638 16736 6644 16748
rect 6696 16736 6702 16788
rect 10594 16736 10600 16788
rect 10652 16776 10658 16788
rect 11149 16779 11207 16785
rect 11149 16776 11161 16779
rect 10652 16748 11161 16776
rect 10652 16736 10658 16748
rect 11149 16745 11161 16748
rect 11195 16745 11207 16779
rect 11149 16739 11207 16745
rect 12345 16779 12403 16785
rect 12345 16745 12357 16779
rect 12391 16776 12403 16779
rect 12526 16776 12532 16788
rect 12391 16748 12532 16776
rect 12391 16745 12403 16748
rect 12345 16739 12403 16745
rect 12526 16736 12532 16748
rect 12584 16736 12590 16788
rect 17126 16736 17132 16788
rect 17184 16776 17190 16788
rect 17313 16779 17371 16785
rect 17313 16776 17325 16779
rect 17184 16748 17325 16776
rect 17184 16736 17190 16748
rect 17313 16745 17325 16748
rect 17359 16745 17371 16779
rect 17313 16739 17371 16745
rect 3234 16708 3240 16720
rect 1780 16680 3240 16708
rect 3234 16668 3240 16680
rect 3292 16668 3298 16720
rect 4893 16711 4951 16717
rect 4893 16677 4905 16711
rect 4939 16708 4951 16711
rect 6549 16711 6607 16717
rect 6549 16708 6561 16711
rect 4939 16680 6561 16708
rect 4939 16677 4951 16680
rect 4893 16671 4951 16677
rect 6549 16677 6561 16680
rect 6595 16677 6607 16711
rect 6549 16671 6607 16677
rect 7552 16711 7610 16717
rect 7552 16677 7564 16711
rect 7598 16708 7610 16711
rect 8294 16708 8300 16720
rect 7598 16680 8300 16708
rect 7598 16677 7610 16680
rect 7552 16671 7610 16677
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 16482 16708 16488 16720
rect 15948 16680 16488 16708
rect 15948 16652 15976 16680
rect 16482 16668 16488 16680
rect 16540 16708 16546 16720
rect 18040 16711 18098 16717
rect 16540 16680 17816 16708
rect 16540 16668 16546 16680
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 2038 16640 2044 16652
rect 1627 16612 2044 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 5534 16640 5540 16652
rect 2179 16612 5540 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5905 16643 5963 16649
rect 5905 16609 5917 16643
rect 5951 16640 5963 16643
rect 7098 16640 7104 16652
rect 5951 16612 7104 16640
rect 5951 16609 5963 16612
rect 5905 16603 5963 16609
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 7285 16643 7343 16649
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 7374 16640 7380 16652
rect 7331 16612 7380 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 9766 16640 9772 16652
rect 9727 16612 9772 16640
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 10036 16643 10094 16649
rect 10036 16609 10048 16643
rect 10082 16640 10094 16643
rect 10778 16640 10784 16652
rect 10082 16612 10784 16640
rect 10082 16609 10094 16612
rect 10036 16603 10094 16609
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 15930 16640 15936 16652
rect 15843 16612 15936 16640
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16206 16649 16212 16652
rect 16200 16640 16212 16649
rect 16167 16612 16212 16640
rect 16200 16603 16212 16612
rect 16206 16600 16212 16603
rect 16264 16600 16270 16652
rect 17788 16649 17816 16680
rect 18040 16677 18052 16711
rect 18086 16708 18098 16711
rect 18598 16708 18604 16720
rect 18086 16680 18604 16708
rect 18086 16677 18098 16680
rect 18040 16671 18098 16677
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 17862 16640 17868 16652
rect 17819 16612 17868 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 1762 16532 1768 16584
rect 1820 16572 1826 16584
rect 2317 16575 2375 16581
rect 2317 16572 2329 16575
rect 1820 16544 2329 16572
rect 1820 16532 1826 16544
rect 2317 16541 2329 16544
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16572 5227 16575
rect 5258 16572 5264 16584
rect 5215 16544 5264 16572
rect 5215 16541 5227 16544
rect 5169 16535 5227 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12805 16575 12863 16581
rect 12805 16572 12817 16575
rect 12492 16544 12817 16572
rect 12492 16532 12498 16544
rect 12805 16541 12817 16544
rect 12851 16541 12863 16575
rect 12805 16535 12863 16541
rect 12989 16575 13047 16581
rect 12989 16541 13001 16575
rect 13035 16572 13047 16575
rect 13078 16572 13084 16584
rect 13035 16544 13084 16572
rect 13035 16541 13047 16544
rect 12989 16535 13047 16541
rect 13078 16532 13084 16544
rect 13136 16532 13142 16584
rect 8662 16436 8668 16448
rect 8623 16408 8668 16436
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 19150 16436 19156 16448
rect 19111 16408 19156 16436
rect 19150 16396 19156 16408
rect 19208 16396 19214 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 5258 16192 5264 16244
rect 5316 16232 5322 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5316 16204 6009 16232
rect 5316 16192 5322 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 7098 16192 7104 16244
rect 7156 16232 7162 16244
rect 10778 16232 10784 16244
rect 7156 16204 7880 16232
rect 10739 16204 10784 16232
rect 7156 16192 7162 16204
rect 2038 16056 2044 16108
rect 2096 16096 2102 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 2096 16068 2145 16096
rect 2096 16056 2102 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 4062 16096 4068 16108
rect 4023 16068 4068 16096
rect 2133 16059 2191 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 7852 16096 7880 16204
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 13078 16192 13084 16244
rect 13136 16232 13142 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13136 16204 13829 16232
rect 13136 16192 13142 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 15289 16235 15347 16241
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15470 16232 15476 16244
rect 15335 16204 15476 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 15565 16235 15623 16241
rect 15565 16201 15577 16235
rect 15611 16232 15623 16235
rect 16942 16232 16948 16244
rect 15611 16204 16948 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 14292 16136 15516 16164
rect 5736 16068 6960 16096
rect 7852 16068 9536 16096
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2498 16028 2504 16040
rect 1995 16000 2504 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 1412 15960 1440 15991
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 2682 16028 2688 16040
rect 2643 16000 2688 16028
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 2924 16000 3801 16028
rect 2924 15988 2930 16000
rect 3789 15997 3801 16000
rect 3835 16028 3847 16031
rect 4522 16028 4528 16040
rect 3835 16000 4528 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 4522 15988 4528 16000
rect 4580 15988 4586 16040
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 4706 16028 4712 16040
rect 4663 16000 4712 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 5736 16028 5764 16068
rect 6932 16040 6960 16068
rect 4816 16000 5764 16028
rect 6825 16031 6883 16037
rect 4816 15960 4844 16000
rect 6825 15997 6837 16031
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 1412 15932 4844 15960
rect 4884 15963 4942 15969
rect 4884 15929 4896 15963
rect 4930 15960 4942 15963
rect 6086 15960 6092 15972
rect 4930 15932 6092 15960
rect 4930 15929 4942 15932
rect 4884 15923 4942 15929
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 6840 15960 6868 15991
rect 6914 15988 6920 16040
rect 6972 15988 6978 16040
rect 7374 16028 7380 16040
rect 7024 16000 7380 16028
rect 7024 15960 7052 16000
rect 7374 15988 7380 16000
rect 7432 16028 7438 16040
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 7432 16000 9413 16028
rect 7432 15988 7438 16000
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 6840 15932 7052 15960
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 8662 15960 8668 15972
rect 7138 15932 8668 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 9508 15960 9536 16068
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11204 16068 11529 16096
rect 11204 16056 11210 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 11609 16099 11667 16105
rect 11609 16065 11621 16099
rect 11655 16065 11667 16099
rect 11609 16059 11667 16065
rect 9668 16031 9726 16037
rect 9668 15997 9680 16031
rect 9714 16028 9726 16031
rect 9950 16028 9956 16040
rect 9714 16000 9956 16028
rect 9714 15997 9726 16000
rect 9668 15991 9726 15997
rect 9950 15988 9956 16000
rect 10008 16028 10014 16040
rect 11624 16028 11652 16059
rect 10008 16000 11652 16028
rect 12437 16031 12495 16037
rect 10008 15988 10014 16000
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12483 16000 12940 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12912 15972 12940 16000
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 14292 16028 14320 16136
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14424 16068 14657 16096
rect 14424 16056 14430 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 15488 16037 15516 16136
rect 16206 16096 16212 16108
rect 16167 16068 16212 16096
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 13320 16000 14320 16028
rect 15473 16031 15531 16037
rect 13320 15988 13326 16000
rect 15473 15997 15485 16031
rect 15519 15997 15531 16031
rect 15473 15991 15531 15997
rect 11425 15963 11483 15969
rect 11425 15960 11437 15963
rect 9508 15932 11437 15960
rect 11425 15929 11437 15932
rect 11471 15929 11483 15963
rect 11425 15923 11483 15929
rect 12618 15920 12624 15972
rect 12676 15969 12682 15972
rect 12676 15963 12740 15969
rect 12676 15929 12694 15963
rect 12728 15929 12740 15963
rect 12676 15923 12740 15929
rect 12676 15920 12682 15923
rect 12894 15920 12900 15972
rect 12952 15920 12958 15972
rect 14553 15963 14611 15969
rect 14553 15960 14565 15963
rect 13004 15932 14565 15960
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 3421 15895 3479 15901
rect 3421 15892 3433 15895
rect 3108 15864 3433 15892
rect 3108 15852 3114 15864
rect 3421 15861 3433 15864
rect 3467 15861 3479 15895
rect 3421 15855 3479 15861
rect 3881 15895 3939 15901
rect 3881 15861 3893 15895
rect 3927 15892 3939 15895
rect 4798 15892 4804 15904
rect 3927 15864 4804 15892
rect 3927 15861 3939 15864
rect 3881 15855 3939 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 6273 15895 6331 15901
rect 6273 15861 6285 15895
rect 6319 15892 6331 15895
rect 6914 15892 6920 15904
rect 6319 15864 6920 15892
rect 6319 15861 6331 15864
rect 6273 15855 6331 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7248 15864 8217 15892
rect 7248 15852 7254 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 8941 15895 8999 15901
rect 8941 15861 8953 15895
rect 8987 15892 8999 15895
rect 10042 15892 10048 15904
rect 8987 15864 10048 15892
rect 8987 15861 8999 15864
rect 8941 15855 8999 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 11054 15892 11060 15904
rect 11015 15864 11060 15892
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12250 15852 12256 15904
rect 12308 15892 12314 15904
rect 13004 15892 13032 15932
rect 14553 15929 14565 15932
rect 14599 15960 14611 15963
rect 16025 15963 16083 15969
rect 16025 15960 16037 15963
rect 14599 15932 16037 15960
rect 14599 15929 14611 15932
rect 14553 15923 14611 15929
rect 16025 15929 16037 15932
rect 16071 15929 16083 15963
rect 16025 15923 16083 15929
rect 14090 15892 14096 15904
rect 12308 15864 13032 15892
rect 14051 15864 14096 15892
rect 12308 15852 12314 15864
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 14458 15892 14464 15904
rect 14419 15864 14464 15892
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15933 15895 15991 15901
rect 15933 15892 15945 15895
rect 15436 15864 15945 15892
rect 15436 15852 15442 15864
rect 15933 15861 15945 15864
rect 15979 15861 15991 15895
rect 15933 15855 15991 15861
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6549 15691 6607 15697
rect 6549 15688 6561 15691
rect 5592 15660 6561 15688
rect 5592 15648 5598 15660
rect 6549 15657 6561 15660
rect 6595 15657 6607 15691
rect 6914 15688 6920 15700
rect 6875 15660 6920 15688
rect 6549 15651 6607 15657
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 7009 15691 7067 15697
rect 7009 15657 7021 15691
rect 7055 15688 7067 15691
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7055 15660 7573 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 7561 15651 7619 15657
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8202 15688 8208 15700
rect 8067 15660 8208 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 11054 15688 11060 15700
rect 10183 15660 11060 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15657 11483 15691
rect 11425 15651 11483 15657
rect 2584 15623 2642 15629
rect 2584 15589 2596 15623
rect 2630 15620 2642 15623
rect 4062 15620 4068 15632
rect 2630 15592 4068 15620
rect 2630 15589 2642 15592
rect 2584 15583 2642 15589
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 4522 15580 4528 15632
rect 4580 15620 4586 15632
rect 7929 15623 7987 15629
rect 7929 15620 7941 15623
rect 4580 15592 7941 15620
rect 4580 15580 4586 15592
rect 7929 15589 7941 15592
rect 7975 15589 7987 15623
rect 11440 15620 11468 15651
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12805 15691 12863 15697
rect 12492 15660 12537 15688
rect 12492 15648 12498 15660
rect 12805 15657 12817 15691
rect 12851 15688 12863 15691
rect 14090 15688 14096 15700
rect 12851 15660 14096 15688
rect 12851 15657 12863 15660
rect 12805 15651 12863 15657
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 16206 15648 16212 15700
rect 16264 15688 16270 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 16264 15660 17141 15688
rect 16264 15648 16270 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17129 15651 17187 15657
rect 12710 15620 12716 15632
rect 11440 15592 12716 15620
rect 7929 15583 7987 15589
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 13716 15623 13774 15629
rect 13716 15589 13728 15623
rect 13762 15620 13774 15623
rect 14366 15620 14372 15632
rect 13762 15592 14372 15620
rect 13762 15589 13774 15592
rect 13716 15583 13774 15589
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 15930 15580 15936 15632
rect 15988 15580 15994 15632
rect 18316 15623 18374 15629
rect 18316 15589 18328 15623
rect 18362 15620 18374 15623
rect 19150 15620 19156 15632
rect 18362 15592 19156 15620
rect 18362 15589 18374 15592
rect 18316 15583 18374 15589
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 1762 15552 1768 15564
rect 1723 15524 1768 15552
rect 1762 15512 1768 15524
rect 1820 15512 1826 15564
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15552 5595 15555
rect 7006 15552 7012 15564
rect 5583 15524 7012 15552
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 11793 15555 11851 15561
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12434 15552 12440 15564
rect 11839 15524 12440 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 13449 15555 13507 15561
rect 13449 15521 13461 15555
rect 13495 15552 13507 15555
rect 15470 15552 15476 15564
rect 13495 15524 15476 15552
rect 13495 15521 13507 15524
rect 13449 15515 13507 15521
rect 15470 15512 15476 15524
rect 15528 15552 15534 15564
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 15528 15524 15761 15552
rect 15528 15512 15534 15524
rect 15749 15521 15761 15524
rect 15795 15552 15807 15555
rect 15948 15552 15976 15580
rect 15795 15524 15976 15552
rect 16016 15555 16074 15561
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 16016 15521 16028 15555
rect 16062 15552 16074 15555
rect 16482 15552 16488 15564
rect 16062 15524 16488 15552
rect 16062 15521 16074 15524
rect 16016 15515 16074 15521
rect 16482 15512 16488 15524
rect 16540 15512 16546 15564
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 4062 15484 4068 15496
rect 4023 15456 4068 15484
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4890 15484 4896 15496
rect 4851 15456 4896 15484
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 7190 15484 7196 15496
rect 7151 15456 7196 15484
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15484 8263 15487
rect 8662 15484 8668 15496
rect 8251 15456 8668 15484
rect 8251 15453 8263 15456
rect 8205 15447 8263 15453
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10778 15484 10784 15496
rect 10367 15456 10784 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12894 15484 12900 15496
rect 12855 15456 12900 15484
rect 12069 15447 12127 15453
rect 9030 15376 9036 15428
rect 9088 15416 9094 15428
rect 11900 15416 11928 15447
rect 9088 15388 11928 15416
rect 12084 15416 12112 15447
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13127 15456 13308 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 12618 15416 12624 15428
rect 12084 15388 12624 15416
rect 9088 15376 9094 15388
rect 12618 15376 12624 15388
rect 12676 15416 12682 15428
rect 13280 15416 13308 15456
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 18012 15456 18061 15484
rect 18012 15444 18018 15456
rect 18049 15453 18061 15456
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 12676 15388 13308 15416
rect 12676 15376 12682 15388
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 3697 15351 3755 15357
rect 3697 15348 3709 15351
rect 3292 15320 3709 15348
rect 3292 15308 3298 15320
rect 3697 15317 3709 15320
rect 3743 15317 3755 15351
rect 3697 15311 3755 15317
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 5353 15351 5411 15357
rect 5353 15348 5365 15351
rect 4764 15320 5365 15348
rect 4764 15308 4770 15320
rect 5353 15317 5365 15320
rect 5399 15348 5411 15351
rect 5442 15348 5448 15360
rect 5399 15320 5448 15348
rect 5399 15317 5411 15320
rect 5353 15311 5411 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 13280 15348 13308 15388
rect 14829 15351 14887 15357
rect 14829 15348 14841 15351
rect 13280 15320 14841 15348
rect 14829 15317 14841 15320
rect 14875 15317 14887 15351
rect 19426 15348 19432 15360
rect 19387 15320 19432 15348
rect 14829 15311 14887 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2498 15104 2504 15156
rect 2556 15144 2562 15156
rect 2593 15147 2651 15153
rect 2593 15144 2605 15147
rect 2556 15116 2605 15144
rect 2556 15104 2562 15116
rect 2593 15113 2605 15116
rect 2639 15113 2651 15147
rect 6086 15144 6092 15156
rect 6047 15116 6092 15144
rect 2593 15107 2651 15113
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 9950 15144 9956 15156
rect 9907 15116 9956 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13725 15147 13783 15153
rect 13725 15144 13737 15147
rect 12952 15116 13737 15144
rect 12952 15104 12958 15116
rect 13725 15113 13737 15116
rect 13771 15113 13783 15147
rect 13725 15107 13783 15113
rect 15933 15147 15991 15153
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 16114 15144 16120 15156
rect 15979 15116 16120 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 10686 15036 10692 15088
rect 10744 15076 10750 15088
rect 10965 15079 11023 15085
rect 10965 15076 10977 15079
rect 10744 15048 10977 15076
rect 10744 15036 10750 15048
rect 10965 15045 10977 15048
rect 11011 15045 11023 15079
rect 12250 15076 12256 15088
rect 10965 15039 11023 15045
rect 11440 15048 12256 15076
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2682 15008 2688 15020
rect 2179 14980 2688 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3050 15008 3056 15020
rect 3011 14980 3056 15008
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 3234 15008 3240 15020
rect 3195 14980 3240 15008
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 7374 14968 7380 15020
rect 7432 15008 7438 15020
rect 8481 15011 8539 15017
rect 8481 15008 8493 15011
rect 7432 14980 8493 15008
rect 7432 14968 7438 14980
rect 8481 14977 8493 14980
rect 8527 14977 8539 15011
rect 8481 14971 8539 14977
rect 10502 14968 10508 15020
rect 10560 15008 10566 15020
rect 11440 15017 11468 15048
rect 12250 15036 12256 15048
rect 12308 15036 12314 15088
rect 13081 15079 13139 15085
rect 13081 15045 13093 15079
rect 13127 15076 13139 15079
rect 13262 15076 13268 15088
rect 13127 15048 13268 15076
rect 13127 15045 13139 15048
rect 13081 15039 13139 15045
rect 13262 15036 13268 15048
rect 13320 15036 13326 15088
rect 11425 15011 11483 15017
rect 11425 15008 11437 15011
rect 10560 14980 11437 15008
rect 10560 14968 10566 14980
rect 11425 14977 11437 14980
rect 11471 14977 11483 15011
rect 11425 14971 11483 14977
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 1846 14943 1904 14949
rect 1846 14909 1858 14943
rect 1892 14909 1904 14943
rect 1846 14903 1904 14909
rect 2961 14943 3019 14949
rect 2961 14909 2973 14943
rect 3007 14940 3019 14943
rect 4062 14940 4068 14952
rect 3007 14912 4068 14940
rect 3007 14909 3019 14912
rect 2961 14903 3019 14909
rect 1863 14872 1891 14903
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 4709 14943 4767 14949
rect 4709 14940 4721 14943
rect 4396 14912 4721 14940
rect 4396 14900 4402 14912
rect 4709 14909 4721 14912
rect 4755 14940 4767 14943
rect 5534 14940 5540 14952
rect 4755 14912 5540 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 7190 14940 7196 14952
rect 7151 14912 7196 14940
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7466 14900 7472 14952
rect 7524 14940 7530 14952
rect 11333 14943 11391 14949
rect 11333 14940 11345 14943
rect 7524 14912 11345 14940
rect 7524 14900 7530 14912
rect 11333 14909 11345 14912
rect 11379 14909 11391 14943
rect 11333 14903 11391 14909
rect 2682 14872 2688 14884
rect 1863 14844 2688 14872
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 4976 14875 5034 14881
rect 4976 14841 4988 14875
rect 5022 14872 5034 14875
rect 5718 14872 5724 14884
rect 5022 14844 5724 14872
rect 5022 14841 5034 14844
rect 4976 14835 5034 14841
rect 5718 14832 5724 14844
rect 5776 14832 5782 14884
rect 8748 14875 8806 14881
rect 8748 14841 8760 14875
rect 8794 14872 8806 14875
rect 9306 14872 9312 14884
rect 8794 14844 9312 14872
rect 8794 14841 8806 14844
rect 8748 14835 8806 14841
rect 9306 14832 9312 14844
rect 9364 14832 9370 14884
rect 658 14764 664 14816
rect 716 14804 722 14816
rect 10778 14804 10784 14816
rect 716 14776 10784 14804
rect 716 14764 722 14776
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11348 14804 11376 14903
rect 11532 14872 11560 14971
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12492 14980 12537 15008
rect 12492 14968 12498 14980
rect 13998 14968 14004 15020
rect 14056 15008 14062 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 14056 14980 14197 15008
rect 14056 14968 14062 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14366 15008 14372 15020
rect 14327 14980 14372 15008
rect 14185 14971 14243 14977
rect 14366 14968 14372 14980
rect 14424 14968 14430 15020
rect 16482 15008 16488 15020
rect 16443 14980 16488 15008
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 19426 15008 19432 15020
rect 18739 14980 19432 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 13262 14940 13268 14952
rect 13223 14912 13268 14940
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 14458 14940 14464 14952
rect 13964 14912 14464 14940
rect 13964 14900 13970 14912
rect 14458 14900 14464 14912
rect 14516 14940 14522 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 14516 14912 18521 14940
rect 14516 14900 14522 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 11606 14872 11612 14884
rect 11532 14844 11612 14872
rect 11606 14832 11612 14844
rect 11664 14832 11670 14884
rect 16301 14875 16359 14881
rect 16301 14841 16313 14875
rect 16347 14872 16359 14875
rect 16945 14875 17003 14881
rect 16945 14872 16957 14875
rect 16347 14844 16957 14872
rect 16347 14841 16359 14844
rect 16301 14835 16359 14841
rect 16945 14841 16957 14844
rect 16991 14841 17003 14875
rect 18877 14875 18935 14881
rect 18877 14872 18889 14875
rect 16945 14835 17003 14841
rect 18432 14844 18889 14872
rect 18432 14816 18460 14844
rect 18877 14841 18889 14844
rect 18923 14841 18935 14875
rect 18877 14835 18935 14841
rect 13906 14804 13912 14816
rect 11348 14776 13912 14804
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 14090 14804 14096 14816
rect 14051 14776 14096 14804
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 15010 14764 15016 14816
rect 15068 14804 15074 14816
rect 16393 14807 16451 14813
rect 16393 14804 16405 14807
rect 15068 14776 16405 14804
rect 15068 14764 15074 14776
rect 16393 14773 16405 14776
rect 16439 14773 16451 14807
rect 16393 14767 16451 14773
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18230 14804 18236 14816
rect 18095 14776 18236 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 18414 14804 18420 14816
rect 18375 14776 18420 14804
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2958 14600 2964 14612
rect 1627 14572 2964 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 5718 14600 5724 14612
rect 5679 14572 5724 14600
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 9033 14603 9091 14609
rect 5828 14572 7236 14600
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2225 14535 2283 14541
rect 2225 14532 2237 14535
rect 1820 14504 2237 14532
rect 1820 14492 1826 14504
rect 2225 14501 2237 14504
rect 2271 14501 2283 14535
rect 2225 14495 2283 14501
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 5828 14532 5856 14572
rect 3752 14504 5856 14532
rect 6540 14535 6598 14541
rect 3752 14492 3758 14504
rect 6540 14501 6552 14535
rect 6586 14532 6598 14535
rect 7098 14532 7104 14544
rect 6586 14504 7104 14532
rect 6586 14501 6598 14504
rect 6540 14495 6598 14501
rect 7098 14492 7104 14504
rect 7156 14492 7162 14544
rect 7208 14532 7236 14572
rect 9033 14569 9045 14603
rect 9079 14600 9091 14603
rect 10870 14600 10876 14612
rect 9079 14572 10876 14600
rect 9079 14569 9091 14572
rect 9033 14563 9091 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 13998 14600 14004 14612
rect 11020 14572 14004 14600
rect 11020 14560 11026 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 14461 14603 14519 14609
rect 14461 14600 14473 14603
rect 14424 14572 14473 14600
rect 14424 14560 14430 14572
rect 14461 14569 14473 14572
rect 14507 14569 14519 14603
rect 14461 14563 14519 14569
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 16540 14572 16865 14600
rect 16540 14560 16546 14572
rect 16853 14569 16865 14572
rect 16899 14569 16911 14603
rect 18414 14600 18420 14612
rect 16853 14563 16911 14569
rect 17420 14572 18420 14600
rect 10772 14535 10830 14541
rect 7208 14504 9720 14532
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1854 14464 1860 14476
rect 1443 14436 1860 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1854 14424 1860 14436
rect 1912 14424 1918 14476
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14433 2007 14467
rect 1949 14427 2007 14433
rect 1964 14260 1992 14427
rect 2314 14424 2320 14476
rect 2372 14464 2378 14476
rect 4338 14464 4344 14476
rect 2372 14436 4344 14464
rect 2372 14424 2378 14436
rect 4338 14424 4344 14436
rect 4396 14424 4402 14476
rect 4608 14467 4666 14473
rect 4608 14433 4620 14467
rect 4654 14464 4666 14467
rect 6086 14464 6092 14476
rect 4654 14436 6092 14464
rect 4654 14433 4666 14436
rect 4608 14427 4666 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 8938 14464 8944 14476
rect 8899 14436 8944 14464
rect 8938 14424 8944 14436
rect 8996 14424 9002 14476
rect 9692 14464 9720 14504
rect 10772 14501 10784 14535
rect 10818 14532 10830 14535
rect 11606 14532 11612 14544
rect 10818 14504 11612 14532
rect 10818 14501 10830 14504
rect 10772 14495 10830 14501
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 17420 14532 17448 14572
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 11716 14504 17448 14532
rect 17497 14535 17555 14541
rect 11716 14464 11744 14504
rect 17497 14501 17509 14535
rect 17543 14532 17555 14535
rect 17954 14532 17960 14544
rect 17543 14504 17960 14532
rect 17543 14501 17555 14504
rect 17497 14495 17555 14501
rect 17954 14492 17960 14504
rect 18012 14492 18018 14544
rect 18224 14535 18282 14541
rect 18224 14501 18236 14535
rect 18270 14532 18282 14535
rect 19426 14532 19432 14544
rect 18270 14504 19432 14532
rect 18270 14501 18282 14504
rect 18224 14495 18282 14501
rect 19426 14492 19432 14504
rect 19484 14492 19490 14544
rect 9692 14436 11744 14464
rect 12345 14467 12403 14473
rect 12345 14433 12357 14467
rect 12391 14464 12403 14467
rect 12618 14464 12624 14476
rect 12391 14436 12624 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13081 14467 13139 14473
rect 13081 14464 13093 14467
rect 13044 14436 13093 14464
rect 13044 14424 13050 14436
rect 13081 14433 13093 14436
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 13348 14467 13406 14473
rect 13348 14433 13360 14467
rect 13394 14464 13406 14467
rect 13906 14464 13912 14476
rect 13394 14436 13912 14464
rect 13394 14433 13406 14436
rect 13348 14427 13406 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 15470 14464 15476 14476
rect 15431 14436 15476 14464
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 15746 14473 15752 14476
rect 15740 14464 15752 14473
rect 15707 14436 15752 14464
rect 15740 14427 15752 14436
rect 15746 14424 15752 14427
rect 15804 14424 15810 14476
rect 18046 14464 18052 14476
rect 17972 14436 18052 14464
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 6178 14396 6184 14408
rect 5592 14368 6184 14396
rect 5592 14356 5598 14368
rect 6178 14356 6184 14368
rect 6236 14396 6242 14408
rect 6273 14399 6331 14405
rect 6273 14396 6285 14399
rect 6236 14368 6285 14396
rect 6236 14356 6242 14368
rect 6273 14365 6285 14368
rect 6319 14365 6331 14399
rect 6273 14359 6331 14365
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8386 14396 8392 14408
rect 8159 14368 8392 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 10505 14399 10563 14405
rect 9180 14368 9225 14396
rect 9180 14356 9186 14368
rect 10505 14365 10517 14399
rect 10551 14365 10563 14399
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 10505 14359 10563 14365
rect 6914 14260 6920 14272
rect 1964 14232 6920 14260
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 7650 14260 7656 14272
rect 7611 14232 7656 14260
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8570 14260 8576 14272
rect 8531 14232 8576 14260
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 10520 14260 10548 14359
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 13004 14328 13032 14424
rect 17972 14405 18000 14436
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 17957 14399 18015 14405
rect 17957 14365 17969 14399
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 11440 14300 13032 14328
rect 11440 14260 11468 14300
rect 11882 14260 11888 14272
rect 10520 14232 11468 14260
rect 11843 14232 11888 14260
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 14090 14260 14096 14272
rect 12032 14232 14096 14260
rect 12032 14220 12038 14232
rect 14090 14220 14096 14232
rect 14148 14260 14154 14272
rect 17402 14260 17408 14272
rect 14148 14232 17408 14260
rect 14148 14220 14154 14232
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 19337 14263 19395 14269
rect 19337 14260 19349 14263
rect 18748 14232 19349 14260
rect 18748 14220 18754 14232
rect 19337 14229 19349 14232
rect 19383 14229 19395 14263
rect 19337 14223 19395 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2682 14016 2688 14068
rect 2740 14056 2746 14068
rect 4525 14059 4583 14065
rect 4525 14056 4537 14059
rect 2740 14028 4537 14056
rect 2740 14016 2746 14028
rect 4525 14025 4537 14028
rect 4571 14025 4583 14059
rect 9306 14056 9312 14068
rect 9267 14028 9312 14056
rect 4525 14019 4583 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 12618 14056 12624 14068
rect 12579 14028 12624 14056
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 13262 14016 13268 14068
rect 13320 14016 13326 14068
rect 15010 14056 15016 14068
rect 14971 14028 15016 14056
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 15746 14056 15752 14068
rect 15659 14028 15752 14056
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 5000 13960 5549 13988
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2314 13880 2320 13932
rect 2372 13920 2378 13932
rect 5000 13929 5028 13960
rect 5537 13957 5549 13960
rect 5583 13957 5595 13991
rect 5537 13951 5595 13957
rect 5810 13948 5816 14000
rect 5868 13988 5874 14000
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 5868 13960 6837 13988
rect 5868 13948 5874 13960
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 6825 13951 6883 13957
rect 7374 13948 7380 14000
rect 7432 13988 7438 14000
rect 7432 13960 7972 13988
rect 7432 13948 7438 13960
rect 2409 13923 2467 13929
rect 2409 13920 2421 13923
rect 2372 13892 2421 13920
rect 2372 13880 2378 13892
rect 2409 13889 2421 13892
rect 2455 13889 2467 13923
rect 2409 13883 2467 13889
rect 4985 13923 5043 13929
rect 4985 13889 4997 13923
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5169 13923 5227 13929
rect 5169 13889 5181 13923
rect 5215 13920 5227 13923
rect 5718 13920 5724 13932
rect 5215 13892 5724 13920
rect 5215 13889 5227 13892
rect 5169 13883 5227 13889
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 6086 13920 6092 13932
rect 6047 13892 6092 13920
rect 6086 13880 6092 13892
rect 6144 13880 6150 13932
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7650 13920 7656 13932
rect 7515 13892 7656 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 7944 13929 7972 13960
rect 10778 13948 10784 14000
rect 10836 13988 10842 14000
rect 10836 13960 11468 13988
rect 10836 13948 10842 13960
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 11146 13920 11152 13932
rect 10551 13892 11152 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 11440 13929 11468 13960
rect 11606 13948 11612 14000
rect 11664 13948 11670 14000
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13988 12127 13991
rect 13280 13988 13308 14016
rect 12115 13960 13308 13988
rect 12115 13957 12127 13960
rect 12069 13951 12127 13957
rect 11425 13923 11483 13929
rect 11425 13889 11437 13923
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13920 11575 13923
rect 11624 13920 11652 13948
rect 13265 13923 13323 13929
rect 11563 13892 12388 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2676 13855 2734 13861
rect 1719 13824 2360 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2332 13784 2360 13824
rect 2676 13821 2688 13855
rect 2722 13852 2734 13855
rect 3234 13852 3240 13864
rect 2722 13824 3240 13852
rect 2722 13821 2734 13824
rect 2676 13815 2734 13821
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 5258 13852 5264 13864
rect 3344 13824 5264 13852
rect 3344 13784 3372 13824
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5997 13855 6055 13861
rect 5997 13821 6009 13855
rect 6043 13852 6055 13855
rect 6822 13852 6828 13864
rect 6043 13824 6828 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7285 13855 7343 13861
rect 7285 13821 7297 13855
rect 7331 13852 7343 13855
rect 7742 13852 7748 13864
rect 7331 13824 7748 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 8196 13855 8254 13861
rect 8196 13821 8208 13855
rect 8242 13852 8254 13855
rect 9122 13852 9128 13864
rect 8242 13824 9128 13852
rect 8242 13821 8254 13824
rect 8196 13815 8254 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13852 10287 13855
rect 11606 13852 11612 13864
rect 10275 13824 11612 13852
rect 10275 13821 10287 13824
rect 10229 13815 10287 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 12250 13852 12256 13864
rect 12211 13824 12256 13852
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12360 13852 12388 13892
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13906 13920 13912 13932
rect 13311 13892 13912 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15672 13929 15700 14028
rect 15746 14016 15752 14028
rect 15804 14056 15810 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 15804 14028 17417 14056
rect 15804 14016 15810 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 17405 14019 17463 14025
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18782 14056 18788 14068
rect 18095 14028 18788 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 15160 13892 15485 13920
rect 15160 13880 15166 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13889 15715 13923
rect 18506 13920 18512 13932
rect 18467 13892 18512 13920
rect 15657 13883 15715 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 18690 13920 18696 13932
rect 18651 13892 18696 13920
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 14550 13852 14556 13864
rect 12360 13824 14556 13852
rect 14550 13812 14556 13824
rect 14608 13812 14614 13864
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 17678 13852 17684 13864
rect 16071 13824 17684 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 4890 13784 4896 13796
rect 2332 13756 3372 13784
rect 4851 13756 4896 13784
rect 4890 13744 4896 13756
rect 4948 13744 4954 13796
rect 4982 13744 4988 13796
rect 5040 13784 5046 13796
rect 5350 13784 5356 13796
rect 5040 13756 5356 13784
rect 5040 13744 5046 13756
rect 5350 13744 5356 13756
rect 5408 13784 5414 13796
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 5408 13756 7205 13784
rect 5408 13744 5414 13756
rect 7193 13753 7205 13756
rect 7239 13753 7251 13787
rect 7193 13747 7251 13753
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 12802 13784 12808 13796
rect 7432 13756 12808 13784
rect 7432 13744 7438 13756
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 16040 13784 16068 13815
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 15344 13756 16068 13784
rect 16292 13787 16350 13793
rect 15344 13744 15350 13756
rect 16292 13753 16304 13787
rect 16338 13784 16350 13787
rect 16390 13784 16396 13796
rect 16338 13756 16396 13784
rect 16338 13753 16350 13756
rect 16292 13747 16350 13753
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 18417 13787 18475 13793
rect 18417 13784 18429 13787
rect 18012 13756 18429 13784
rect 18012 13744 18018 13756
rect 18417 13753 18429 13756
rect 18463 13753 18475 13787
rect 18417 13747 18475 13753
rect 3694 13676 3700 13728
rect 3752 13716 3758 13728
rect 3789 13719 3847 13725
rect 3789 13716 3801 13719
rect 3752 13688 3801 13716
rect 3752 13676 3758 13688
rect 3789 13685 3801 13688
rect 3835 13685 3847 13719
rect 3789 13679 3847 13685
rect 5905 13719 5963 13725
rect 5905 13685 5917 13719
rect 5951 13716 5963 13719
rect 8938 13716 8944 13728
rect 5951 13688 8944 13716
rect 5951 13685 5963 13688
rect 5905 13679 5963 13685
rect 8938 13676 8944 13688
rect 8996 13676 9002 13728
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 11146 13716 11152 13728
rect 11011 13688 11152 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11333 13719 11391 13725
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 11974 13716 11980 13728
rect 11379 13688 11980 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12986 13716 12992 13728
rect 12947 13688 12992 13716
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13136 13688 13181 13716
rect 13136 13676 13142 13688
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 14332 13688 15393 13716
rect 14332 13676 14338 13688
rect 15381 13685 15393 13688
rect 15427 13685 15439 13719
rect 15381 13679 15439 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1394 13472 1400 13524
rect 1452 13512 1458 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 1452 13484 1593 13512
rect 1452 13472 1458 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 2685 13515 2743 13521
rect 2685 13481 2697 13515
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 3145 13515 3203 13521
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3191 13484 4077 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1949 13379 2007 13385
rect 1949 13345 1961 13379
rect 1995 13376 2007 13379
rect 2700 13376 2728 13475
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4212 13484 4537 13512
rect 4212 13472 4218 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 5258 13512 5264 13524
rect 5219 13484 5264 13512
rect 4525 13475 4583 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 5810 13512 5816 13524
rect 5767 13484 5816 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 6972 13484 8033 13512
rect 6972 13472 6978 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8021 13475 8079 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8570 13512 8576 13524
rect 8527 13484 8576 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 13906 13512 13912 13524
rect 13867 13484 13912 13512
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 14182 13472 14188 13524
rect 14240 13512 14246 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14240 13484 14565 13512
rect 14240 13472 14246 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 14553 13475 14611 13481
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 15102 13512 15108 13524
rect 14691 13484 15108 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 15838 13512 15844 13524
rect 15795 13484 15844 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 4982 13444 4988 13456
rect 4479 13416 4988 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 4982 13404 4988 13416
rect 5040 13404 5046 13456
rect 6540 13447 6598 13453
rect 5092 13416 6316 13444
rect 1995 13348 2728 13376
rect 3053 13379 3111 13385
rect 1995 13345 2007 13348
rect 1949 13339 2007 13345
rect 3053 13345 3065 13379
rect 3099 13376 3111 13379
rect 3510 13376 3516 13388
rect 3099 13348 3516 13376
rect 3099 13345 3111 13348
rect 3053 13339 3111 13345
rect 1412 13308 1440 13339
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 5092 13376 5120 13416
rect 4120 13348 5120 13376
rect 5629 13379 5687 13385
rect 4120 13336 4126 13348
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 6178 13376 6184 13388
rect 5675 13348 6184 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 6288 13376 6316 13416
rect 6540 13413 6552 13447
rect 6586 13444 6598 13447
rect 7650 13444 7656 13456
rect 6586 13416 7656 13444
rect 6586 13413 6598 13416
rect 6540 13407 6598 13413
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 16574 13444 16580 13456
rect 12728 13416 16580 13444
rect 7374 13376 7380 13388
rect 6288 13348 7380 13376
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 12728 13376 12756 13416
rect 16574 13404 16580 13416
rect 16632 13404 16638 13456
rect 17948 13447 18006 13453
rect 17948 13413 17960 13447
rect 17994 13444 18006 13447
rect 18690 13444 18696 13456
rect 17994 13416 18696 13444
rect 17994 13413 18006 13416
rect 17948 13407 18006 13413
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 12802 13385 12808 13388
rect 10284 13348 12756 13376
rect 10284 13336 10290 13348
rect 12796 13339 12808 13385
rect 12860 13376 12866 13388
rect 16117 13379 16175 13385
rect 12860 13348 12896 13376
rect 12802 13336 12808 13339
rect 12860 13336 12866 13348
rect 16117 13345 16129 13379
rect 16163 13376 16175 13379
rect 16761 13379 16819 13385
rect 16761 13376 16773 13379
rect 16163 13348 16773 13376
rect 16163 13345 16175 13348
rect 16117 13339 16175 13345
rect 16761 13345 16773 13348
rect 16807 13345 16819 13379
rect 17678 13376 17684 13388
rect 17639 13348 17684 13376
rect 16761 13339 16819 13345
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 1412 13280 2145 13308
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13308 3387 13311
rect 4246 13308 4252 13320
rect 3375 13280 4252 13308
rect 3375 13277 3387 13280
rect 3329 13271 3387 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 3694 13200 3700 13252
rect 3752 13240 3758 13252
rect 4632 13240 4660 13271
rect 3752 13212 4660 13240
rect 3752 13200 3758 13212
rect 5920 13172 5948 13271
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6144 13280 6285 13308
rect 6144 13268 6150 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 8665 13311 8723 13317
rect 8665 13277 8677 13311
rect 8711 13308 8723 13311
rect 9306 13308 9312 13320
rect 8711 13280 9312 13308
rect 8711 13277 8723 13280
rect 8665 13271 8723 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 10042 13308 10048 13320
rect 9723 13280 10048 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 12526 13308 12532 13320
rect 12487 13280 12532 13308
rect 12526 13268 12532 13280
rect 12584 13268 12590 13320
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15010 13308 15016 13320
rect 14875 13280 15016 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13277 16267 13311
rect 16390 13308 16396 13320
rect 16351 13280 16396 13308
rect 16209 13271 16267 13277
rect 16224 13240 16252 13271
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 16942 13240 16948 13252
rect 16224 13212 16948 13240
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 6086 13172 6092 13184
rect 5920 13144 6092 13172
rect 6086 13132 6092 13144
rect 6144 13172 6150 13184
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 6144 13144 7665 13172
rect 6144 13132 6150 13144
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 7653 13135 7711 13141
rect 8478 13132 8484 13184
rect 8536 13172 8542 13184
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 8536 13144 11437 13172
rect 8536 13132 8542 13144
rect 11425 13141 11437 13144
rect 11471 13172 11483 13175
rect 12250 13172 12256 13184
rect 11471 13144 12256 13172
rect 11471 13141 11483 13144
rect 11425 13135 11483 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 14182 13172 14188 13184
rect 14143 13144 14188 13172
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 19058 13172 19064 13184
rect 19019 13144 19064 13172
rect 19058 13132 19064 13144
rect 19116 13132 19122 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 2222 12928 2228 12980
rect 2280 12968 2286 12980
rect 2501 12971 2559 12977
rect 2501 12968 2513 12971
rect 2280 12940 2513 12968
rect 2280 12928 2286 12940
rect 2501 12937 2513 12940
rect 2547 12937 2559 12971
rect 2501 12931 2559 12937
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7558 12968 7564 12980
rect 7248 12940 7564 12968
rect 7248 12928 7254 12940
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 10226 12968 10232 12980
rect 7668 12940 10232 12968
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 2774 12900 2780 12912
rect 1995 12872 2780 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 4246 12860 4252 12912
rect 4304 12900 4310 12912
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 4304 12872 4629 12900
rect 4304 12860 4310 12872
rect 4617 12869 4629 12872
rect 4663 12900 4675 12903
rect 7668 12900 7696 12940
rect 10226 12928 10232 12940
rect 10284 12928 10290 12980
rect 10689 12971 10747 12977
rect 10689 12937 10701 12971
rect 10735 12968 10747 12971
rect 10870 12968 10876 12980
rect 10735 12940 10876 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12968 11575 12971
rect 11606 12968 11612 12980
rect 11563 12940 11612 12968
rect 11563 12937 11575 12940
rect 11517 12931 11575 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 13078 12968 13084 12980
rect 12483 12940 13084 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 14369 12971 14427 12977
rect 14369 12968 14381 12971
rect 13320 12940 14381 12968
rect 13320 12928 13326 12940
rect 14369 12937 14381 12940
rect 14415 12937 14427 12971
rect 16022 12968 16028 12980
rect 14369 12931 14427 12937
rect 14476 12940 16028 12968
rect 10594 12900 10600 12912
rect 4663 12872 7696 12900
rect 10555 12872 10600 12900
rect 4663 12869 4675 12872
rect 4617 12863 4675 12869
rect 10594 12860 10600 12872
rect 10652 12860 10658 12912
rect 11882 12900 11888 12912
rect 11339 12872 11888 12900
rect 11339 12844 11367 12872
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 14476 12900 14504 12940
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 16448 12940 16681 12968
rect 16448 12928 16454 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 16942 12968 16948 12980
rect 16903 12940 16948 12968
rect 16669 12931 16727 12937
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18598 12968 18604 12980
rect 18095 12940 18604 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 13872 12872 14504 12900
rect 13872 12860 13878 12872
rect 6178 12832 6184 12844
rect 6139 12804 6184 12832
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 9030 12832 9036 12844
rect 6512 12804 9036 12832
rect 6512 12792 6518 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11204 12804 11249 12832
rect 11204 12792 11210 12804
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11388 12804 11481 12832
rect 11388 12792 11394 12804
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 12032 12804 12081 12832
rect 12032 12792 12038 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12860 12804 13001 12832
rect 12860 12792 12866 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12832 14151 12835
rect 15010 12832 15016 12844
rect 14139 12804 15016 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15286 12832 15292 12844
rect 15247 12804 15292 12832
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 16724 12804 17509 12832
rect 16724 12792 16730 12804
rect 17497 12801 17509 12804
rect 17543 12801 17555 12835
rect 18690 12832 18696 12844
rect 18651 12804 18696 12832
rect 17497 12795 17555 12801
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2317 12767 2375 12773
rect 2317 12733 2329 12767
rect 2363 12764 2375 12767
rect 3050 12764 3056 12776
rect 2363 12736 3056 12764
rect 2363 12733 2375 12736
rect 2317 12727 2375 12733
rect 3050 12724 3056 12736
rect 3108 12724 3114 12776
rect 3237 12767 3295 12773
rect 3237 12733 3249 12767
rect 3283 12764 3295 12767
rect 3786 12764 3792 12776
rect 3283 12736 3792 12764
rect 3283 12733 3295 12736
rect 3237 12727 3295 12733
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 8478 12764 8484 12776
rect 7791 12736 8484 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8478 12724 8484 12736
rect 8536 12724 8542 12776
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 8628 12736 9229 12764
rect 8628 12724 8634 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 9484 12767 9542 12773
rect 9484 12733 9496 12767
rect 9530 12764 9542 12767
rect 9530 12736 9628 12764
rect 9530 12733 9542 12736
rect 9484 12727 9542 12733
rect 3504 12699 3562 12705
rect 3504 12665 3516 12699
rect 3550 12696 3562 12699
rect 3694 12696 3700 12708
rect 3550 12668 3700 12696
rect 3550 12665 3562 12668
rect 3504 12659 3562 12665
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 9600 12696 9628 12736
rect 11606 12724 11612 12776
rect 11664 12764 11670 12776
rect 13909 12767 13967 12773
rect 13909 12764 13921 12767
rect 11664 12736 13921 12764
rect 11664 12724 11670 12736
rect 13909 12733 13921 12736
rect 13955 12764 13967 12767
rect 14369 12767 14427 12773
rect 13955 12736 14320 12764
rect 13955 12733 13967 12736
rect 13909 12727 13967 12733
rect 10318 12696 10324 12708
rect 9600 12668 10324 12696
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 10686 12656 10692 12708
rect 10744 12696 10750 12708
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 10744 12668 11069 12696
rect 10744 12656 10750 12668
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11057 12659 11115 12665
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 11977 12699 12035 12705
rect 11977 12696 11989 12699
rect 11204 12668 11989 12696
rect 11204 12656 11210 12668
rect 11977 12665 11989 12668
rect 12023 12665 12035 12699
rect 11977 12659 12035 12665
rect 12805 12699 12863 12705
rect 12805 12665 12817 12699
rect 12851 12696 12863 12699
rect 14182 12696 14188 12708
rect 12851 12668 14188 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 14292 12696 14320 12736
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 14645 12767 14703 12773
rect 14645 12764 14657 12767
rect 14415 12736 14657 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 14645 12733 14657 12736
rect 14691 12733 14703 12767
rect 14645 12727 14703 12733
rect 15556 12767 15614 12773
rect 15556 12733 15568 12767
rect 15602 12764 15614 12767
rect 16684 12764 16712 12792
rect 17402 12764 17408 12776
rect 15602 12736 16712 12764
rect 17363 12736 17408 12764
rect 15602 12733 15614 12736
rect 15556 12727 15614 12733
rect 17402 12724 17408 12736
rect 17460 12724 17466 12776
rect 15654 12696 15660 12708
rect 14292 12668 15660 12696
rect 15654 12656 15660 12668
rect 15712 12696 15718 12708
rect 17126 12696 17132 12708
rect 15712 12668 17132 12696
rect 15712 12656 15718 12668
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 17954 12656 17960 12708
rect 18012 12696 18018 12708
rect 18417 12699 18475 12705
rect 18417 12696 18429 12699
rect 18012 12668 18429 12696
rect 18012 12656 18018 12668
rect 18417 12665 18429 12668
rect 18463 12665 18475 12699
rect 18417 12659 18475 12665
rect 11882 12628 11888 12640
rect 11843 12600 11888 12628
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 12943 12600 13461 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13814 12628 13820 12640
rect 13775 12600 13820 12628
rect 13449 12591 13507 12597
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 14458 12628 14464 12640
rect 14419 12600 14464 12628
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 14550 12588 14556 12640
rect 14608 12628 14614 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 14608 12600 17325 12628
rect 14608 12588 14614 12600
rect 17313 12597 17325 12600
rect 17359 12597 17371 12631
rect 17313 12591 17371 12597
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 18564 12600 18609 12628
rect 18564 12588 18570 12600
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 3510 12424 3516 12436
rect 3471 12396 3516 12424
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 5629 12427 5687 12433
rect 3620 12396 5304 12424
rect 1762 12316 1768 12368
rect 1820 12356 1826 12368
rect 2317 12359 2375 12365
rect 2317 12356 2329 12359
rect 1820 12328 2329 12356
rect 1820 12316 1826 12328
rect 2317 12325 2329 12328
rect 2363 12325 2375 12359
rect 3050 12356 3056 12368
rect 3011 12328 3056 12356
rect 2317 12319 2375 12325
rect 3050 12316 3056 12328
rect 3108 12316 3114 12368
rect 3234 12316 3240 12368
rect 3292 12356 3298 12368
rect 3620 12356 3648 12396
rect 3292 12328 3648 12356
rect 3292 12316 3298 12328
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 5276 12356 5304 12396
rect 5629 12393 5641 12427
rect 5675 12424 5687 12427
rect 5994 12424 6000 12436
rect 5675 12396 6000 12424
rect 5675 12393 5687 12396
rect 5629 12387 5687 12393
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 7650 12424 7656 12436
rect 6104 12396 7656 12424
rect 6104 12356 6132 12396
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 9122 12424 9128 12436
rect 9083 12396 9128 12424
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 10042 12424 10048 12436
rect 10003 12396 10048 12424
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 12986 12384 12992 12436
rect 13044 12424 13050 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13044 12396 13645 12424
rect 13044 12384 13050 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15286 12424 15292 12436
rect 14967 12396 15292 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 16666 12424 16672 12436
rect 16627 12396 16672 12424
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 18506 12424 18512 12436
rect 17635 12396 18512 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 6178 12365 6184 12368
rect 4120 12328 5212 12356
rect 5276 12328 6132 12356
rect 4120 12316 4126 12328
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2056 12084 2084 12251
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 4516 12291 4574 12297
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 4516 12257 4528 12291
rect 4562 12288 4574 12291
rect 5074 12288 5080 12300
rect 4562 12260 5080 12288
rect 4562 12257 4574 12260
rect 4516 12251 4574 12257
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5184 12288 5212 12328
rect 6172 12319 6184 12365
rect 6236 12356 6242 12368
rect 10137 12359 10195 12365
rect 10137 12356 10149 12359
rect 6236 12328 6272 12356
rect 6472 12328 10149 12356
rect 6178 12316 6184 12319
rect 6236 12316 6242 12328
rect 6472 12288 6500 12328
rect 10137 12325 10149 12328
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 12244 12359 12302 12365
rect 12244 12325 12256 12359
rect 12290 12356 12302 12359
rect 14182 12356 14188 12368
rect 12290 12328 14188 12356
rect 12290 12325 12302 12328
rect 12244 12319 12302 12325
rect 14182 12316 14188 12328
rect 14240 12316 14246 12368
rect 15556 12359 15614 12365
rect 15556 12325 15568 12359
rect 15602 12356 15614 12359
rect 15746 12356 15752 12368
rect 15602 12328 15752 12356
rect 15602 12325 15614 12328
rect 15556 12319 15614 12325
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 17957 12359 18015 12365
rect 17957 12356 17969 12359
rect 17828 12328 17969 12356
rect 17828 12316 17834 12328
rect 17957 12325 17969 12328
rect 18003 12325 18015 12359
rect 17957 12319 18015 12325
rect 5184 12260 6500 12288
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 8001 12291 8059 12297
rect 8001 12288 8013 12291
rect 7524 12260 8013 12288
rect 7524 12248 7530 12260
rect 8001 12257 8013 12260
rect 8047 12257 8059 12291
rect 8001 12251 8059 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12526 12288 12532 12300
rect 12023 12260 12532 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12526 12248 12532 12260
rect 12584 12288 12590 12300
rect 13262 12288 13268 12300
rect 12584 12260 13268 12288
rect 12584 12248 12590 12260
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 14001 12291 14059 12297
rect 14001 12288 14013 12291
rect 13504 12260 14013 12288
rect 13504 12248 13510 12260
rect 14001 12257 14013 12260
rect 14047 12257 14059 12291
rect 14001 12251 14059 12257
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 15102 12288 15108 12300
rect 14516 12260 15108 12288
rect 14516 12248 14522 12260
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 15286 12288 15292 12300
rect 15199 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12288 15350 12300
rect 15930 12288 15936 12300
rect 15344 12260 15936 12288
rect 15344 12248 15350 12260
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 18049 12291 18107 12297
rect 18049 12288 18061 12291
rect 17184 12260 18061 12288
rect 17184 12248 17190 12260
rect 18049 12257 18061 12260
rect 18095 12257 18107 12291
rect 18049 12251 18107 12257
rect 3602 12180 3608 12232
rect 3660 12220 3666 12232
rect 3786 12220 3792 12232
rect 3660 12192 3792 12220
rect 3660 12180 3666 12192
rect 3786 12180 3792 12192
rect 3844 12220 3850 12232
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 3844 12192 4261 12220
rect 3844 12180 3850 12192
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 5810 12180 5816 12232
rect 5868 12220 5874 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5868 12192 5917 12220
rect 5868 12180 5874 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 10318 12220 10324 12232
rect 10231 12192 10324 12220
rect 7745 12183 7803 12189
rect 4890 12084 4896 12096
rect 2056 12056 4896 12084
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 7285 12087 7343 12093
rect 7285 12084 7297 12087
rect 6604 12056 7297 12084
rect 6604 12044 6610 12056
rect 7285 12053 7297 12056
rect 7331 12053 7343 12087
rect 7285 12047 7343 12053
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7760 12084 7788 12183
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 11330 12220 11336 12232
rect 10376 12192 11336 12220
rect 10376 12180 10382 12192
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 14090 12220 14096 12232
rect 14051 12192 14096 12220
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12189 14243 12223
rect 14185 12183 14243 12189
rect 18233 12223 18291 12229
rect 18233 12189 18245 12223
rect 18279 12220 18291 12223
rect 18506 12220 18512 12232
rect 18279 12192 18512 12220
rect 18279 12189 18291 12192
rect 18233 12183 18291 12189
rect 9677 12155 9735 12161
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 11882 12152 11888 12164
rect 9723 12124 11888 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 14200 12152 14228 12183
rect 18506 12180 18512 12192
rect 18564 12220 18570 12232
rect 19058 12220 19064 12232
rect 18564 12192 19064 12220
rect 18564 12180 18570 12192
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 13372 12124 14228 12152
rect 8478 12084 8484 12096
rect 7432 12056 8484 12084
rect 7432 12044 7438 12056
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13372 12093 13400 12124
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 12952 12056 13369 12084
rect 12952 12044 12958 12056
rect 13357 12053 13369 12056
rect 13403 12053 13415 12087
rect 13357 12047 13415 12053
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 3142 11880 3148 11892
rect 2915 11852 3148 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 5132 11852 5181 11880
rect 5132 11840 5138 11852
rect 5169 11849 5181 11852
rect 5215 11849 5227 11883
rect 7558 11880 7564 11892
rect 5169 11843 5227 11849
rect 7208 11852 7564 11880
rect 4890 11772 4896 11824
rect 4948 11812 4954 11824
rect 6822 11812 6828 11824
rect 4948 11784 6828 11812
rect 4948 11772 4954 11784
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 1964 11716 3924 11744
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 1964 11685 1992 11716
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2225 11679 2283 11685
rect 2225 11645 2237 11679
rect 2271 11676 2283 11679
rect 2685 11679 2743 11685
rect 2685 11676 2697 11679
rect 2271 11648 2697 11676
rect 2271 11645 2283 11648
rect 2225 11639 2283 11645
rect 2685 11645 2697 11648
rect 2731 11645 2743 11679
rect 2685 11639 2743 11645
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3789 11679 3847 11685
rect 3789 11676 3801 11679
rect 3660 11648 3801 11676
rect 3660 11636 3666 11648
rect 3789 11645 3801 11648
rect 3835 11645 3847 11679
rect 3789 11639 3847 11645
rect 3896 11608 3924 11716
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 6236 11716 6377 11744
rect 6236 11704 6242 11716
rect 6365 11713 6377 11716
rect 6411 11744 6423 11747
rect 6546 11744 6552 11756
rect 6411 11716 6552 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 6546 11704 6552 11716
rect 6604 11704 6610 11756
rect 4056 11679 4114 11685
rect 4056 11645 4068 11679
rect 4102 11676 4114 11679
rect 6196 11676 6224 11704
rect 7208 11685 7236 11852
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 12437 11883 12495 11889
rect 7708 11852 10732 11880
rect 7708 11840 7714 11852
rect 10704 11812 10732 11852
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 14090 11880 14096 11892
rect 12483 11852 14096 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 15010 11880 15016 11892
rect 14240 11852 15016 11880
rect 14240 11840 14246 11852
rect 15010 11840 15016 11852
rect 15068 11880 15074 11892
rect 16945 11883 17003 11889
rect 15068 11852 15332 11880
rect 15068 11840 15074 11852
rect 15304 11812 15332 11852
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 17954 11880 17960 11892
rect 16991 11852 17960 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 19981 11883 20039 11889
rect 19981 11880 19993 11883
rect 18064 11852 19993 11880
rect 18064 11812 18092 11852
rect 19981 11849 19993 11852
rect 20027 11849 20039 11883
rect 19981 11843 20039 11849
rect 10704 11784 14412 11812
rect 15304 11784 18092 11812
rect 7374 11744 7380 11756
rect 7335 11716 7380 11744
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 8628 11716 9781 11744
rect 8628 11704 8634 11716
rect 9769 11713 9781 11716
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13446 11744 13452 11756
rect 13127 11716 13216 11744
rect 13407 11716 13452 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 4102 11648 6224 11676
rect 7193 11679 7251 11685
rect 4102 11645 4114 11648
rect 4056 11639 4114 11645
rect 7193 11645 7205 11679
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7926 11636 7932 11688
rect 7984 11676 7990 11688
rect 9858 11676 9864 11688
rect 7984 11648 9864 11676
rect 7984 11636 7990 11648
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 10036 11679 10094 11685
rect 10036 11645 10048 11679
rect 10082 11676 10094 11679
rect 10594 11676 10600 11688
rect 10082 11648 10600 11676
rect 10082 11645 10094 11648
rect 10036 11639 10094 11645
rect 10594 11636 10600 11648
rect 10652 11636 10658 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 12066 11676 12072 11688
rect 11112 11648 12072 11676
rect 11112 11636 11118 11648
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 4798 11608 4804 11620
rect 3896 11580 4804 11608
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 6086 11608 6092 11620
rect 6047 11580 6092 11608
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 6181 11611 6239 11617
rect 6181 11577 6193 11611
rect 6227 11608 6239 11611
rect 6270 11608 6276 11620
rect 6227 11580 6276 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 7644 11611 7702 11617
rect 7644 11577 7656 11611
rect 7690 11608 7702 11611
rect 7742 11608 7748 11620
rect 7690 11580 7748 11608
rect 7690 11577 7702 11580
rect 7644 11571 7702 11577
rect 7742 11568 7748 11580
rect 7800 11568 7806 11620
rect 11606 11568 11612 11620
rect 11664 11608 11670 11620
rect 13188 11608 13216 11716
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 14384 11744 14412 11784
rect 17589 11747 17647 11753
rect 14384 11716 14504 11744
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 13320 11648 14381 11676
rect 13320 11636 13326 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 14476 11676 14504 11716
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 17954 11744 17960 11756
rect 17635 11716 17960 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 17954 11704 17960 11716
rect 18012 11744 18018 11756
rect 18506 11744 18512 11756
rect 18012 11716 18512 11744
rect 18012 11704 18018 11716
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 14476 11648 17417 11676
rect 14369 11639 14427 11645
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 18598 11676 18604 11688
rect 18559 11648 18604 11676
rect 17405 11639 17463 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 14182 11608 14188 11620
rect 11664 11580 12940 11608
rect 13188 11580 14188 11608
rect 11664 11568 11670 11580
rect 5718 11540 5724 11552
rect 5679 11512 5724 11540
rect 5718 11500 5724 11512
rect 5776 11500 5782 11552
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8757 11543 8815 11549
rect 8757 11540 8769 11543
rect 7524 11512 8769 11540
rect 7524 11500 7530 11512
rect 8757 11509 8769 11512
rect 8803 11509 8815 11543
rect 8757 11503 8815 11509
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 10836 11512 11161 11540
rect 10836 11500 10842 11512
rect 11149 11509 11161 11512
rect 11195 11509 11207 11543
rect 11149 11503 11207 11509
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 12912 11549 12940 11580
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 14550 11568 14556 11620
rect 14608 11617 14614 11620
rect 18874 11617 18880 11620
rect 14608 11611 14672 11617
rect 14608 11577 14626 11611
rect 14660 11577 14672 11611
rect 17313 11611 17371 11617
rect 14608 11571 14672 11577
rect 15304 11580 16804 11608
rect 14608 11568 14614 11571
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12676 11512 12817 11540
rect 12676 11500 12682 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12897 11543 12955 11549
rect 12897 11509 12909 11543
rect 12943 11540 12955 11543
rect 15304 11540 15332 11580
rect 15746 11540 15752 11552
rect 12943 11512 15332 11540
rect 15707 11512 15752 11540
rect 12943 11509 12955 11512
rect 12897 11503 12955 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16666 11540 16672 11552
rect 16071 11512 16672 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16776 11540 16804 11580
rect 17313 11577 17325 11611
rect 17359 11608 17371 11611
rect 18049 11611 18107 11617
rect 18049 11608 18061 11611
rect 17359 11580 18061 11608
rect 17359 11577 17371 11580
rect 17313 11571 17371 11577
rect 18049 11577 18061 11580
rect 18095 11577 18107 11611
rect 18868 11608 18880 11617
rect 18835 11580 18880 11608
rect 18049 11571 18107 11577
rect 18868 11571 18880 11580
rect 18874 11568 18880 11571
rect 18932 11568 18938 11620
rect 17770 11540 17776 11552
rect 16776 11512 17776 11540
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 2832 11308 4537 11336
rect 2832 11296 2838 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 4893 11339 4951 11345
rect 4893 11305 4905 11339
rect 4939 11336 4951 11339
rect 5537 11339 5595 11345
rect 5537 11336 5549 11339
rect 4939 11308 5549 11336
rect 4939 11305 4951 11308
rect 4893 11299 4951 11305
rect 5537 11305 5549 11308
rect 5583 11305 5595 11339
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 5537 11299 5595 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7285 11339 7343 11345
rect 7285 11305 7297 11339
rect 7331 11336 7343 11339
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 7331 11308 7849 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 7837 11299 7895 11305
rect 10229 11339 10287 11345
rect 10229 11305 10241 11339
rect 10275 11336 10287 11339
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 10275 11308 12633 11336
rect 10275 11305 10287 11308
rect 10229 11299 10287 11305
rect 12621 11305 12633 11308
rect 12667 11305 12679 11339
rect 12621 11299 12679 11305
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13354 11336 13360 11348
rect 13311 11308 13360 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 15749 11339 15807 11345
rect 15749 11305 15761 11339
rect 15795 11336 15807 11339
rect 16022 11336 16028 11348
rect 15795 11308 16028 11336
rect 15795 11305 15807 11308
rect 15749 11299 15807 11305
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11305 16359 11339
rect 16666 11336 16672 11348
rect 16627 11308 16672 11336
rect 16301 11299 16359 11305
rect 4985 11271 5043 11277
rect 4985 11237 4997 11271
rect 5031 11268 5043 11271
rect 5718 11268 5724 11280
rect 5031 11240 5724 11268
rect 5031 11237 5043 11240
rect 4985 11231 5043 11237
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 6730 11228 6736 11280
rect 6788 11268 6794 11280
rect 11146 11268 11152 11280
rect 6788 11240 11152 11268
rect 6788 11228 6794 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 12250 11228 12256 11280
rect 12308 11228 12314 11280
rect 15562 11228 15568 11280
rect 15620 11268 15626 11280
rect 16316 11268 16344 11299
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 15620 11240 16344 11268
rect 17580 11271 17638 11277
rect 15620 11228 15626 11240
rect 17580 11237 17592 11271
rect 17626 11268 17638 11271
rect 17954 11268 17960 11280
rect 17626 11240 17960 11268
rect 17626 11237 17638 11240
rect 17580 11231 17638 11237
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 2406 11200 2412 11212
rect 2367 11172 2412 11200
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5905 11203 5963 11209
rect 5905 11200 5917 11203
rect 5592 11172 5917 11200
rect 5592 11160 5598 11172
rect 5905 11169 5917 11172
rect 5951 11169 5963 11203
rect 7190 11200 7196 11212
rect 7151 11172 7196 11200
rect 5905 11163 5963 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 7300 11172 8217 11200
rect 2498 11132 2504 11144
rect 2459 11104 2504 11132
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2590 11092 2596 11144
rect 2648 11132 2654 11144
rect 5074 11132 5080 11144
rect 2648 11104 2693 11132
rect 5035 11104 5080 11132
rect 2648 11092 2654 11104
rect 5074 11092 5080 11104
rect 5132 11092 5138 11144
rect 5994 11132 6000 11144
rect 5955 11104 6000 11132
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7300 11132 7328 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11200 8355 11203
rect 9769 11203 9827 11209
rect 8343 11172 8524 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 7466 11132 7472 11144
rect 6880 11104 7328 11132
rect 7427 11104 7472 11132
rect 6880 11092 6886 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 8404 11064 8432 11095
rect 7800 11036 8432 11064
rect 8496 11064 8524 11172
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 9815 11172 10609 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 10597 11163 10655 11169
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11698 11160 11704 11212
rect 11756 11200 11762 11212
rect 11756 11172 11801 11200
rect 11756 11160 11762 11172
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 9916 11104 10701 11132
rect 9916 11092 9922 11104
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 11793 11135 11851 11141
rect 11793 11132 11805 11135
rect 10836 11104 11805 11132
rect 10836 11092 10842 11104
rect 11793 11101 11805 11104
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 11054 11064 11060 11076
rect 8496 11036 11060 11064
rect 7800 11024 7806 11036
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 11238 11064 11244 11076
rect 11199 11036 11244 11064
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 12268 11073 12296 11228
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 12952 11172 13645 11200
rect 12952 11160 12958 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 15654 11200 15660 11212
rect 15615 11172 15660 11200
rect 13633 11163 13691 11169
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15746 11160 15752 11212
rect 15804 11200 15810 11212
rect 17313 11203 17371 11209
rect 15804 11172 16896 11200
rect 15804 11160 15810 11172
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13722 11132 13728 11144
rect 12860 11104 12905 11132
rect 13683 11104 13728 11132
rect 12860 11092 12866 11104
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13817 11135 13875 11141
rect 13817 11101 13829 11135
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 12253 11067 12311 11073
rect 12253 11033 12265 11067
rect 12299 11033 12311 11067
rect 12253 11027 12311 11033
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 13832 11064 13860 11095
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 16868 11141 16896 11172
rect 17313 11169 17325 11203
rect 17359 11200 17371 11203
rect 18598 11200 18604 11212
rect 17359 11172 18604 11200
rect 17359 11169 17371 11172
rect 17313 11163 17371 11169
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 14608 11104 15853 11132
rect 14608 11092 14614 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 16761 11135 16819 11141
rect 16761 11101 16773 11135
rect 16807 11101 16819 11135
rect 16761 11095 16819 11101
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 13688 11036 13860 11064
rect 15289 11067 15347 11073
rect 13688 11024 13694 11036
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 16776 11064 16804 11095
rect 17328 11064 17356 11163
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 15335 11036 16804 11064
rect 16868 11036 17356 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 2041 10999 2099 11005
rect 2041 10996 2053 10999
rect 1820 10968 2053 10996
rect 1820 10956 1826 10968
rect 2041 10965 2053 10968
rect 2087 10965 2099 10999
rect 2041 10959 2099 10965
rect 6086 10956 6092 11008
rect 6144 10996 6150 11008
rect 6822 10996 6828 11008
rect 6144 10968 6828 10996
rect 6144 10956 6150 10968
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 15654 10996 15660 11008
rect 10376 10968 15660 10996
rect 10376 10956 10382 10968
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 16022 10956 16028 11008
rect 16080 10996 16086 11008
rect 16868 10996 16896 11036
rect 16080 10968 16896 10996
rect 16080 10956 16086 10968
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7469 10795 7527 10801
rect 7469 10792 7481 10795
rect 7248 10764 7481 10792
rect 7248 10752 7254 10764
rect 7469 10761 7481 10764
rect 7515 10761 7527 10795
rect 10318 10792 10324 10804
rect 7469 10755 7527 10761
rect 7576 10764 10324 10792
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 7576 10724 7604 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11425 10795 11483 10801
rect 11425 10761 11437 10795
rect 11471 10792 11483 10795
rect 12802 10792 12808 10804
rect 11471 10764 12808 10792
rect 11471 10761 11483 10764
rect 11425 10755 11483 10761
rect 4028 10696 7604 10724
rect 4028 10684 4034 10696
rect 11330 10684 11336 10736
rect 11388 10724 11394 10736
rect 11440 10724 11468 10755
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 14274 10792 14280 10804
rect 12912 10764 14280 10792
rect 12912 10724 12940 10764
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14550 10752 14556 10804
rect 14608 10792 14614 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 14608 10764 14749 10792
rect 14608 10752 14614 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 16298 10792 16304 10804
rect 16259 10764 16304 10792
rect 14737 10755 14795 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 16592 10764 19441 10792
rect 11388 10696 11468 10724
rect 12544 10696 12940 10724
rect 11388 10684 11394 10696
rect 1394 10616 1400 10668
rect 1452 10656 1458 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1452 10628 1961 10656
rect 1452 10616 1458 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 3142 10656 3148 10668
rect 3103 10628 3148 10656
rect 1949 10619 2007 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3844 10628 4077 10656
rect 3844 10616 3850 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5534 10656 5540 10668
rect 5307 10628 5540 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7800 10628 8033 10656
rect 7800 10616 7806 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 1762 10588 1768 10600
rect 1723 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 3326 10548 3332 10600
rect 3384 10588 3390 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3384 10560 3985 10588
rect 3384 10548 3390 10560
rect 3973 10557 3985 10560
rect 4019 10557 4031 10591
rect 3973 10551 4031 10557
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10588 5963 10591
rect 7006 10588 7012 10600
rect 5951 10560 7012 10588
rect 5951 10557 5963 10560
rect 5905 10551 5963 10557
rect 7006 10548 7012 10560
rect 7064 10588 7070 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 7064 10560 9137 10588
rect 7064 10548 7070 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9953 10591 10011 10597
rect 9272 10560 9904 10588
rect 9272 10548 9278 10560
rect 2869 10523 2927 10529
rect 2869 10489 2881 10523
rect 2915 10520 2927 10523
rect 3418 10520 3424 10532
rect 2915 10492 3424 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 7837 10523 7895 10529
rect 7837 10489 7849 10523
rect 7883 10520 7895 10523
rect 8481 10523 8539 10529
rect 8481 10520 8493 10523
rect 7883 10492 8493 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8481 10489 8493 10492
rect 8527 10489 8539 10523
rect 9876 10520 9904 10560
rect 9953 10557 9965 10591
rect 9999 10588 10011 10591
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9999 10560 10057 10588
rect 9999 10557 10011 10560
rect 9953 10551 10011 10557
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10312 10591 10370 10597
rect 10312 10557 10324 10591
rect 10358 10588 10370 10591
rect 10778 10588 10784 10600
rect 10358 10560 10784 10588
rect 10358 10557 10370 10560
rect 10312 10551 10370 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 12544 10588 12572 10696
rect 12894 10656 12900 10668
rect 12855 10628 12900 10656
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13262 10616 13268 10668
rect 13320 10656 13326 10668
rect 13357 10659 13415 10665
rect 13357 10656 13369 10659
rect 13320 10628 13369 10656
rect 13320 10616 13326 10628
rect 13357 10625 13369 10628
rect 13403 10625 13415 10659
rect 13357 10619 13415 10625
rect 15010 10616 15016 10668
rect 15068 10656 15074 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15068 10628 15485 10656
rect 15068 10616 15074 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15654 10656 15660 10668
rect 15567 10628 15660 10656
rect 15473 10619 15531 10625
rect 15654 10616 15660 10628
rect 15712 10656 15718 10668
rect 16592 10656 16620 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 16850 10656 16856 10668
rect 15712 10628 16620 10656
rect 16811 10628 16856 10656
rect 15712 10616 15718 10628
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 10888 10560 12572 10588
rect 12805 10591 12863 10597
rect 10888 10520 10916 10560
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 15102 10588 15108 10600
rect 12805 10551 12863 10557
rect 13464 10560 15108 10588
rect 9876 10492 10916 10520
rect 8481 10483 8539 10489
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 12526 10520 12532 10532
rect 11204 10492 12532 10520
rect 11204 10480 11210 10492
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 12820 10520 12848 10551
rect 13464 10520 13492 10560
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18316 10591 18374 10597
rect 18316 10557 18328 10591
rect 18362 10588 18374 10591
rect 18690 10588 18696 10600
rect 18362 10560 18696 10588
rect 18362 10557 18374 10560
rect 18316 10551 18374 10557
rect 13630 10529 13636 10532
rect 13624 10520 13636 10529
rect 12820 10492 13492 10520
rect 13591 10492 13636 10520
rect 13624 10483 13636 10492
rect 13630 10480 13636 10483
rect 13688 10480 13694 10532
rect 16761 10523 16819 10529
rect 16761 10520 16773 10523
rect 15028 10492 16773 10520
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3513 10455 3571 10461
rect 3513 10452 3525 10455
rect 3007 10424 3525 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3513 10421 3525 10424
rect 3559 10421 3571 10455
rect 3513 10415 3571 10421
rect 3881 10455 3939 10461
rect 3881 10421 3893 10455
rect 3927 10452 3939 10455
rect 5534 10452 5540 10464
rect 3927 10424 5540 10452
rect 3927 10421 3939 10424
rect 3881 10415 3939 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 7374 10452 7380 10464
rect 6052 10424 7380 10452
rect 6052 10412 6058 10424
rect 7374 10412 7380 10424
rect 7432 10452 7438 10464
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7432 10424 7941 10452
rect 7432 10412 7438 10424
rect 7929 10421 7941 10424
rect 7975 10421 7987 10455
rect 7929 10415 7987 10421
rect 8570 10412 8576 10464
rect 8628 10452 8634 10464
rect 8941 10455 8999 10461
rect 8941 10452 8953 10455
rect 8628 10424 8953 10452
rect 8628 10412 8634 10424
rect 8941 10421 8953 10424
rect 8987 10452 8999 10455
rect 9953 10455 10011 10461
rect 9953 10452 9965 10455
rect 8987 10424 9965 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9953 10421 9965 10424
rect 9999 10421 10011 10455
rect 9953 10415 10011 10421
rect 12621 10455 12679 10461
rect 12621 10421 12633 10455
rect 12667 10452 12679 10455
rect 12710 10452 12716 10464
rect 12667 10424 12716 10452
rect 12667 10421 12679 10424
rect 12621 10415 12679 10421
rect 12710 10412 12716 10424
rect 12768 10452 12774 10464
rect 13262 10452 13268 10464
rect 12768 10424 13268 10452
rect 12768 10412 12774 10424
rect 13262 10412 13268 10424
rect 13320 10412 13326 10464
rect 15028 10461 15056 10492
rect 16761 10489 16773 10492
rect 16807 10489 16819 10523
rect 18064 10520 18092 10551
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 18598 10520 18604 10532
rect 18064 10492 18604 10520
rect 16761 10483 16819 10489
rect 18598 10480 18604 10492
rect 18656 10480 18662 10532
rect 15013 10455 15071 10461
rect 15013 10421 15025 10455
rect 15059 10421 15071 10455
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 15013 10415 15071 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 16666 10452 16672 10464
rect 16627 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 3200 10220 5457 10248
rect 3200 10208 3206 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6086 10248 6092 10260
rect 5592 10220 6092 10248
rect 5592 10208 5598 10220
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 12437 10251 12495 10257
rect 7852 10220 12204 10248
rect 1848 10183 1906 10189
rect 1848 10149 1860 10183
rect 1894 10180 1906 10183
rect 3160 10180 3188 10208
rect 1894 10152 3188 10180
rect 1894 10149 1906 10152
rect 1848 10143 1906 10149
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4332 10183 4390 10189
rect 4332 10180 4344 10183
rect 3844 10152 4344 10180
rect 3844 10140 3850 10152
rect 4332 10149 4344 10152
rect 4378 10180 4390 10183
rect 7852 10180 7880 10220
rect 4378 10152 7880 10180
rect 11072 10152 12112 10180
rect 4378 10149 4390 10152
rect 4332 10143 4390 10149
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 2774 10112 2780 10124
rect 1627 10084 2780 10112
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 2774 10072 2780 10084
rect 2832 10112 2838 10124
rect 3602 10112 3608 10124
rect 2832 10084 3608 10112
rect 2832 10072 2838 10084
rect 3602 10072 3608 10084
rect 3660 10112 3666 10124
rect 3970 10112 3976 10124
rect 3660 10084 3976 10112
rect 3660 10072 3666 10084
rect 3970 10072 3976 10084
rect 4028 10112 4034 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 4028 10084 4077 10112
rect 4028 10072 4034 10084
rect 4065 10081 4077 10084
rect 4111 10081 4123 10115
rect 4065 10075 4123 10081
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10112 6423 10115
rect 6454 10112 6460 10124
rect 6411 10084 6460 10112
rect 6411 10081 6423 10084
rect 6365 10075 6423 10081
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 6638 10121 6644 10124
rect 6632 10112 6644 10121
rect 6599 10084 6644 10112
rect 6632 10075 6644 10084
rect 6638 10072 6644 10075
rect 6696 10072 6702 10124
rect 8386 10112 8392 10124
rect 8347 10084 8392 10112
rect 8386 10072 8392 10084
rect 8444 10072 8450 10124
rect 8481 10115 8539 10121
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 10226 10112 10232 10124
rect 8527 10084 10232 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11072 10121 11100 10152
rect 11330 10121 11336 10124
rect 11057 10115 11115 10121
rect 11057 10081 11069 10115
rect 11103 10081 11115 10115
rect 11324 10112 11336 10121
rect 11291 10084 11336 10112
rect 11057 10075 11115 10081
rect 11324 10075 11336 10084
rect 11330 10072 11336 10075
rect 11388 10072 11394 10124
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2924 10016 3249 10044
rect 2924 10004 2930 10016
rect 3237 10013 3249 10016
rect 3283 10013 3295 10047
rect 8662 10044 8668 10056
rect 8575 10016 8668 10044
rect 3237 10007 3295 10013
rect 8662 10004 8668 10016
rect 8720 10044 8726 10056
rect 9582 10044 9588 10056
rect 8720 10016 9588 10044
rect 8720 10004 8726 10016
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 12084 10044 12112 10152
rect 12176 10112 12204 10220
rect 12437 10217 12449 10251
rect 12483 10217 12495 10251
rect 12437 10211 12495 10217
rect 12452 10180 12480 10211
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13688 10220 14105 10248
rect 13688 10208 13694 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 12986 10189 12992 10192
rect 12958 10183 12992 10189
rect 12958 10180 12970 10183
rect 12452 10152 12970 10180
rect 12958 10149 12970 10152
rect 13044 10180 13050 10192
rect 16292 10183 16350 10189
rect 13044 10152 13106 10180
rect 12958 10143 12992 10149
rect 12986 10140 12992 10143
rect 13044 10140 13050 10152
rect 16292 10149 16304 10183
rect 16338 10180 16350 10183
rect 16850 10180 16856 10192
rect 16338 10152 16856 10180
rect 16338 10149 16350 10152
rect 16292 10143 16350 10149
rect 16850 10140 16856 10152
rect 16908 10140 16914 10192
rect 12176 10084 17448 10112
rect 12710 10044 12716 10056
rect 12084 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 17420 9985 17448 10084
rect 17405 9979 17463 9985
rect 7300 9948 8156 9976
rect 2590 9868 2596 9920
rect 2648 9908 2654 9920
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2648 9880 2973 9908
rect 2648 9868 2654 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 7300 9908 7328 9948
rect 8018 9908 8024 9920
rect 3936 9880 7328 9908
rect 7979 9880 8024 9908
rect 3936 9868 3942 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8128 9908 8156 9948
rect 17405 9945 17417 9979
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 15378 9908 15384 9920
rect 8128 9880 15384 9908
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 3513 9707 3571 9713
rect 3513 9704 3525 9707
rect 3476 9676 3525 9704
rect 3476 9664 3482 9676
rect 3513 9673 3525 9676
rect 3559 9673 3571 9707
rect 5718 9704 5724 9716
rect 3513 9667 3571 9673
rect 5092 9676 5724 9704
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 1949 9639 2007 9645
rect 1949 9636 1961 9639
rect 1728 9608 1961 9636
rect 1728 9596 1734 9608
rect 1949 9605 1961 9608
rect 1995 9605 2007 9639
rect 1949 9599 2007 9605
rect 3970 9596 3976 9648
rect 4028 9636 4034 9648
rect 5092 9636 5120 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 16022 9704 16028 9716
rect 15396 9676 16028 9704
rect 4028 9608 5120 9636
rect 4028 9596 4034 9608
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 3786 9568 3792 9580
rect 3191 9540 3792 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3786 9528 3792 9540
rect 3844 9568 3850 9580
rect 5092 9577 5120 9608
rect 6457 9639 6515 9645
rect 6457 9605 6469 9639
rect 6503 9605 6515 9639
rect 6457 9599 6515 9605
rect 4065 9571 4123 9577
rect 4065 9568 4077 9571
rect 3844 9540 4077 9568
rect 3844 9528 3850 9540
rect 4065 9537 4077 9540
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 6472 9568 6500 9599
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 9953 9639 10011 9645
rect 9953 9636 9965 9639
rect 9640 9608 9965 9636
rect 9640 9596 9646 9608
rect 9953 9605 9965 9608
rect 9999 9605 10011 9639
rect 10226 9636 10232 9648
rect 10187 9608 10232 9636
rect 9953 9599 10011 9605
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 13722 9636 13728 9648
rect 12483 9608 13728 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 6638 9568 6644 9580
rect 6472 9540 6644 9568
rect 5077 9531 5135 9537
rect 6638 9528 6644 9540
rect 6696 9568 6702 9580
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 6696 9540 7389 9568
rect 6696 9528 6702 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 12986 9568 12992 9580
rect 12947 9540 12992 9568
rect 10781 9531 10839 9537
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 4706 9500 4712 9512
rect 1811 9472 4712 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 7190 9500 7196 9512
rect 5276 9472 7196 9500
rect 2869 9435 2927 9441
rect 2869 9401 2881 9435
rect 2915 9432 2927 9435
rect 3050 9432 3056 9444
rect 2915 9404 3056 9432
rect 2915 9401 2927 9404
rect 2869 9395 2927 9401
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 3973 9435 4031 9441
rect 3973 9432 3985 9435
rect 3844 9404 3985 9432
rect 3844 9392 3850 9404
rect 3973 9401 3985 9404
rect 4019 9432 4031 9435
rect 5276 9432 5304 9472
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9500 7343 9503
rect 8018 9500 8024 9512
rect 7331 9472 8024 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8840 9503 8898 9509
rect 8840 9469 8852 9503
rect 8886 9500 8898 9503
rect 9122 9500 9128 9512
rect 8886 9472 9128 9500
rect 8886 9469 8898 9472
rect 8840 9463 8898 9469
rect 9122 9460 9128 9472
rect 9180 9500 9186 9512
rect 10796 9500 10824 9531
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 15396 9577 15424 9676
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 16761 9707 16819 9713
rect 16761 9673 16773 9707
rect 16807 9704 16819 9707
rect 16850 9704 16856 9716
rect 16807 9676 16856 9704
rect 16807 9673 16819 9676
rect 16761 9667 16819 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 15381 9571 15439 9577
rect 15381 9537 15393 9571
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16724 9540 17049 9568
rect 16724 9528 16730 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 9180 9472 10824 9500
rect 9180 9460 9186 9472
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 12805 9503 12863 9509
rect 12805 9500 12817 9503
rect 12584 9472 12817 9500
rect 12584 9460 12590 9472
rect 12805 9469 12817 9472
rect 12851 9469 12863 9503
rect 12805 9463 12863 9469
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13998 9500 14004 9512
rect 12943 9472 14004 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13998 9460 14004 9472
rect 14056 9500 14062 9512
rect 15010 9500 15016 9512
rect 14056 9472 15016 9500
rect 14056 9460 14062 9472
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15654 9509 15660 9512
rect 15648 9500 15660 9509
rect 15615 9472 15660 9500
rect 15648 9463 15660 9472
rect 15654 9460 15660 9463
rect 15712 9460 15718 9512
rect 4019 9404 5304 9432
rect 5344 9435 5402 9441
rect 4019 9401 4031 9404
rect 3973 9395 4031 9401
rect 5344 9401 5356 9435
rect 5390 9432 5402 9435
rect 6730 9432 6736 9444
rect 5390 9404 6736 9432
rect 5390 9401 5402 9404
rect 5344 9395 5402 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 7208 9432 7236 9460
rect 8478 9432 8484 9444
rect 7208 9404 8484 9432
rect 8478 9392 8484 9404
rect 8536 9392 8542 9444
rect 10689 9435 10747 9441
rect 10689 9401 10701 9435
rect 10735 9432 10747 9435
rect 12342 9432 12348 9444
rect 10735 9404 12348 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 2498 9364 2504 9376
rect 2459 9336 2504 9364
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2958 9364 2964 9376
rect 2919 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3881 9367 3939 9373
rect 3881 9364 3893 9367
rect 3660 9336 3893 9364
rect 3660 9324 3666 9336
rect 3881 9333 3893 9336
rect 3927 9333 3939 9367
rect 3881 9327 3939 9333
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 4856 9336 6837 9364
rect 4856 9324 4862 9336
rect 6825 9333 6837 9336
rect 6871 9333 6883 9367
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 6825 9327 6883 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 9306 9364 9312 9376
rect 7524 9336 9312 9364
rect 7524 9324 7530 9336
rect 9306 9324 9312 9336
rect 9364 9364 9370 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 9364 9336 10609 9364
rect 9364 9324 9370 9336
rect 10597 9333 10609 9336
rect 10643 9333 10655 9367
rect 10597 9327 10655 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2556 9132 2973 9160
rect 2556 9120 2562 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 6089 9163 6147 9169
rect 6089 9129 6101 9163
rect 6135 9160 6147 9163
rect 7190 9160 7196 9172
rect 6135 9132 7196 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8386 9160 8392 9172
rect 8347 9132 8392 9160
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 2866 9092 2872 9104
rect 2827 9064 2872 9092
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 18966 9092 18972 9104
rect 4120 9064 18972 9092
rect 4120 9052 4126 9064
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 6503 8996 7113 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 7101 8993 7113 8996
rect 7147 8993 7159 9027
rect 8754 9024 8760 9036
rect 8715 8996 8760 9024
rect 7101 8987 7159 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 9398 9024 9404 9036
rect 8864 8996 9404 9024
rect 8864 8968 8892 8996
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 5408 8928 6561 8956
rect 5408 8916 5414 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6730 8956 6736 8968
rect 6643 8928 6736 8956
rect 6549 8919 6607 8925
rect 6730 8916 6736 8928
rect 6788 8956 6794 8968
rect 8662 8956 8668 8968
rect 6788 8928 8668 8956
rect 6788 8916 6794 8928
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 8846 8956 8852 8968
rect 8807 8928 8852 8956
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8956 9091 8959
rect 9122 8956 9128 8968
rect 9079 8928 9128 8956
rect 9079 8925 9091 8928
rect 9033 8919 9091 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2501 8891 2559 8897
rect 2501 8888 2513 8891
rect 2464 8860 2513 8888
rect 2464 8848 2470 8860
rect 2501 8857 2513 8860
rect 2547 8857 2559 8891
rect 2501 8851 2559 8857
rect 4154 8848 4160 8900
rect 4212 8888 4218 8900
rect 8754 8888 8760 8900
rect 4212 8860 8760 8888
rect 4212 8848 4218 8860
rect 8754 8848 8760 8860
rect 8812 8848 8818 8900
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 15286 8820 15292 8832
rect 4028 8792 15292 8820
rect 4028 8780 4034 8792
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2774 8616 2780 8628
rect 1780 8588 2780 8616
rect 1780 8489 1808 8588
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 7374 8616 7380 8628
rect 3108 8588 7380 8616
rect 3108 8576 3114 8588
rect 7374 8576 7380 8588
rect 7432 8576 7438 8628
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9217 8619 9275 8625
rect 9217 8616 9229 8619
rect 9180 8588 9229 8616
rect 9180 8576 9186 8588
rect 9217 8585 9229 8588
rect 9263 8585 9275 8619
rect 9217 8579 9275 8585
rect 3789 8551 3847 8557
rect 3789 8517 3801 8551
rect 3835 8548 3847 8551
rect 5442 8548 5448 8560
rect 3835 8520 5448 8548
rect 3835 8517 3847 8520
rect 3789 8511 3847 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1780 8412 1808 8443
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 4338 8480 4344 8492
rect 3200 8452 4344 8480
rect 3200 8440 3206 8452
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 4764 8452 5641 8480
rect 4764 8440 4770 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7742 8480 7748 8492
rect 7515 8452 7748 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7742 8440 7748 8452
rect 7800 8480 7806 8492
rect 7800 8452 7972 8480
rect 7800 8440 7806 8452
rect 1854 8412 1860 8424
rect 1780 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2032 8415 2090 8421
rect 2032 8381 2044 8415
rect 2078 8412 2090 8415
rect 2590 8412 2596 8424
rect 2078 8384 2596 8412
rect 2078 8381 2090 8384
rect 2032 8375 2090 8381
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 4154 8344 4160 8356
rect 4115 8316 4160 8344
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 5460 8344 5488 8375
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7837 8415 7895 8421
rect 7837 8412 7849 8415
rect 6972 8384 7849 8412
rect 6972 8372 6978 8384
rect 7837 8381 7849 8384
rect 7883 8381 7895 8415
rect 7944 8412 7972 8452
rect 8093 8415 8151 8421
rect 8093 8412 8105 8415
rect 7944 8384 8105 8412
rect 7837 8375 7895 8381
rect 8093 8381 8105 8384
rect 8139 8381 8151 8415
rect 8093 8375 8151 8381
rect 7190 8344 7196 8356
rect 5460 8316 6868 8344
rect 7151 8316 7196 8344
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 4246 8276 4252 8288
rect 4207 8248 4252 8276
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 6840 8285 6868 8316
rect 7190 8304 7196 8316
rect 7248 8304 7254 8356
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 7852 8344 7880 8375
rect 8570 8344 8576 8356
rect 7340 8316 7385 8344
rect 7852 8316 8576 8344
rect 7340 8304 7346 8316
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 6825 8279 6883 8285
rect 6825 8245 6837 8279
rect 6871 8245 6883 8279
rect 6825 8239 6883 8245
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 13538 8276 13544 8288
rect 7064 8248 13544 8276
rect 7064 8236 7070 8248
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4798 8072 4804 8084
rect 4571 8044 4804 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 2124 8007 2182 8013
rect 2124 7973 2136 8007
rect 2170 8004 2182 8007
rect 3142 8004 3148 8016
rect 2170 7976 3148 8004
rect 2170 7973 2182 7976
rect 2124 7967 2182 7973
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 4080 8004 4108 8035
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5442 8072 5448 8084
rect 5403 8044 5448 8072
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 7006 8072 7012 8084
rect 6503 8044 7012 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7800 8044 7941 8072
rect 7800 8032 7806 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8849 8075 8907 8081
rect 8849 8072 8861 8075
rect 8343 8044 8861 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8849 8041 8861 8044
rect 8895 8072 8907 8075
rect 11790 8072 11796 8084
rect 8895 8044 11796 8072
rect 8895 8041 8907 8044
rect 8849 8035 8907 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 19061 8075 19119 8081
rect 12268 8044 18920 8072
rect 5537 8007 5595 8013
rect 5537 8004 5549 8007
rect 4080 7976 5549 8004
rect 5537 7973 5549 7976
rect 5583 7973 5595 8007
rect 5537 7967 5595 7973
rect 6816 8007 6874 8013
rect 6816 7973 6828 8007
rect 6862 8004 6874 8007
rect 6914 8004 6920 8016
rect 6862 7976 6920 8004
rect 6862 7973 6874 7976
rect 6816 7967 6874 7973
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 7466 7964 7472 8016
rect 7524 7964 7530 8016
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 12268 8004 12296 8044
rect 7708 7976 12296 8004
rect 7708 7964 7714 7976
rect 1854 7936 1860 7948
rect 1815 7908 1860 7936
rect 1854 7896 1860 7908
rect 1912 7896 1918 7948
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4028 7908 4445 7936
rect 4028 7896 4034 7908
rect 4433 7905 4445 7908
rect 4479 7936 4491 7939
rect 7484 7936 7512 7964
rect 18892 7945 18920 8044
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19334 8072 19340 8084
rect 19107 8044 19340 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 8757 7939 8815 7945
rect 8757 7936 8769 7939
rect 4479 7908 7512 7936
rect 7576 7908 8769 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 4617 7831 4675 7837
rect 4724 7840 5641 7868
rect 4338 7760 4344 7812
rect 4396 7800 4402 7812
rect 4632 7800 4660 7831
rect 4396 7772 4660 7800
rect 4396 7760 4402 7772
rect 3234 7732 3240 7744
rect 3147 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7732 3298 7744
rect 4724 7732 4752 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 5629 7831 5687 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 4798 7760 4804 7812
rect 4856 7800 4862 7812
rect 4985 7803 5043 7809
rect 4985 7800 4997 7803
rect 4856 7772 4997 7800
rect 4856 7760 4862 7772
rect 4985 7769 4997 7772
rect 5031 7800 5043 7803
rect 6457 7803 6515 7809
rect 6457 7800 6469 7803
rect 5031 7772 6469 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 6457 7769 6469 7772
rect 6503 7769 6515 7803
rect 6457 7763 6515 7769
rect 5074 7732 5080 7744
rect 3292 7704 4752 7732
rect 5035 7704 5080 7732
rect 3292 7692 3298 7704
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 6086 7692 6092 7744
rect 6144 7732 6150 7744
rect 7576 7732 7604 7908
rect 8757 7905 8769 7908
rect 8803 7905 8815 7939
rect 8757 7899 8815 7905
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 8938 7868 8944 7880
rect 8899 7840 8944 7868
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 8386 7732 8392 7744
rect 6144 7704 7604 7732
rect 8347 7704 8392 7732
rect 6144 7692 6150 7704
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 4249 7531 4307 7537
rect 4249 7528 4261 7531
rect 2516 7500 4261 7528
rect 2516 7401 2544 7500
rect 4249 7497 4261 7500
rect 4295 7497 4307 7531
rect 19518 7528 19524 7540
rect 19479 7500 19524 7528
rect 4249 7491 4307 7497
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7361 2559 7395
rect 4264 7392 4292 7491
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 6822 7460 6828 7472
rect 6420 7432 6828 7460
rect 6420 7420 6426 7432
rect 6822 7420 6828 7432
rect 6880 7460 6886 7472
rect 8294 7460 8300 7472
rect 6880 7432 8300 7460
rect 6880 7420 6886 7432
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 4264 7364 4660 7392
rect 2501 7355 2559 7361
rect 1854 7284 1860 7336
rect 1912 7324 1918 7336
rect 2869 7327 2927 7333
rect 2869 7324 2881 7327
rect 1912 7296 2881 7324
rect 1912 7284 1918 7296
rect 2869 7293 2881 7296
rect 2915 7324 2927 7327
rect 4522 7324 4528 7336
rect 2915 7296 4528 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 4522 7284 4528 7296
rect 4580 7284 4586 7336
rect 4632 7324 4660 7364
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 7653 7395 7711 7401
rect 7653 7392 7665 7395
rect 6052 7364 7665 7392
rect 6052 7352 6058 7364
rect 7653 7361 7665 7364
rect 7699 7392 7711 7395
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 7699 7364 8677 7392
rect 7699 7361 7711 7364
rect 7653 7355 7711 7361
rect 8665 7361 8677 7364
rect 8711 7392 8723 7395
rect 8938 7392 8944 7404
rect 8711 7364 8944 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 4781 7327 4839 7333
rect 4781 7324 4793 7327
rect 4632 7296 4793 7324
rect 4781 7293 4793 7296
rect 4827 7293 4839 7327
rect 7374 7324 7380 7336
rect 7335 7296 7380 7324
rect 4781 7287 4839 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 19343 7327 19401 7333
rect 19343 7293 19355 7327
rect 19389 7293 19401 7327
rect 19343 7287 19401 7293
rect 2225 7259 2283 7265
rect 2225 7225 2237 7259
rect 2271 7256 2283 7259
rect 2958 7256 2964 7268
rect 2271 7228 2964 7256
rect 2271 7225 2283 7228
rect 2225 7219 2283 7225
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 3136 7259 3194 7265
rect 3136 7225 3148 7259
rect 3182 7256 3194 7259
rect 3234 7256 3240 7268
rect 3182 7228 3240 7256
rect 3182 7225 3194 7228
rect 3136 7219 3194 7225
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 5718 7216 5724 7268
rect 5776 7256 5782 7268
rect 7469 7259 7527 7265
rect 7469 7256 7481 7259
rect 5776 7228 7481 7256
rect 5776 7216 5782 7228
rect 7469 7225 7481 7228
rect 7515 7225 7527 7259
rect 7469 7219 7527 7225
rect 7742 7216 7748 7268
rect 7800 7256 7806 7268
rect 12342 7256 12348 7268
rect 7800 7228 12348 7256
rect 7800 7216 7806 7228
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 1854 7188 1860 7200
rect 1815 7160 1860 7188
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 5074 7188 5080 7200
rect 2363 7160 5080 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 5994 7188 6000 7200
rect 5951 7160 6000 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6270 7188 6276 7200
rect 6231 7160 6276 7188
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 7006 7188 7012 7200
rect 6967 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 8021 7191 8079 7197
rect 8021 7188 8033 7191
rect 7616 7160 8033 7188
rect 7616 7148 7622 7160
rect 8021 7157 8033 7160
rect 8067 7157 8079 7191
rect 8021 7151 8079 7157
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8352 7160 8401 7188
rect 8352 7148 8358 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 8389 7151 8447 7157
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 19352 7188 19380 7287
rect 12492 7160 19380 7188
rect 12492 7148 12498 7160
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 2958 6984 2964 6996
rect 2919 6956 2964 6984
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 6822 6984 6828 6996
rect 3660 6956 6828 6984
rect 3660 6944 3666 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7745 6987 7803 6993
rect 7745 6984 7757 6987
rect 7064 6956 7757 6984
rect 7064 6944 7070 6956
rect 7745 6953 7757 6956
rect 7791 6953 7803 6987
rect 7745 6947 7803 6953
rect 2866 6876 2872 6928
rect 2924 6916 2930 6928
rect 5718 6916 5724 6928
rect 2924 6888 5724 6916
rect 2924 6876 2930 6888
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 5896 6919 5954 6925
rect 5896 6885 5908 6919
rect 5942 6916 5954 6919
rect 5994 6916 6000 6928
rect 5942 6888 6000 6916
rect 5942 6885 5954 6888
rect 5896 6879 5954 6885
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 6328 6888 7665 6916
rect 6328 6876 6334 6888
rect 7653 6885 7665 6888
rect 7699 6885 7711 6919
rect 7653 6879 7711 6885
rect 1854 6848 1860 6860
rect 1815 6820 1860 6848
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 3375 6820 4077 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 4065 6817 4077 6820
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4522 6808 4528 6860
rect 4580 6848 4586 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 4580 6820 5641 6848
rect 4580 6808 4586 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 19702 6848 19708 6860
rect 19663 6820 19708 6848
rect 5629 6811 5687 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 20257 6851 20315 6857
rect 20257 6817 20269 6851
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 1762 6740 1768 6792
rect 1820 6780 1826 6792
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1820 6752 2053 6780
rect 1820 6740 1826 6752
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3421 6783 3479 6789
rect 3421 6780 3433 6783
rect 3200 6752 3433 6780
rect 3200 6740 3206 6752
rect 3421 6749 3433 6752
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 7650 6780 7656 6792
rect 3605 6743 3663 6749
rect 7024 6752 7656 6780
rect 3234 6672 3240 6724
rect 3292 6712 3298 6724
rect 3620 6712 3648 6743
rect 5350 6712 5356 6724
rect 3292 6684 3648 6712
rect 3804 6684 5356 6712
rect 3292 6672 3298 6684
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3804 6644 3832 6684
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 7024 6721 7052 6752
rect 7650 6740 7656 6752
rect 7708 6780 7714 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7708 6752 7849 6780
rect 7708 6740 7714 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 7009 6715 7067 6721
rect 7009 6712 7021 6715
rect 6972 6684 7021 6712
rect 6972 6672 6978 6684
rect 7009 6681 7021 6684
rect 7055 6681 7067 6715
rect 7009 6675 7067 6681
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7285 6715 7343 6721
rect 7285 6712 7297 6715
rect 7248 6684 7297 6712
rect 7248 6672 7254 6684
rect 7285 6681 7297 6684
rect 7331 6681 7343 6715
rect 19886 6712 19892 6724
rect 19847 6684 19892 6712
rect 7285 6675 7343 6681
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 3200 6616 3832 6644
rect 3200 6604 3206 6616
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 20272 6644 20300 6811
rect 20441 6715 20499 6721
rect 20441 6681 20453 6715
rect 20487 6712 20499 6715
rect 20990 6712 20996 6724
rect 20487 6684 20996 6712
rect 20487 6681 20499 6684
rect 20441 6675 20499 6681
rect 20990 6672 20996 6684
rect 21048 6672 21054 6724
rect 3936 6616 20300 6644
rect 3936 6604 3942 6616
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7282 6440 7288 6452
rect 7147 6412 7288 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 20717 6443 20775 6449
rect 20717 6409 20729 6443
rect 20763 6440 20775 6443
rect 20898 6440 20904 6452
rect 20763 6412 20904 6440
rect 20763 6409 20775 6412
rect 20717 6403 20775 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 19702 6372 19708 6384
rect 4120 6344 19708 6372
rect 4120 6332 4126 6344
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 7650 6304 7656 6316
rect 7611 6276 7656 6304
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6236 7527 6239
rect 7558 6236 7564 6248
rect 7515 6208 7564 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 20539 6239 20597 6245
rect 12268 6208 14504 6236
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 12268 6168 12296 6208
rect 4764 6140 12296 6168
rect 4764 6128 4770 6140
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 8386 6100 8392 6112
rect 7607 6072 8392 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 14476 6100 14504 6208
rect 20539 6205 20551 6239
rect 20585 6205 20597 6239
rect 20539 6199 20597 6205
rect 20548 6100 20576 6199
rect 14476 6072 20576 6100
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 12618 5352 12624 5364
rect 3752 5324 12624 5352
rect 3752 5312 3758 5324
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20806 5352 20812 5364
rect 20763 5324 20812 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 20533 5151 20591 5157
rect 20533 5148 20545 5151
rect 4120 5120 20545 5148
rect 4120 5108 4126 5120
rect 20533 5117 20545 5120
rect 20579 5117 20591 5151
rect 20533 5111 20591 5117
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 10134 4128 10140 4140
rect 5776 4100 10140 4128
rect 5776 4088 5782 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 6086 1340 6092 1352
rect 3384 1312 6092 1340
rect 3384 1300 3390 1312
rect 6086 1300 6092 1312
rect 6144 1300 6150 1352
rect 16574 552 16580 604
rect 16632 592 16638 604
rect 17126 592 17132 604
rect 16632 564 17132 592
rect 16632 552 16638 564
rect 17126 552 17132 564
rect 17184 552 17190 604
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 5724 20000 5776 20052
rect 9496 20000 9548 20052
rect 13636 20000 13688 20052
rect 15200 20000 15252 20052
rect 16580 20000 16632 20052
rect 17408 20000 17460 20052
rect 18328 20000 18380 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 6368 19864 6420 19916
rect 11612 19864 11664 19916
rect 12808 19864 12860 19916
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 6460 19796 6512 19848
rect 2872 19728 2924 19780
rect 2964 19660 3016 19712
rect 8852 19660 8904 19712
rect 10324 19796 10376 19848
rect 13360 19796 13412 19848
rect 15200 19864 15252 19916
rect 16580 19907 16632 19916
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 16580 19873 16589 19907
rect 16589 19873 16623 19907
rect 16623 19873 16632 19907
rect 16580 19864 16632 19873
rect 16672 19864 16724 19916
rect 18788 19864 18840 19916
rect 15568 19728 15620 19780
rect 9864 19660 9916 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 2504 19456 2556 19508
rect 6460 19499 6512 19508
rect 6460 19465 6469 19499
rect 6469 19465 6503 19499
rect 6503 19465 6512 19499
rect 6460 19456 6512 19465
rect 7196 19456 7248 19508
rect 13820 19456 13872 19508
rect 1768 19320 1820 19372
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 2964 19252 3016 19304
rect 204 19184 256 19236
rect 2412 19184 2464 19236
rect 3148 19252 3200 19304
rect 1676 19116 1728 19168
rect 5080 19295 5132 19304
rect 5080 19261 5089 19295
rect 5089 19261 5123 19295
rect 5123 19261 5132 19295
rect 5080 19252 5132 19261
rect 6736 19252 6788 19304
rect 7380 19252 7432 19304
rect 5724 19184 5776 19236
rect 6460 19184 6512 19236
rect 7196 19184 7248 19236
rect 10508 19252 10560 19304
rect 11060 19252 11112 19304
rect 12624 19252 12676 19304
rect 13820 19320 13872 19372
rect 9496 19227 9548 19236
rect 9496 19193 9530 19227
rect 9530 19193 9548 19227
rect 9496 19184 9548 19193
rect 9588 19184 9640 19236
rect 13912 19252 13964 19304
rect 15016 19320 15068 19372
rect 15752 19252 15804 19304
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 16856 19295 16908 19304
rect 16856 19261 16865 19295
rect 16865 19261 16899 19295
rect 16899 19261 16908 19295
rect 16856 19252 16908 19261
rect 3700 19116 3752 19168
rect 3792 19116 3844 19168
rect 4712 19116 4764 19168
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 9680 19116 9732 19168
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 11796 19116 11848 19168
rect 12348 19116 12400 19168
rect 13176 19116 13228 19168
rect 17960 19252 18012 19304
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 18144 19184 18196 19236
rect 18880 19184 18932 19236
rect 14004 19159 14056 19168
rect 14004 19125 14013 19159
rect 14013 19125 14047 19159
rect 14047 19125 14056 19159
rect 14004 19116 14056 19125
rect 14280 19116 14332 19168
rect 16028 19116 16080 19168
rect 17132 19116 17184 19168
rect 17868 19116 17920 19168
rect 19248 19116 19300 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 5264 18912 5316 18964
rect 6736 18912 6788 18964
rect 8760 18955 8812 18964
rect 2320 18887 2372 18896
rect 2320 18853 2329 18887
rect 2329 18853 2363 18887
rect 2363 18853 2372 18887
rect 2320 18844 2372 18853
rect 2412 18776 2464 18828
rect 8760 18921 8769 18955
rect 8769 18921 8803 18955
rect 8803 18921 8812 18955
rect 8760 18912 8812 18921
rect 8852 18955 8904 18964
rect 8852 18921 8861 18955
rect 8861 18921 8895 18955
rect 8895 18921 8904 18955
rect 8852 18912 8904 18921
rect 3148 18819 3200 18828
rect 3148 18785 3157 18819
rect 3157 18785 3191 18819
rect 3191 18785 3200 18819
rect 3148 18776 3200 18785
rect 4252 18776 4304 18828
rect 1492 18708 1544 18760
rect 2688 18708 2740 18760
rect 3332 18751 3384 18760
rect 3332 18717 3341 18751
rect 3341 18717 3375 18751
rect 3375 18717 3384 18751
rect 3332 18708 3384 18717
rect 3792 18708 3844 18760
rect 5172 18640 5224 18692
rect 9864 18844 9916 18896
rect 11704 18912 11756 18964
rect 14556 18912 14608 18964
rect 11980 18844 12032 18896
rect 12808 18887 12860 18896
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 5724 18751 5776 18760
rect 5724 18717 5733 18751
rect 5733 18717 5767 18751
rect 5767 18717 5776 18751
rect 5724 18708 5776 18717
rect 6460 18708 6512 18760
rect 9404 18776 9456 18828
rect 9588 18776 9640 18828
rect 9128 18708 9180 18760
rect 12164 18776 12216 18828
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 12808 18853 12817 18887
rect 12817 18853 12851 18887
rect 12851 18853 12860 18887
rect 12808 18844 12860 18853
rect 15200 18844 15252 18896
rect 16856 18844 16908 18896
rect 18604 18912 18656 18964
rect 18144 18844 18196 18896
rect 18788 18887 18840 18896
rect 18788 18853 18797 18887
rect 18797 18853 18831 18887
rect 18831 18853 18840 18887
rect 18788 18844 18840 18853
rect 13820 18819 13872 18828
rect 13820 18785 13854 18819
rect 13854 18785 13872 18819
rect 13820 18776 13872 18785
rect 15568 18776 15620 18828
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 16672 18776 16724 18828
rect 11152 18708 11204 18760
rect 12072 18708 12124 18760
rect 12440 18708 12492 18760
rect 16396 18708 16448 18760
rect 11888 18640 11940 18692
rect 9496 18572 9548 18624
rect 11152 18572 11204 18624
rect 15660 18640 15712 18692
rect 18788 18708 18840 18760
rect 18512 18640 18564 18692
rect 15016 18572 15068 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 3608 18368 3660 18420
rect 2412 18300 2464 18352
rect 3700 18300 3752 18352
rect 4712 18300 4764 18352
rect 6460 18343 6512 18352
rect 6460 18309 6469 18343
rect 6469 18309 6503 18343
rect 6503 18309 6512 18343
rect 6460 18300 6512 18309
rect 1584 18232 1636 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 9036 18232 9088 18284
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 2320 18164 2372 18216
rect 1124 18096 1176 18148
rect 3792 18164 3844 18216
rect 4712 18164 4764 18216
rect 5080 18207 5132 18216
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 9772 18164 9824 18216
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 3516 18096 3568 18148
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 5908 18096 5960 18148
rect 11152 18164 11204 18216
rect 10600 18139 10652 18148
rect 10600 18105 10634 18139
rect 10634 18105 10652 18139
rect 10600 18096 10652 18105
rect 14188 18368 14240 18420
rect 14004 18300 14056 18352
rect 15200 18275 15252 18284
rect 12256 18164 12308 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 14096 18207 14148 18216
rect 14096 18173 14105 18207
rect 14105 18173 14139 18207
rect 14139 18173 14148 18207
rect 14096 18164 14148 18173
rect 12992 18096 13044 18148
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 17776 18300 17828 18352
rect 22468 18300 22520 18352
rect 16580 18275 16632 18284
rect 16580 18241 16589 18275
rect 16589 18241 16623 18275
rect 16623 18241 16632 18275
rect 16580 18232 16632 18241
rect 17960 18232 18012 18284
rect 14372 18164 14424 18216
rect 15844 18164 15896 18216
rect 19064 18164 19116 18216
rect 15108 18139 15160 18148
rect 6276 18028 6328 18080
rect 7564 18028 7616 18080
rect 8760 18071 8812 18080
rect 8760 18037 8769 18071
rect 8769 18037 8803 18071
rect 8803 18037 8812 18071
rect 8760 18028 8812 18037
rect 9036 18071 9088 18080
rect 9036 18037 9045 18071
rect 9045 18037 9079 18071
rect 9079 18037 9088 18071
rect 9036 18028 9088 18037
rect 9404 18071 9456 18080
rect 9404 18037 9413 18071
rect 9413 18037 9447 18071
rect 9447 18037 9456 18071
rect 9404 18028 9456 18037
rect 10416 18028 10468 18080
rect 11152 18028 11204 18080
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 13820 18071 13872 18080
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 15108 18105 15117 18139
rect 15117 18105 15151 18139
rect 15151 18105 15160 18139
rect 15108 18096 15160 18105
rect 19524 18096 19576 18148
rect 20168 18096 20220 18148
rect 20812 18096 20864 18148
rect 22008 18096 22060 18148
rect 14556 18028 14608 18080
rect 19892 18028 19944 18080
rect 20628 18028 20680 18080
rect 20904 18028 20956 18080
rect 21548 18028 21600 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 2780 17824 2832 17876
rect 3056 17867 3108 17876
rect 3056 17833 3065 17867
rect 3065 17833 3099 17867
rect 3099 17833 3108 17867
rect 3056 17824 3108 17833
rect 3148 17824 3200 17876
rect 5540 17824 5592 17876
rect 6184 17824 6236 17876
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 2412 17688 2464 17740
rect 3332 17688 3384 17740
rect 4068 17688 4120 17740
rect 9036 17824 9088 17876
rect 9956 17824 10008 17876
rect 13912 17824 13964 17876
rect 14280 17824 14332 17876
rect 14556 17867 14608 17876
rect 14556 17833 14565 17867
rect 14565 17833 14599 17867
rect 14599 17833 14608 17867
rect 14556 17824 14608 17833
rect 15660 17867 15712 17876
rect 15660 17833 15669 17867
rect 15669 17833 15703 17867
rect 15703 17833 15712 17867
rect 15660 17824 15712 17833
rect 16028 17824 16080 17876
rect 9404 17756 9456 17808
rect 9772 17756 9824 17808
rect 12256 17756 12308 17808
rect 15200 17756 15252 17808
rect 7932 17731 7984 17740
rect 7932 17697 7941 17731
rect 7941 17697 7975 17731
rect 7975 17697 7984 17731
rect 7932 17688 7984 17697
rect 9956 17688 10008 17740
rect 12808 17731 12860 17740
rect 5908 17620 5960 17672
rect 8300 17620 8352 17672
rect 8760 17620 8812 17672
rect 5816 17484 5868 17536
rect 9404 17620 9456 17672
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 17132 17756 17184 17808
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 12992 17663 13044 17672
rect 12992 17629 13001 17663
rect 13001 17629 13035 17663
rect 13035 17629 13044 17663
rect 12992 17620 13044 17629
rect 13820 17620 13872 17672
rect 15660 17620 15712 17672
rect 17776 17688 17828 17740
rect 16488 17620 16540 17672
rect 10416 17484 10468 17536
rect 18604 17484 18656 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 5816 17280 5868 17332
rect 5908 17280 5960 17332
rect 7380 17280 7432 17332
rect 9956 17323 10008 17332
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 12716 17280 12768 17332
rect 13544 17280 13596 17332
rect 14372 17280 14424 17332
rect 2412 17144 2464 17196
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 11704 17144 11756 17196
rect 12440 17144 12492 17196
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 3332 17076 3384 17128
rect 4712 17076 4764 17128
rect 7012 17076 7064 17128
rect 9680 17076 9732 17128
rect 10968 17076 11020 17128
rect 13268 17076 13320 17128
rect 5264 17008 5316 17060
rect 6920 17008 6972 17060
rect 13084 17008 13136 17060
rect 15016 17076 15068 17128
rect 16304 17280 16356 17332
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 15476 17008 15528 17060
rect 18972 17076 19024 17128
rect 19156 17076 19208 17128
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 4068 16940 4120 16992
rect 12440 16940 12492 16992
rect 12900 16940 12952 16992
rect 12992 16940 13044 16992
rect 14556 16940 14608 16992
rect 16948 16983 17000 16992
rect 16948 16949 16957 16983
rect 16957 16949 16991 16983
rect 16991 16949 17000 16983
rect 16948 16940 17000 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 2044 16736 2096 16788
rect 6644 16736 6696 16788
rect 10600 16736 10652 16788
rect 12532 16736 12584 16788
rect 17132 16736 17184 16788
rect 3240 16668 3292 16720
rect 8300 16668 8352 16720
rect 16488 16668 16540 16720
rect 2044 16600 2096 16652
rect 5540 16600 5592 16652
rect 7104 16600 7156 16652
rect 7380 16600 7432 16652
rect 9772 16643 9824 16652
rect 9772 16609 9781 16643
rect 9781 16609 9815 16643
rect 9815 16609 9824 16643
rect 9772 16600 9824 16609
rect 10784 16600 10836 16652
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 16212 16643 16264 16652
rect 16212 16609 16246 16643
rect 16246 16609 16264 16643
rect 16212 16600 16264 16609
rect 18604 16668 18656 16720
rect 17868 16600 17920 16652
rect 1768 16532 1820 16584
rect 5264 16532 5316 16584
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 12440 16532 12492 16584
rect 13084 16532 13136 16584
rect 8668 16439 8720 16448
rect 8668 16405 8677 16439
rect 8677 16405 8711 16439
rect 8711 16405 8720 16439
rect 8668 16396 8720 16405
rect 19156 16439 19208 16448
rect 19156 16405 19165 16439
rect 19165 16405 19199 16439
rect 19199 16405 19208 16439
rect 19156 16396 19208 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 5264 16192 5316 16244
rect 7104 16192 7156 16244
rect 10784 16235 10836 16244
rect 2044 16056 2096 16108
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 13084 16192 13136 16244
rect 15476 16192 15528 16244
rect 16948 16192 17000 16244
rect 2504 15988 2556 16040
rect 2688 16031 2740 16040
rect 2688 15997 2697 16031
rect 2697 15997 2731 16031
rect 2731 15997 2740 16031
rect 2688 15988 2740 15997
rect 2872 15988 2924 16040
rect 4528 15988 4580 16040
rect 4712 15988 4764 16040
rect 6092 15920 6144 15972
rect 6920 15988 6972 16040
rect 7380 15988 7432 16040
rect 8668 15920 8720 15972
rect 11152 16056 11204 16108
rect 9956 15988 10008 16040
rect 13268 15988 13320 16040
rect 14372 16056 14424 16108
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 12624 15920 12676 15972
rect 12900 15920 12952 15972
rect 3056 15852 3108 15904
rect 4804 15852 4856 15904
rect 6920 15852 6972 15904
rect 7196 15852 7248 15904
rect 10048 15852 10100 15904
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 12256 15852 12308 15904
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 14464 15852 14516 15861
rect 15384 15852 15436 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 5540 15648 5592 15700
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 8208 15648 8260 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 11060 15648 11112 15700
rect 4068 15580 4120 15632
rect 4528 15580 4580 15632
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 14096 15648 14148 15700
rect 16212 15648 16264 15700
rect 12716 15580 12768 15632
rect 14372 15580 14424 15632
rect 15936 15580 15988 15632
rect 19156 15580 19208 15632
rect 1768 15555 1820 15564
rect 1768 15521 1777 15555
rect 1777 15521 1811 15555
rect 1811 15521 1820 15555
rect 1768 15512 1820 15521
rect 7012 15512 7064 15564
rect 12440 15512 12492 15564
rect 15476 15512 15528 15564
rect 16488 15512 16540 15564
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 4068 15487 4120 15496
rect 4068 15453 4077 15487
rect 4077 15453 4111 15487
rect 4111 15453 4120 15487
rect 4068 15444 4120 15453
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 8668 15444 8720 15496
rect 10784 15444 10836 15496
rect 12900 15487 12952 15496
rect 9036 15376 9088 15428
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 12624 15376 12676 15428
rect 17960 15444 18012 15496
rect 3240 15308 3292 15360
rect 4712 15308 4764 15360
rect 5448 15308 5500 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2504 15104 2556 15156
rect 6092 15147 6144 15156
rect 6092 15113 6101 15147
rect 6101 15113 6135 15147
rect 6135 15113 6144 15147
rect 6092 15104 6144 15113
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 9956 15104 10008 15156
rect 12900 15104 12952 15156
rect 16120 15104 16172 15156
rect 10692 15036 10744 15088
rect 2688 14968 2740 15020
rect 3056 15011 3108 15020
rect 3056 14977 3065 15011
rect 3065 14977 3099 15011
rect 3099 14977 3108 15011
rect 3056 14968 3108 14977
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 7380 14968 7432 15020
rect 10508 14968 10560 15020
rect 12256 15036 12308 15088
rect 13268 15036 13320 15088
rect 4068 14900 4120 14952
rect 4344 14900 4396 14952
rect 5540 14900 5592 14952
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 7472 14900 7524 14952
rect 2688 14832 2740 14884
rect 5724 14832 5776 14884
rect 9312 14832 9364 14884
rect 664 14764 716 14816
rect 10784 14764 10836 14816
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 14004 14968 14056 15020
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 16488 15011 16540 15020
rect 16488 14977 16497 15011
rect 16497 14977 16531 15011
rect 16531 14977 16540 15011
rect 16488 14968 16540 14977
rect 19432 14968 19484 15020
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13912 14900 13964 14952
rect 14464 14900 14516 14952
rect 11612 14832 11664 14884
rect 13912 14764 13964 14816
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 15016 14764 15068 14816
rect 18236 14764 18288 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 2964 14560 3016 14612
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 1768 14492 1820 14544
rect 3700 14492 3752 14544
rect 7104 14492 7156 14544
rect 10876 14560 10928 14612
rect 10968 14560 11020 14612
rect 14004 14560 14056 14612
rect 14372 14560 14424 14612
rect 16488 14560 16540 14612
rect 1860 14424 1912 14476
rect 2320 14424 2372 14476
rect 4344 14467 4396 14476
rect 4344 14433 4353 14467
rect 4353 14433 4387 14467
rect 4387 14433 4396 14467
rect 4344 14424 4396 14433
rect 6092 14424 6144 14476
rect 8944 14467 8996 14476
rect 8944 14433 8953 14467
rect 8953 14433 8987 14467
rect 8987 14433 8996 14467
rect 8944 14424 8996 14433
rect 11612 14492 11664 14544
rect 18420 14560 18472 14612
rect 17960 14492 18012 14544
rect 19432 14492 19484 14544
rect 12624 14424 12676 14476
rect 12992 14424 13044 14476
rect 13912 14424 13964 14476
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 15752 14467 15804 14476
rect 15752 14433 15786 14467
rect 15786 14433 15804 14467
rect 15752 14424 15804 14433
rect 5540 14356 5592 14408
rect 6184 14356 6236 14408
rect 8392 14356 8444 14408
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 12532 14399 12584 14408
rect 6920 14220 6972 14272
rect 7656 14263 7708 14272
rect 7656 14229 7665 14263
rect 7665 14229 7699 14263
rect 7699 14229 7708 14263
rect 7656 14220 7708 14229
rect 8576 14263 8628 14272
rect 8576 14229 8585 14263
rect 8585 14229 8619 14263
rect 8619 14229 8628 14263
rect 8576 14220 8628 14229
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 18052 14424 18104 14476
rect 11888 14263 11940 14272
rect 11888 14229 11897 14263
rect 11897 14229 11931 14263
rect 11931 14229 11940 14263
rect 11888 14220 11940 14229
rect 11980 14220 12032 14272
rect 14096 14220 14148 14272
rect 17408 14220 17460 14272
rect 18696 14220 18748 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2688 14016 2740 14068
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 12624 14059 12676 14068
rect 12624 14025 12633 14059
rect 12633 14025 12667 14059
rect 12667 14025 12676 14059
rect 12624 14016 12676 14025
rect 13268 14016 13320 14068
rect 15016 14059 15068 14068
rect 15016 14025 15025 14059
rect 15025 14025 15059 14059
rect 15059 14025 15068 14059
rect 15016 14016 15068 14025
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 2320 13880 2372 13932
rect 5816 13948 5868 14000
rect 7380 13948 7432 14000
rect 5724 13880 5776 13932
rect 6092 13923 6144 13932
rect 6092 13889 6101 13923
rect 6101 13889 6135 13923
rect 6135 13889 6144 13923
rect 6092 13880 6144 13889
rect 7656 13880 7708 13932
rect 10784 13948 10836 14000
rect 11152 13880 11204 13932
rect 11612 13948 11664 14000
rect 3240 13812 3292 13864
rect 5264 13812 5316 13864
rect 6828 13812 6880 13864
rect 7748 13812 7800 13864
rect 9128 13812 9180 13864
rect 11612 13812 11664 13864
rect 12256 13855 12308 13864
rect 12256 13821 12265 13855
rect 12265 13821 12299 13855
rect 12299 13821 12308 13855
rect 12256 13812 12308 13821
rect 13912 13880 13964 13932
rect 15108 13880 15160 13932
rect 15752 14016 15804 14068
rect 18788 14016 18840 14068
rect 18512 13923 18564 13932
rect 18512 13889 18521 13923
rect 18521 13889 18555 13923
rect 18555 13889 18564 13923
rect 18512 13880 18564 13889
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 14556 13812 14608 13864
rect 4896 13787 4948 13796
rect 4896 13753 4905 13787
rect 4905 13753 4939 13787
rect 4939 13753 4948 13787
rect 4896 13744 4948 13753
rect 4988 13744 5040 13796
rect 5356 13744 5408 13796
rect 7380 13744 7432 13796
rect 12808 13744 12860 13796
rect 15292 13744 15344 13796
rect 17684 13812 17736 13864
rect 16396 13744 16448 13796
rect 17960 13744 18012 13796
rect 3700 13676 3752 13728
rect 8944 13676 8996 13728
rect 11152 13676 11204 13728
rect 11980 13676 12032 13728
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 13084 13719 13136 13728
rect 13084 13685 13093 13719
rect 13093 13685 13127 13719
rect 13127 13685 13136 13719
rect 13084 13676 13136 13685
rect 14280 13676 14332 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1400 13472 1452 13524
rect 4160 13472 4212 13524
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5816 13472 5868 13524
rect 6920 13472 6972 13524
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 8576 13472 8628 13524
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 14188 13472 14240 13524
rect 15108 13472 15160 13524
rect 15844 13472 15896 13524
rect 4988 13404 5040 13456
rect 3516 13336 3568 13388
rect 4068 13336 4120 13388
rect 6184 13336 6236 13388
rect 7656 13404 7708 13456
rect 7380 13336 7432 13388
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10232 13336 10284 13388
rect 16580 13404 16632 13456
rect 18696 13404 18748 13456
rect 12808 13379 12860 13388
rect 12808 13345 12842 13379
rect 12842 13345 12860 13379
rect 12808 13336 12860 13345
rect 17684 13379 17736 13388
rect 17684 13345 17693 13379
rect 17693 13345 17727 13379
rect 17727 13345 17736 13379
rect 17684 13336 17736 13345
rect 4252 13268 4304 13320
rect 3700 13200 3752 13252
rect 6092 13268 6144 13320
rect 9312 13268 9364 13320
rect 10048 13268 10100 13320
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 15016 13268 15068 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 16948 13200 17000 13252
rect 6092 13132 6144 13184
rect 8484 13132 8536 13184
rect 12256 13132 12308 13184
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2228 12928 2280 12980
rect 7196 12928 7248 12980
rect 7564 12971 7616 12980
rect 7564 12937 7573 12971
rect 7573 12937 7607 12971
rect 7607 12937 7616 12971
rect 7564 12928 7616 12937
rect 2780 12860 2832 12912
rect 4252 12860 4304 12912
rect 10232 12928 10284 12980
rect 10876 12928 10928 12980
rect 11612 12928 11664 12980
rect 13084 12928 13136 12980
rect 13268 12928 13320 12980
rect 10600 12903 10652 12912
rect 10600 12869 10609 12903
rect 10609 12869 10643 12903
rect 10643 12869 10652 12903
rect 10600 12860 10652 12869
rect 11888 12860 11940 12912
rect 13820 12860 13872 12912
rect 16028 12928 16080 12980
rect 16396 12928 16448 12980
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 18604 12928 18656 12980
rect 6184 12835 6236 12844
rect 6184 12801 6193 12835
rect 6193 12801 6227 12835
rect 6227 12801 6236 12835
rect 6184 12792 6236 12801
rect 6460 12792 6512 12844
rect 9036 12792 9088 12844
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 11336 12835 11388 12844
rect 11336 12801 11345 12835
rect 11345 12801 11379 12835
rect 11379 12801 11388 12835
rect 11336 12792 11388 12801
rect 11980 12792 12032 12844
rect 12808 12792 12860 12844
rect 15016 12792 15068 12844
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 16672 12792 16724 12844
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 3056 12724 3108 12776
rect 3792 12724 3844 12776
rect 8484 12724 8536 12776
rect 8576 12724 8628 12776
rect 3700 12656 3752 12708
rect 11612 12724 11664 12776
rect 10324 12656 10376 12708
rect 10692 12656 10744 12708
rect 11152 12656 11204 12708
rect 14188 12656 14240 12708
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 15660 12656 15712 12708
rect 17132 12656 17184 12708
rect 17960 12656 18012 12708
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 14556 12588 14608 12640
rect 18512 12631 18564 12640
rect 18512 12597 18521 12631
rect 18521 12597 18555 12631
rect 18555 12597 18564 12631
rect 18512 12588 18564 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 3516 12427 3568 12436
rect 3516 12393 3525 12427
rect 3525 12393 3559 12427
rect 3559 12393 3568 12427
rect 3516 12384 3568 12393
rect 1768 12316 1820 12368
rect 3056 12359 3108 12368
rect 3056 12325 3065 12359
rect 3065 12325 3099 12359
rect 3099 12325 3108 12359
rect 3056 12316 3108 12325
rect 3240 12316 3292 12368
rect 4068 12316 4120 12368
rect 6000 12384 6052 12436
rect 7656 12384 7708 12436
rect 9128 12427 9180 12436
rect 9128 12393 9137 12427
rect 9137 12393 9171 12427
rect 9171 12393 9180 12427
rect 9128 12384 9180 12393
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 12992 12384 13044 12436
rect 15292 12384 15344 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 18512 12384 18564 12436
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 5080 12248 5132 12300
rect 6184 12359 6236 12368
rect 6184 12325 6218 12359
rect 6218 12325 6236 12359
rect 6184 12316 6236 12325
rect 14188 12316 14240 12368
rect 15752 12316 15804 12368
rect 17776 12316 17828 12368
rect 7472 12248 7524 12300
rect 12532 12248 12584 12300
rect 13268 12248 13320 12300
rect 13452 12248 13504 12300
rect 14464 12248 14516 12300
rect 15108 12291 15160 12300
rect 15108 12257 15117 12291
rect 15117 12257 15151 12291
rect 15151 12257 15160 12291
rect 15108 12248 15160 12257
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 15936 12248 15988 12300
rect 17132 12248 17184 12300
rect 3608 12180 3660 12232
rect 3792 12180 3844 12232
rect 5816 12180 5868 12232
rect 10324 12223 10376 12232
rect 4896 12044 4948 12096
rect 6552 12044 6604 12096
rect 7380 12044 7432 12096
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 11336 12180 11388 12232
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 11888 12112 11940 12164
rect 18512 12180 18564 12232
rect 19064 12180 19116 12232
rect 8484 12044 8536 12096
rect 12900 12044 12952 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 3148 11840 3200 11892
rect 5080 11840 5132 11892
rect 4896 11772 4948 11824
rect 6828 11772 6880 11824
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 3608 11636 3660 11688
rect 6184 11704 6236 11756
rect 6552 11704 6604 11756
rect 7564 11840 7616 11892
rect 7656 11840 7708 11892
rect 14096 11840 14148 11892
rect 14188 11840 14240 11892
rect 15016 11840 15068 11892
rect 17960 11840 18012 11892
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8576 11704 8628 11756
rect 13452 11747 13504 11756
rect 7932 11636 7984 11688
rect 9864 11636 9916 11688
rect 10600 11636 10652 11688
rect 11060 11636 11112 11688
rect 12072 11636 12124 11688
rect 4804 11568 4856 11620
rect 6092 11611 6144 11620
rect 6092 11577 6101 11611
rect 6101 11577 6135 11611
rect 6135 11577 6144 11611
rect 6092 11568 6144 11577
rect 6276 11568 6328 11620
rect 7748 11568 7800 11620
rect 11612 11568 11664 11620
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 13268 11636 13320 11688
rect 17960 11704 18012 11756
rect 18512 11704 18564 11756
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 5724 11543 5776 11552
rect 5724 11509 5733 11543
rect 5733 11509 5767 11543
rect 5767 11509 5776 11543
rect 5724 11500 5776 11509
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 7472 11500 7524 11552
rect 10784 11500 10836 11552
rect 12624 11500 12676 11552
rect 14188 11568 14240 11620
rect 14556 11568 14608 11620
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 16672 11500 16724 11552
rect 18880 11611 18932 11620
rect 18880 11577 18914 11611
rect 18914 11577 18932 11611
rect 18880 11568 18932 11577
rect 17776 11500 17828 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2780 11296 2832 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 13360 11296 13412 11348
rect 16028 11296 16080 11348
rect 16672 11339 16724 11348
rect 5724 11228 5776 11280
rect 6736 11228 6788 11280
rect 11152 11228 11204 11280
rect 12256 11228 12308 11280
rect 15568 11228 15620 11280
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 17960 11228 18012 11280
rect 2412 11203 2464 11212
rect 2412 11169 2421 11203
rect 2421 11169 2455 11203
rect 2455 11169 2464 11203
rect 2412 11160 2464 11169
rect 5540 11160 5592 11212
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 2596 11135 2648 11144
rect 2596 11101 2605 11135
rect 2605 11101 2639 11135
rect 2639 11101 2648 11135
rect 5080 11135 5132 11144
rect 2596 11092 2648 11101
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 6828 11092 6880 11144
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7748 11024 7800 11076
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 9864 11092 9916 11144
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 11060 11024 11112 11076
rect 11244 11067 11296 11076
rect 11244 11033 11253 11067
rect 11253 11033 11287 11067
rect 11287 11033 11296 11067
rect 11244 11024 11296 11033
rect 12900 11160 12952 11212
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 15752 11160 15804 11212
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 12808 11135 12860 11144
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 13728 11135 13780 11144
rect 12808 11092 12860 11101
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 13636 11024 13688 11076
rect 14556 11092 14608 11144
rect 18604 11160 18656 11212
rect 1768 10956 1820 11008
rect 6092 10956 6144 11008
rect 6828 10956 6880 11008
rect 10324 10956 10376 11008
rect 15660 10956 15712 11008
rect 16028 10956 16080 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 7196 10752 7248 10804
rect 3976 10684 4028 10736
rect 10324 10752 10376 10804
rect 11336 10684 11388 10736
rect 12808 10752 12860 10804
rect 14280 10752 14332 10804
rect 14556 10752 14608 10804
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 1400 10616 1452 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3792 10616 3844 10668
rect 5540 10616 5592 10668
rect 7748 10616 7800 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 3332 10548 3384 10600
rect 7012 10548 7064 10600
rect 9220 10548 9272 10600
rect 3424 10480 3476 10532
rect 10784 10548 10836 10600
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 13268 10616 13320 10668
rect 15016 10616 15068 10668
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 16856 10659 16908 10668
rect 15660 10616 15712 10625
rect 16856 10625 16865 10659
rect 16865 10625 16899 10659
rect 16899 10625 16908 10659
rect 16856 10616 16908 10625
rect 11152 10480 11204 10532
rect 12532 10480 12584 10532
rect 15108 10548 15160 10600
rect 13636 10523 13688 10532
rect 13636 10489 13670 10523
rect 13670 10489 13688 10523
rect 13636 10480 13688 10489
rect 5540 10412 5592 10464
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6000 10412 6052 10464
rect 7380 10412 7432 10464
rect 8576 10412 8628 10464
rect 12716 10412 12768 10464
rect 13268 10412 13320 10464
rect 18696 10548 18748 10600
rect 18604 10480 18656 10532
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 3148 10208 3200 10260
rect 5540 10208 5592 10260
rect 6092 10208 6144 10260
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 3792 10140 3844 10192
rect 2780 10072 2832 10124
rect 3608 10072 3660 10124
rect 3976 10072 4028 10124
rect 6460 10072 6512 10124
rect 6644 10115 6696 10124
rect 6644 10081 6678 10115
rect 6678 10081 6696 10115
rect 6644 10072 6696 10081
rect 8392 10115 8444 10124
rect 8392 10081 8401 10115
rect 8401 10081 8435 10115
rect 8435 10081 8444 10115
rect 8392 10072 8444 10081
rect 10232 10072 10284 10124
rect 11336 10115 11388 10124
rect 11336 10081 11370 10115
rect 11370 10081 11388 10115
rect 11336 10072 11388 10081
rect 2872 10004 2924 10056
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 9588 10004 9640 10056
rect 13636 10208 13688 10260
rect 12992 10183 13044 10192
rect 12992 10149 13004 10183
rect 13004 10149 13044 10183
rect 12992 10140 13044 10149
rect 16856 10140 16908 10192
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 2596 9868 2648 9920
rect 3884 9868 3936 9920
rect 8024 9911 8076 9920
rect 8024 9877 8033 9911
rect 8033 9877 8067 9911
rect 8067 9877 8076 9911
rect 8024 9868 8076 9877
rect 15384 9868 15436 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3424 9664 3476 9716
rect 1676 9596 1728 9648
rect 3976 9596 4028 9648
rect 5724 9664 5776 9716
rect 3792 9528 3844 9580
rect 9588 9596 9640 9648
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 13728 9596 13780 9648
rect 6644 9528 6696 9580
rect 12992 9571 13044 9580
rect 4712 9460 4764 9512
rect 3056 9392 3108 9444
rect 3792 9392 3844 9444
rect 7196 9460 7248 9512
rect 8024 9460 8076 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9128 9460 9180 9512
rect 12992 9537 13001 9571
rect 13001 9537 13035 9571
rect 13035 9537 13044 9571
rect 12992 9528 13044 9537
rect 16028 9664 16080 9716
rect 16856 9664 16908 9716
rect 16672 9528 16724 9580
rect 12532 9460 12584 9512
rect 14004 9460 14056 9512
rect 15016 9460 15068 9512
rect 15660 9503 15712 9512
rect 15660 9469 15694 9503
rect 15694 9469 15712 9503
rect 15660 9460 15712 9469
rect 6736 9392 6788 9444
rect 8484 9392 8536 9444
rect 12348 9392 12400 9444
rect 2504 9367 2556 9376
rect 2504 9333 2513 9367
rect 2513 9333 2547 9367
rect 2547 9333 2556 9367
rect 2504 9324 2556 9333
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3608 9324 3660 9376
rect 4804 9324 4856 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 7472 9324 7524 9376
rect 9312 9324 9364 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 2504 9120 2556 9172
rect 7196 9120 7248 9172
rect 8392 9163 8444 9172
rect 8392 9129 8401 9163
rect 8401 9129 8435 9163
rect 8435 9129 8444 9163
rect 8392 9120 8444 9129
rect 2872 9095 2924 9104
rect 2872 9061 2881 9095
rect 2881 9061 2915 9095
rect 2915 9061 2924 9095
rect 2872 9052 2924 9061
rect 4068 9052 4120 9104
rect 18972 9052 19024 9104
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 8760 9027 8812 9036
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 8760 8984 8812 8993
rect 9404 8984 9456 9036
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 5356 8916 5408 8968
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 8668 8916 8720 8968
rect 8852 8959 8904 8968
rect 8852 8925 8861 8959
rect 8861 8925 8895 8959
rect 8895 8925 8904 8959
rect 8852 8916 8904 8925
rect 9128 8916 9180 8968
rect 2412 8848 2464 8900
rect 4160 8848 4212 8900
rect 8760 8848 8812 8900
rect 3976 8780 4028 8832
rect 15292 8780 15344 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2780 8576 2832 8628
rect 3056 8576 3108 8628
rect 7380 8576 7432 8628
rect 9128 8576 9180 8628
rect 5448 8508 5500 8560
rect 3148 8440 3200 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4712 8440 4764 8492
rect 7748 8440 7800 8492
rect 1860 8372 1912 8424
rect 2596 8372 2648 8424
rect 4160 8347 4212 8356
rect 4160 8313 4169 8347
rect 4169 8313 4203 8347
rect 4203 8313 4212 8347
rect 4160 8304 4212 8313
rect 6920 8372 6972 8424
rect 7196 8347 7248 8356
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 7196 8313 7205 8347
rect 7205 8313 7239 8347
rect 7239 8313 7248 8347
rect 7196 8304 7248 8313
rect 7288 8347 7340 8356
rect 7288 8313 7297 8347
rect 7297 8313 7331 8347
rect 7331 8313 7340 8347
rect 7288 8304 7340 8313
rect 8576 8304 8628 8356
rect 7012 8236 7064 8288
rect 13544 8236 13596 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3148 7964 3200 8016
rect 4804 8032 4856 8084
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 7012 8032 7064 8084
rect 7748 8032 7800 8084
rect 11796 8032 11848 8084
rect 6920 7964 6972 8016
rect 7472 7964 7524 8016
rect 7656 7964 7708 8016
rect 1860 7939 1912 7948
rect 1860 7905 1869 7939
rect 1869 7905 1903 7939
rect 1903 7905 1912 7939
rect 1860 7896 1912 7905
rect 3976 7896 4028 7948
rect 19340 8032 19392 8084
rect 4344 7760 4396 7812
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 4804 7760 4856 7812
rect 5080 7735 5132 7744
rect 3240 7692 3292 7701
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 6092 7692 6144 7744
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 19524 7531 19576 7540
rect 19524 7497 19533 7531
rect 19533 7497 19567 7531
rect 19567 7497 19576 7531
rect 19524 7488 19576 7497
rect 6368 7420 6420 7472
rect 6828 7420 6880 7472
rect 8300 7420 8352 7472
rect 1860 7284 1912 7336
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 6000 7352 6052 7404
rect 8944 7352 8996 7404
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 2964 7216 3016 7268
rect 3240 7216 3292 7268
rect 5724 7216 5776 7268
rect 7748 7216 7800 7268
rect 12348 7216 12400 7268
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 5080 7148 5132 7200
rect 6000 7148 6052 7200
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 7564 7148 7616 7200
rect 8300 7148 8352 7200
rect 12440 7148 12492 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 2964 6987 3016 6996
rect 2964 6953 2973 6987
rect 2973 6953 3007 6987
rect 3007 6953 3016 6987
rect 2964 6944 3016 6953
rect 3608 6944 3660 6996
rect 6828 6944 6880 6996
rect 7012 6944 7064 6996
rect 2872 6876 2924 6928
rect 5724 6876 5776 6928
rect 6000 6876 6052 6928
rect 6276 6876 6328 6928
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 4528 6808 4580 6860
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 1768 6740 1820 6792
rect 3148 6740 3200 6792
rect 3240 6672 3292 6724
rect 3148 6604 3200 6656
rect 5356 6672 5408 6724
rect 6920 6672 6972 6724
rect 7656 6740 7708 6792
rect 7196 6672 7248 6724
rect 19892 6715 19944 6724
rect 19892 6681 19901 6715
rect 19901 6681 19935 6715
rect 19935 6681 19944 6715
rect 19892 6672 19944 6681
rect 3884 6604 3936 6656
rect 20996 6672 21048 6724
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 7288 6400 7340 6452
rect 20904 6400 20956 6452
rect 4068 6332 4120 6384
rect 19708 6332 19760 6384
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 7564 6196 7616 6248
rect 4712 6128 4764 6180
rect 8392 6060 8444 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 3700 5312 3752 5364
rect 12624 5312 12676 5364
rect 20812 5312 20864 5364
rect 4068 5108 4120 5160
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 5724 4088 5776 4140
rect 10140 4088 10192 4140
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 3332 1300 3384 1352
rect 6092 1300 6144 1352
rect 16580 552 16632 604
rect 17132 552 17184 604
<< metal2 >>
rect 202 22320 258 22800
rect 662 22320 718 22800
rect 1122 22320 1178 22800
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 216 19242 244 22320
rect 204 19236 256 19242
rect 204 19178 256 19184
rect 676 14822 704 22320
rect 1136 18154 1164 22320
rect 1124 18148 1176 18154
rect 1124 18090 1176 18096
rect 664 14816 716 14822
rect 664 14758 716 14764
rect 1412 13530 1440 22471
rect 1582 22320 1638 22800
rect 2042 22320 2098 22800
rect 2502 22320 2558 22800
rect 2962 22320 3018 22800
rect 3422 22320 3478 22800
rect 3882 22320 3938 22800
rect 4342 22320 4398 22800
rect 4802 22320 4858 22800
rect 5262 22320 5318 22800
rect 5722 22320 5778 22800
rect 6182 22320 6238 22800
rect 6642 22320 6698 22800
rect 7102 22320 7158 22800
rect 7562 22320 7618 22800
rect 8114 22320 8170 22800
rect 8574 22320 8630 22800
rect 9034 22320 9090 22800
rect 9494 22320 9550 22800
rect 9954 22320 10010 22800
rect 10414 22320 10470 22800
rect 10874 22320 10930 22800
rect 11334 22320 11390 22800
rect 11794 22320 11850 22800
rect 12254 22320 12310 22800
rect 12714 22320 12770 22800
rect 13174 22320 13230 22800
rect 13634 22320 13690 22800
rect 14094 22320 14150 22800
rect 14554 22320 14610 22800
rect 15014 22320 15070 22800
rect 15566 22320 15622 22800
rect 16026 22320 16082 22800
rect 16486 22320 16542 22800
rect 16946 22320 17002 22800
rect 17406 22320 17462 22800
rect 17866 22320 17922 22800
rect 18326 22320 18382 22800
rect 18786 22320 18842 22800
rect 19246 22320 19302 22800
rect 19706 22320 19762 22800
rect 20166 22320 20222 22800
rect 20626 22320 20682 22800
rect 21086 22320 21142 22800
rect 21546 22320 21602 22800
rect 22006 22320 22062 22800
rect 22466 22320 22522 22800
rect 1596 19394 1624 22320
rect 1674 20632 1730 20641
rect 1674 20567 1730 20576
rect 1504 19366 1624 19394
rect 1504 18766 1532 19366
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1596 18290 1624 19246
rect 1688 19174 1716 20567
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 19378 1808 19858
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1950 18320 2006 18329
rect 1584 18284 1636 18290
rect 1950 18255 2006 18264
rect 1584 18226 1636 18232
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17377 1624 18022
rect 1964 17882 1992 18255
rect 2056 18193 2084 22320
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2226 19272 2282 19281
rect 2226 19207 2282 19216
rect 2042 18184 2098 18193
rect 2042 18119 2098 18128
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1582 17368 1638 17377
rect 1582 17303 1638 17312
rect 1676 16992 1728 16998
rect 1674 16960 1676 16969
rect 1728 16960 1730 16969
rect 1674 16895 1730 16904
rect 1780 16590 1808 17682
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2056 16794 2084 17070
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1768 16584 1820 16590
rect 1582 16552 1638 16561
rect 1768 16526 1820 16532
rect 1582 16487 1638 16496
rect 1596 16250 1624 16487
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 2056 16114 2084 16594
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1964 15706 1992 15943
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1674 14648 1730 14657
rect 1674 14583 1730 14592
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1400 13524 1452 13530
rect 1400 13466 1452 13472
rect 1596 11898 1624 13631
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 10674 1440 11630
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1688 9654 1716 14583
rect 1780 14550 1808 15506
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1860 14476 1912 14482
rect 1860 14418 1912 14424
rect 1872 13938 1900 14418
rect 1950 14104 2006 14113
rect 1950 14039 2006 14048
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 12374 1808 12718
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10606 1808 10950
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1964 9178 1992 14039
rect 2240 12986 2268 19207
rect 2332 18902 2360 19858
rect 2516 19514 2544 22320
rect 2870 21584 2926 21593
rect 2870 21519 2926 21528
rect 2778 21176 2834 21185
rect 2778 21111 2834 21120
rect 2792 20058 2820 21111
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2778 19816 2834 19825
rect 2884 19786 2912 21519
rect 2976 20346 3004 22320
rect 3238 22128 3294 22137
rect 3238 22063 3294 22072
rect 2976 20318 3188 20346
rect 3054 20224 3110 20233
rect 3054 20159 3110 20168
rect 2778 19751 2834 19760
rect 2872 19780 2924 19786
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2410 19272 2466 19281
rect 2410 19207 2412 19216
rect 2464 19207 2466 19216
rect 2412 19178 2464 19184
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2424 18358 2452 18770
rect 2688 18760 2740 18766
rect 2686 18728 2688 18737
rect 2740 18728 2742 18737
rect 2686 18663 2742 18672
rect 2412 18352 2464 18358
rect 2318 18320 2374 18329
rect 2412 18294 2464 18300
rect 2318 18255 2374 18264
rect 2332 18222 2360 18255
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2792 18034 2820 19751
rect 2872 19722 2924 19728
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 2976 19310 3004 19654
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 2962 18864 3018 18873
rect 2962 18799 3018 18808
rect 2792 18006 2912 18034
rect 2778 17912 2834 17921
rect 2778 17847 2780 17856
rect 2832 17847 2834 17856
rect 2780 17818 2832 17824
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2424 17202 2452 17682
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2884 16250 2912 18006
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2332 14482 2360 15438
rect 2516 15162 2544 15982
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2700 15026 2728 15982
rect 2778 15600 2834 15609
rect 2778 15535 2834 15544
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 2332 13938 2360 14418
rect 2700 14074 2728 14826
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2792 12918 2820 15535
rect 2884 14498 2912 15982
rect 2976 14618 3004 18799
rect 3068 17882 3096 20159
rect 3160 19310 3188 20318
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3160 17882 3188 18770
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3252 16726 3280 22063
rect 3436 18873 3464 22320
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 3792 19168 3844 19174
rect 3792 19110 3844 19116
rect 3422 18864 3478 18873
rect 3422 18799 3478 18808
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3344 17746 3372 18702
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3620 18193 3648 18362
rect 3712 18358 3740 19110
rect 3804 18766 3832 19110
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 3606 18184 3662 18193
rect 3516 18148 3568 18154
rect 3606 18119 3662 18128
rect 3516 18090 3568 18096
rect 3528 18034 3556 18090
rect 3712 18034 3740 18294
rect 3804 18222 3832 18702
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3528 18006 3740 18034
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3344 17134 3372 17682
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3896 16810 3924 22320
rect 4356 19802 4384 22320
rect 4172 19774 4384 19802
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4080 17746 4108 18022
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3344 16782 3924 16810
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15026 3096 15846
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3146 15056 3202 15065
rect 3056 15020 3108 15026
rect 3252 15026 3280 15302
rect 3146 14991 3202 15000
rect 3240 15020 3292 15026
rect 3056 14962 3108 14968
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2884 14470 3004 14498
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11354 2820 12242
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1780 6798 1808 8978
rect 2424 8906 2452 11154
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2516 10810 2544 11086
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2608 9926 2636 11086
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2516 9178 2544 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2608 8430 2636 9862
rect 2792 8634 2820 10066
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 9110 2912 9998
rect 2976 9382 3004 14470
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3068 12374 3096 12718
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 3160 11898 3188 14991
rect 3240 14962 3292 14968
rect 3252 13870 3280 14962
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10266 3188 10610
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 1872 7954 1900 8366
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1872 7342 1900 7890
rect 2976 7392 3004 9318
rect 3068 8634 3096 9386
rect 3160 8974 3188 10202
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2884 7364 3004 7392
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1872 6866 1900 7142
rect 2884 6934 2912 7364
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2976 7002 3004 7210
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 2884 2961 2912 6870
rect 3068 3913 3096 8570
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3160 8294 3188 8434
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3160 8022 3188 8230
rect 3252 8129 3280 12310
rect 3344 10606 3372 16782
rect 4080 16114 4108 16934
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15638 4108 16050
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4080 14958 4108 15438
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3712 13818 3740 14486
rect 3620 13790 3740 13818
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 12442 3556 13330
rect 3620 12594 3648 13790
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3712 13258 3740 13670
rect 4172 13530 4200 19774
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4724 19174 4752 19790
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4264 13410 4292 18770
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4724 18222 4752 18294
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4724 17134 4752 18158
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4724 16046 4752 17070
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4540 15638 4568 15982
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4724 15366 4752 15982
rect 4816 15910 4844 22320
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5092 18222 5120 19246
rect 5276 18970 5304 22320
rect 5736 20058 5764 22320
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5736 18766 5764 19178
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5184 18329 5212 18634
rect 5170 18320 5226 18329
rect 5170 18255 5226 18264
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5552 17882 5580 18702
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5920 17678 5948 18090
rect 6196 17882 6224 22320
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5828 17338 5856 17478
rect 5920 17338 5948 17614
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 5276 16590 5304 17002
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 16250 5304 16526
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 5552 15706 5580 16594
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6104 15978 6132 16526
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4356 14482 4384 14894
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4908 13802 4936 15438
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15178 5488 15302
rect 5460 15150 5580 15178
rect 6104 15162 6132 15914
rect 5552 14958 5580 15150
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5552 14414 5580 14894
rect 5724 14884 5776 14890
rect 5724 14826 5776 14832
rect 5736 14618 5764 14826
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5736 13938 5764 14554
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5000 13462 5028 13738
rect 5276 13530 5304 13806
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4172 13382 4292 13410
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3712 12714 3740 13194
rect 3792 12776 3844 12782
rect 4080 12753 4108 13330
rect 3792 12718 3844 12724
rect 4066 12744 4122 12753
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3620 12566 3740 12594
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3620 11694 3648 12174
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 9722 3464 10474
rect 3620 10130 3648 11630
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3238 8120 3294 8129
rect 3238 8055 3294 8064
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7274 3280 7686
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3160 6662 3188 6734
rect 3252 6730 3280 7210
rect 3620 7002 3648 9318
rect 3712 8537 3740 12566
rect 3804 12238 3832 12718
rect 4066 12679 4122 12688
rect 4068 12368 4120 12374
rect 4066 12336 4068 12345
rect 4120 12336 4122 12345
rect 4066 12271 4122 12280
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3974 10840 4030 10849
rect 3974 10775 4030 10784
rect 3988 10742 4016 10775
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3804 10198 3832 10610
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3804 9586 3832 10134
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3792 9444 3844 9450
rect 3792 9386 3844 9392
rect 3698 8528 3754 8537
rect 3698 8463 3754 8472
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3054 3904 3110 3913
rect 3054 3839 3110 3848
rect 3160 3505 3188 6598
rect 3620 5522 3648 6938
rect 3804 5658 3832 9386
rect 3896 7585 3924 9862
rect 3988 9654 4016 10066
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3974 9480 4030 9489
rect 3974 9415 4030 9424
rect 3988 8838 4016 9415
rect 4068 9104 4120 9110
rect 4066 9072 4068 9081
rect 4120 9072 4122 9081
rect 4066 9007 4122 9016
rect 4172 8906 4200 13382
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 12918 4292 13262
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4252 12912 4304 12918
rect 4252 12854 4304 12860
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4908 11830 4936 12038
rect 5092 11898 5120 12242
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4804 11620 4856 11626
rect 4804 11562 4856 11568
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4250 8936 4306 8945
rect 4160 8900 4212 8906
rect 4250 8871 4306 8880
rect 4160 8842 4212 8848
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 4172 8362 4200 8842
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3882 7576 3938 7585
rect 3882 7511 3938 7520
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 5817 3924 6598
rect 3882 5808 3938 5817
rect 3882 5743 3938 5752
rect 3804 5630 3924 5658
rect 3620 5494 3832 5522
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3712 4321 3740 5306
rect 3698 4312 3754 4321
rect 3698 4247 3754 4256
rect 3146 3496 3202 3505
rect 3146 3431 3202 3440
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 3804 2009 3832 5494
rect 3790 2000 3846 2009
rect 3790 1935 3846 1944
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 241 3372 1294
rect 3896 1057 3924 5630
rect 3882 1048 3938 1057
rect 3882 983 3938 992
rect 3988 649 4016 7890
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4080 6225 4108 6326
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4865 4108 5102
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 4172 2553 4200 8298
rect 4264 8294 4292 8871
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8498 4752 9454
rect 4816 9382 4844 11562
rect 5092 11150 5120 11834
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 5368 8974 5396 13738
rect 5828 13530 5856 13942
rect 6104 13938 6132 14418
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6092 13932 6144 13938
rect 6012 13892 6092 13920
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6012 12442 6040 13892
rect 6092 13874 6144 13880
rect 6196 13818 6224 14350
rect 6104 13790 6224 13818
rect 6104 13326 6132 13790
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6104 12356 6132 13126
rect 6196 12850 6224 13330
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6184 12368 6236 12374
rect 6104 12328 6184 12356
rect 6184 12310 6236 12316
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5736 11286 5764 11494
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10674 5580 11154
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5724 10464 5776 10470
rect 5828 10452 5856 12174
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6012 10470 6040 11086
rect 6104 11014 6132 11562
rect 6196 11150 6224 11698
rect 6288 11626 6316 18022
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 5776 10424 5856 10452
rect 6000 10464 6052 10470
rect 5724 10406 5776 10412
rect 6000 10406 6052 10412
rect 5552 10266 5580 10406
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5736 9722 5764 10406
rect 6104 10266 6132 10950
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4158 2544 4214 2553
rect 4158 2479 4214 2488
rect 4264 1601 4292 8230
rect 4356 7818 4384 8434
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4816 7818 4844 8026
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4540 6866 4568 7278
rect 5092 7206 5120 7686
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 5368 6730 5396 8910
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5460 8090 5488 8502
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 6104 7750 6132 10202
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5736 6934 5764 7210
rect 6012 7206 6040 7346
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6012 6934 6040 7142
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4724 5273 4752 6122
rect 4710 5264 4766 5273
rect 4710 5199 4766 5208
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4250 1592 4306 1601
rect 4250 1527 4306 1536
rect 3974 640 4030 649
rect 3974 575 4030 584
rect 5736 480 5764 4082
rect 6104 1358 6132 7686
rect 6380 7478 6408 19858
rect 6460 19848 6512 19854
rect 6460 19790 6512 19796
rect 6472 19514 6500 19790
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6472 19242 6500 19450
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6472 18358 6500 18702
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6656 16794 6684 22320
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6748 18970 6776 19246
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 7116 18034 7144 22320
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7208 19242 7236 19450
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 7392 18290 7420 19246
rect 7470 18864 7526 18873
rect 7470 18799 7526 18808
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 6840 18006 7144 18034
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6840 13870 6868 18006
rect 7392 17338 7420 18226
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6932 16046 6960 17002
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6932 15706 6960 15846
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7024 15570 7052 17070
rect 7392 16658 7420 17274
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7116 16250 7144 16594
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7116 15994 7144 16186
rect 7392 16046 7420 16594
rect 7380 16040 7432 16046
rect 7116 15966 7328 15994
rect 7380 15982 7432 15988
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7024 15162 7052 15506
rect 7208 15502 7236 15846
rect 7196 15496 7248 15502
rect 7116 15456 7196 15484
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7116 14550 7144 15456
rect 7196 15438 7248 15444
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6932 13530 6960 14214
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6458 13288 6514 13297
rect 6458 13223 6514 13232
rect 6472 12850 6500 13223
rect 7208 12986 7236 14894
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11762 6592 12038
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6734 11384 6790 11393
rect 6840 11354 6868 11766
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6734 11319 6790 11328
rect 6828 11348 6880 11354
rect 6748 11286 6776 11319
rect 6828 11290 6880 11296
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6840 11014 6868 11086
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 7024 10606 7052 11494
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7208 10810 7236 11154
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6472 8378 6500 10066
rect 6656 9586 6684 10066
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 7196 9512 7248 9518
rect 7300 9500 7328 15966
rect 7392 15026 7420 15982
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7392 14006 7420 14962
rect 7484 14958 7512 18799
rect 7576 18086 7604 22320
rect 8128 20346 8156 22320
rect 7760 20318 8156 20346
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7668 13938 7696 14214
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13394 7420 13738
rect 7668 13462 7696 13874
rect 7760 13870 7788 20318
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8588 18204 8616 22320
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8772 18970 8800 19110
rect 8864 18970 8892 19654
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 9048 18290 9076 22320
rect 9508 20058 9536 22320
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9586 19272 9642 19281
rect 9496 19236 9548 19242
rect 9586 19207 9588 19216
rect 9496 19178 9548 19184
rect 9640 19207 9642 19216
rect 9588 19178 9640 19184
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9128 18760 9180 18766
rect 9126 18728 9128 18737
rect 9180 18728 9182 18737
rect 9126 18663 9182 18672
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8220 18176 8616 18204
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 7944 17202 7972 17682
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15706 8248 18176
rect 9416 18086 9444 18770
rect 9508 18630 9536 19178
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9600 18170 9628 18770
rect 9692 18290 9720 19110
rect 9876 18902 9904 19654
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9772 18216 9824 18222
rect 9600 18164 9772 18170
rect 9600 18158 9824 18164
rect 9600 18142 9812 18158
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 8772 17678 8800 18022
rect 9048 17882 9076 18022
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9784 17814 9812 18142
rect 9968 17882 9996 22320
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10336 18222 10364 19790
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10428 18086 10456 22320
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9416 17678 9444 17750
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8760 17672 8812 17678
rect 8760 17614 8812 17620
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 8312 16726 8340 17614
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8680 15978 8708 16390
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8680 15502 8708 15914
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 8404 13530 8432 14350
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8588 13530 8616 14214
rect 8956 13734 8984 14418
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11762 7420 12038
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7484 11558 7512 12242
rect 7576 11898 7604 12922
rect 8496 12782 8524 13126
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 11898 7696 12378
rect 8484 12096 8536 12102
rect 8588 12050 8616 12718
rect 8536 12044 8616 12050
rect 8484 12038 8616 12044
rect 8496 12022 8616 12038
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7930 11792 7986 11801
rect 8588 11762 8616 12022
rect 7930 11727 7986 11736
rect 8576 11756 8628 11762
rect 7944 11694 7972 11727
rect 8576 11698 8628 11704
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11150 7512 11494
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7760 11082 7788 11562
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7760 10674 7788 11018
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7248 9472 7328 9500
rect 7196 9454 7248 9460
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 8974 6776 9386
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 9178 7236 9318
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7392 8634 7420 10406
rect 7760 10266 7788 10610
rect 8588 10470 8616 11698
rect 8576 10464 8628 10470
rect 8576 10406 8628 10412
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 9518 8064 9862
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 6920 8424 6972 8430
rect 6748 8384 6920 8412
rect 6748 8378 6776 8384
rect 6472 8350 6776 8378
rect 6920 8366 6972 8372
rect 7196 8356 7248 8362
rect 6564 7886 6592 8350
rect 7196 8298 7248 8304
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 8090 7052 8230
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6934 6316 7142
rect 6840 7002 6868 7414
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6932 6730 6960 7958
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7024 7002 7052 7142
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 7208 6730 7236 8298
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7300 6458 7328 8298
rect 7392 7342 7420 8570
rect 7484 8022 7512 9318
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8404 9178 8432 10066
rect 8588 9518 8616 10406
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8484 9444 8536 9450
rect 8484 9386 8536 9392
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7760 8090 7788 8434
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7564 7200 7616 7206
rect 7668 7177 7696 7958
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7564 7142 7616 7148
rect 7654 7168 7710 7177
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7576 6254 7604 7142
rect 7654 7103 7710 7112
rect 7656 6792 7708 6798
rect 7760 6769 7788 7210
rect 8312 7206 8340 7414
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7656 6734 7708 6740
rect 7746 6760 7802 6769
rect 7668 6322 7696 6734
rect 7746 6695 7802 6704
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 8404 6118 8432 7686
rect 8496 7342 8524 9386
rect 8588 8362 8616 9454
rect 8680 8974 8708 9998
rect 8956 9761 8984 13670
rect 9048 12850 9076 15370
rect 9312 14884 9364 14890
rect 9312 14826 9364 14832
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9140 13870 9168 14350
rect 9324 14074 9352 14826
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9140 12442 9168 13806
rect 9324 13326 9352 14010
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9232 10033 9260 10542
rect 9218 10024 9274 10033
rect 9218 9959 9274 9968
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 9310 9616 9366 9625
rect 9310 9551 9366 9560
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8772 8906 8800 8978
rect 9140 8974 9168 9454
rect 9324 9382 9352 9551
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 9416 9042 9444 17614
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9692 15706 9720 17070
rect 9784 16658 9812 17750
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 17338 9996 17682
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10428 17202 10456 17478
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9968 15162 9996 15982
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15706 10088 15846
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10520 15026 10548 19246
rect 10600 18148 10652 18154
rect 10600 18090 10652 18096
rect 10612 17678 10640 18090
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10612 16794 10640 17614
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10796 16250 10824 16594
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10796 15502 10824 16186
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9508 12668 9812 12696
rect 9508 10577 9536 12668
rect 9784 12617 9812 12668
rect 9770 12608 9826 12617
rect 9770 12543 9826 12552
rect 10060 12442 10088 13262
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 11150 9904 11630
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9494 10568 9550 10577
rect 9494 10503 9550 10512
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9654 9628 9998
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 8852 8968 8904 8974
rect 8850 8936 8852 8945
rect 9128 8968 9180 8974
rect 8904 8936 8906 8945
rect 8760 8900 8812 8906
rect 9128 8910 9180 8916
rect 8850 8871 8906 8880
rect 8760 8842 8812 8848
rect 9140 8634 9168 8910
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7410 8984 7822
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 10152 4146 10180 13330
rect 10244 12986 10272 13330
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 10600 12912 10652 12918
rect 10598 12880 10600 12889
rect 10652 12880 10654 12889
rect 10598 12815 10654 12824
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10336 12238 10364 12650
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10612 11694 10640 12815
rect 10704 12714 10732 15030
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14498 10824 14758
rect 10888 14618 10916 22320
rect 11348 19802 11376 22320
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11164 19774 11376 19802
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10980 17134 11008 17614
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 11072 15994 11100 19246
rect 11164 18766 11192 19774
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11624 18850 11652 19858
rect 11808 19174 11836 22320
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11716 18970 11744 19110
rect 12268 18986 12296 22320
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 11704 18964 11756 18970
rect 11704 18906 11756 18912
rect 11808 18958 12296 18986
rect 11624 18822 11744 18850
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18222 11192 18566
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11716 18086 11744 18822
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11164 16114 11192 18022
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11716 17202 11744 18022
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11072 15966 11192 15994
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15706 11100 15846
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10980 14498 11008 14554
rect 10796 14470 11008 14498
rect 10796 14006 10824 14470
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 11164 13938 11192 15966
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11624 14550 11652 14826
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11624 14006 11652 14486
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10888 12730 10916 12922
rect 11164 12850 11192 13670
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11624 12986 11652 13806
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 10888 12714 11192 12730
rect 10692 12708 10744 12714
rect 10888 12708 11204 12714
rect 10888 12702 11152 12708
rect 10692 12650 10744 12656
rect 11152 12650 11204 12656
rect 11348 12238 11376 12786
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 12458 11652 12718
rect 11624 12430 11744 12458
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10796 11150 10824 11494
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10810 10364 10950
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10796 10606 10824 11086
rect 11072 11082 11100 11630
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 11164 10538 11192 11222
rect 11624 11218 11652 11562
rect 11716 11218 11744 12430
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11242 11112 11298 11121
rect 11242 11047 11244 11056
rect 11296 11047 11298 11056
rect 11244 11018 11296 11024
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11348 10130 11376 10678
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 10244 9654 10272 10066
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11808 8090 11836 18958
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11992 18737 12020 18838
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12072 18760 12124 18766
rect 11978 18728 12034 18737
rect 11888 18692 11940 18698
rect 12072 18702 12124 18708
rect 11978 18663 12034 18672
rect 11888 18634 11940 18640
rect 11900 14362 11928 18634
rect 11900 14334 12020 14362
rect 11992 14278 12020 14334
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11900 12918 11928 14214
rect 11992 13734 12020 14214
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11978 12880 12034 12889
rect 11978 12815 11980 12824
rect 12032 12815 12034 12824
rect 11980 12786 12032 12792
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12170 11928 12582
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 12084 11694 12112 18702
rect 12176 12458 12204 18770
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12268 17814 12296 18158
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15094 12296 15846
rect 12256 15088 12308 15094
rect 12256 15030 12308 15036
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12268 13190 12296 13806
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12176 12430 12287 12458
rect 12259 12424 12287 12430
rect 12259 12396 12296 12424
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12268 11286 12296 12396
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12360 9450 12388 19110
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12452 18222 12480 18702
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12452 17202 12480 18158
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12452 16998 12480 17138
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12544 16794 12572 18770
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12636 16674 12664 19246
rect 12728 17338 12756 22320
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12820 18902 12848 19858
rect 13188 19174 13216 22320
rect 13648 20058 13676 22320
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 14108 19938 14136 22320
rect 13820 19916 13872 19922
rect 14108 19910 14228 19938
rect 13820 19858 13872 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12544 16646 12664 16674
rect 12716 16652 12768 16658
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12452 15706 12480 16526
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 15026 12480 15506
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12544 14414 12572 16646
rect 12716 16594 12768 16600
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12636 15434 12664 15914
rect 12728 15638 12756 16594
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12636 14074 12664 14418
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12820 13802 12848 17682
rect 13004 17678 13032 18090
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 16998 13032 17614
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12912 15978 12940 16934
rect 13096 16590 13124 17002
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 13096 16250 13124 16526
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13280 16046 13308 17070
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12912 15586 12940 15914
rect 12912 15558 13032 15586
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12912 15162 12940 15438
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13004 14482 13032 15558
rect 13280 15094 13308 15982
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 13280 14074 13308 14894
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12544 12306 12572 13262
rect 12820 12850 12848 13330
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12730 12848 12786
rect 12820 12702 12940 12730
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12912 12102 12940 12702
rect 13004 12442 13032 13670
rect 13096 12986 13124 13670
rect 13280 12986 13308 14010
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 13280 11694 13308 12242
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12544 9518 12572 10474
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12348 9444 12400 9450
rect 12348 9386 12400 9392
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 12360 7274 12480 7290
rect 12348 7268 12480 7274
rect 12400 7262 12480 7268
rect 12348 7210 12400 7216
rect 12452 7206 12480 7262
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 12636 5370 12664 11494
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12716 11144 12768 11150
rect 12714 11112 12716 11121
rect 12808 11144 12860 11150
rect 12768 11112 12770 11121
rect 12808 11086 12860 11092
rect 12714 11047 12770 11056
rect 12820 10810 12848 11086
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12912 10674 12940 11154
rect 13280 10674 13308 11630
rect 13372 11354 13400 19790
rect 13832 19514 13860 19858
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13832 18834 13860 19314
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 18086 13860 18770
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17678 13860 18022
rect 13924 17882 13952 19246
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18358 14044 19110
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14108 18222 14136 19790
rect 14200 18426 14228 19910
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14292 17882 14320 19110
rect 14568 18970 14596 22320
rect 15028 20618 15056 22320
rect 15028 20590 15240 20618
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 15212 20058 15240 20590
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14370 18728 14426 18737
rect 14370 18663 14426 18672
rect 14384 18222 14412 18663
rect 15028 18630 15056 19314
rect 15212 18902 15240 19858
rect 15580 19786 15608 22320
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 14384 17338 14412 18158
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17882 14596 18022
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13464 11762 13492 12242
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13280 10470 13308 10610
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 12728 10062 12756 10406
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 13004 9586 13032 10134
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 13556 8294 13584 17274
rect 14384 16402 14412 17274
rect 15028 17134 15056 18566
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14200 16374 14412 16402
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14108 15706 14136 15846
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14822 13952 14894
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 14016 14618 14044 14962
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13924 13938 13952 14418
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13924 13530 13952 13874
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13832 12646 13860 12854
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13648 10538 13676 11018
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13648 10266 13676 10474
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 9654 13768 11086
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 14016 9518 14044 14554
rect 14108 14278 14136 14758
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14200 13530 14228 16374
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 15638 14412 16050
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14384 15026 14412 15574
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14618 14412 14962
rect 14476 14958 14504 15846
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14568 13870 14596 16934
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 15028 14074 15056 14758
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15120 13938 15148 18090
rect 15212 17814 15240 18226
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15488 16250 15516 17002
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14188 13524 14240 13530
rect 14188 13466 14240 13472
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12714 14228 13126
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11898 14136 12174
rect 14200 11898 14228 12310
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14200 11626 14228 11834
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14292 10810 14320 13670
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15120 13530 15148 13874
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 15028 12850 15056 13262
rect 15304 12850 15332 13738
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14384 12702 14596 12730
rect 14384 12617 14412 12702
rect 14568 12646 14596 12702
rect 14464 12640 14516 12646
rect 14370 12608 14426 12617
rect 14464 12582 14516 12588
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14370 12543 14426 12552
rect 14476 12306 14504 12582
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 15028 11898 15056 12786
rect 15304 12442 15332 12786
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15304 12306 15332 12378
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14568 11150 14596 11562
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14568 10810 14596 11086
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 15028 9518 15056 10610
rect 15120 10606 15148 12242
rect 15108 10600 15160 10606
rect 15396 10554 15424 15846
rect 15488 15570 15516 16186
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15488 14482 15516 15506
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15580 11286 15608 18770
rect 15660 18692 15712 18698
rect 15660 18634 15712 18640
rect 15672 17882 15700 18634
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15660 17672 15712 17678
rect 15764 17660 15792 19246
rect 16040 19174 16068 22320
rect 16500 20074 16528 22320
rect 16500 20058 16620 20074
rect 16500 20052 16632 20058
rect 16500 20046 16580 20052
rect 16580 19994 16632 20000
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16672 19916 16724 19922
rect 16672 19858 16724 19864
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15712 17632 15792 17660
rect 15660 17614 15712 17620
rect 15672 12714 15700 17614
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 14074 15792 14418
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15856 13530 15884 18158
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15948 15638 15976 16594
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 16040 12986 16068 17818
rect 16132 15162 16160 19246
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16316 17338 16344 18770
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 16114 16252 16594
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16224 15706 16252 16050
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16408 15586 16436 18702
rect 16592 18290 16620 19858
rect 16684 18834 16712 19858
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16960 19258 16988 22320
rect 17420 20058 17448 22320
rect 17408 20052 17460 20058
rect 17408 19994 17460 20000
rect 16868 18902 16896 19246
rect 16960 19230 17172 19258
rect 17144 19174 17172 19230
rect 17880 19174 17908 22320
rect 18340 20058 18368 22320
rect 18800 20074 18828 22320
rect 18328 20052 18380 20058
rect 18800 20046 18920 20074
rect 18328 19994 18380 20000
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 16672 18828 16724 18834
rect 16672 18770 16724 18776
rect 17776 18352 17828 18358
rect 17776 18294 17828 18300
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 17132 17808 17184 17814
rect 17132 17750 17184 17756
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 16726 16528 17614
rect 17144 17202 17172 17750
rect 17788 17746 17816 18294
rect 17972 18290 18000 19246
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18156 18902 18184 19178
rect 18616 18970 18644 19246
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18800 18902 18828 19858
rect 18892 19242 18920 20046
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 19260 19174 19288 22320
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 18144 18896 18196 18902
rect 18144 18838 18196 18844
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16960 16250 16988 16934
rect 17144 16794 17172 17138
rect 17132 16788 17184 16794
rect 17132 16730 17184 16736
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16316 15558 16436 15586
rect 16488 15564 16540 15570
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15764 11558 15792 12310
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15764 11218 15792 11494
rect 15948 11234 15976 12242
rect 16040 11354 16068 12922
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15752 11212 15804 11218
rect 15948 11206 16068 11234
rect 15752 11154 15804 11160
rect 15672 11014 15700 11154
rect 16040 11014 16068 11206
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15108 10542 15160 10548
rect 15304 10526 15424 10554
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15304 8838 15332 10526
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15396 9926 15424 10406
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15672 9518 15700 10610
rect 16040 10062 16068 10950
rect 16316 10810 16344 15558
rect 16488 15506 16540 15512
rect 16500 15026 16528 15506
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16500 14618 16528 14962
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16408 13326 16436 13738
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12986 16436 13262
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9722 16068 9998
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 16592 610 16620 13398
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12986 16988 13194
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16684 12442 16712 12786
rect 17420 12782 17448 14214
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17696 13394 17724 13806
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 17144 12306 17172 12650
rect 17788 12374 17816 17682
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17880 16538 17908 16594
rect 17880 16510 18000 16538
rect 17972 15502 18000 16510
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 15042 18000 15438
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17972 15014 18092 15042
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17972 13802 18000 14486
rect 18064 14482 18092 15014
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18248 14260 18276 14758
rect 18432 14618 18460 14758
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18524 14362 18552 18634
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17202 18644 17478
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18616 16726 18644 17138
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18524 14334 18644 14362
rect 18248 14232 18552 14260
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18524 13938 18552 14232
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18616 12986 18644 14334
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 13938 18736 14214
rect 18800 14074 18828 18702
rect 19720 18306 19748 22320
rect 19352 18278 19748 18306
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 19076 17338 19104 18158
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18708 13462 18736 13874
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17788 11558 17816 12310
rect 17972 11898 18000 12650
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18524 12442 18552 12582
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18524 11762 18552 12174
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 16684 11354 16712 11494
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 17972 11286 18000 11698
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 18616 11218 18644 11630
rect 18708 11354 18736 12786
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18892 11529 18920 11562
rect 18878 11520 18934 11529
rect 18878 11455 18934 11464
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 9586 16712 10406
rect 16868 10198 16896 10610
rect 18616 10538 18644 11154
rect 18708 10606 18736 11290
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16868 9722 16896 10134
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 18984 9110 19012 17070
rect 19168 16454 19196 17070
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19168 15638 19196 16390
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19076 12238 19104 13126
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 19352 8090 19380 18278
rect 20180 18154 20208 22320
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15026 19472 15302
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19444 14550 19472 14962
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 19536 7546 19564 18090
rect 20640 18086 20668 22320
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 19720 6390 19748 6802
rect 19904 6730 19932 18022
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 20824 5370 20852 18090
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20916 6458 20944 18022
rect 21100 16130 21128 22320
rect 21560 18086 21588 22320
rect 22020 18154 22048 22320
rect 22480 18358 22508 22320
rect 22468 18352 22520 18358
rect 22468 18294 22520 18300
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21008 16102 21128 16130
rect 21008 6730 21036 16102
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 16580 604 16632 610
rect 16580 546 16632 552
rect 17132 604 17184 610
rect 17132 546 17184 552
rect 17144 480 17172 546
rect 3330 232 3386 241
rect 3330 167 3386 176
rect 5722 0 5778 480
rect 17130 0 17186 480
<< via2 >>
rect 1398 22480 1454 22536
rect 1674 20576 1730 20632
rect 1950 18264 2006 18320
rect 2226 19216 2282 19272
rect 2042 18128 2098 18184
rect 1582 17312 1638 17368
rect 1674 16940 1676 16960
rect 1676 16940 1728 16960
rect 1728 16940 1730 16960
rect 1674 16904 1730 16940
rect 1582 16496 1638 16552
rect 1950 15952 2006 16008
rect 1674 14592 1730 14648
rect 1582 13640 1638 13696
rect 1950 14048 2006 14104
rect 2870 21528 2926 21584
rect 2778 21120 2834 21176
rect 2778 19760 2834 19816
rect 3238 22072 3294 22128
rect 3054 20168 3110 20224
rect 2410 19236 2466 19272
rect 2410 19216 2412 19236
rect 2412 19216 2464 19236
rect 2464 19216 2466 19236
rect 2686 18708 2688 18728
rect 2688 18708 2740 18728
rect 2740 18708 2742 18728
rect 2686 18672 2742 18708
rect 2318 18264 2374 18320
rect 2962 18808 3018 18864
rect 2778 17876 2834 17912
rect 2778 17856 2780 17876
rect 2780 17856 2832 17876
rect 2832 17856 2834 17876
rect 2778 15544 2834 15600
rect 3422 18808 3478 18864
rect 3606 18128 3662 18184
rect 3146 15000 3202 15056
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 5170 18264 5226 18320
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3238 8064 3294 8120
rect 4066 12688 4122 12744
rect 4066 12316 4068 12336
rect 4068 12316 4120 12336
rect 4120 12316 4122 12336
rect 4066 12280 4122 12316
rect 3974 10784 4030 10840
rect 3698 8472 3754 8528
rect 3054 3848 3110 3904
rect 3974 9424 4030 9480
rect 4066 9052 4068 9072
rect 4068 9052 4120 9072
rect 4120 9052 4122 9072
rect 4066 9016 4122 9052
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4250 8880 4306 8936
rect 3882 7520 3938 7576
rect 3882 5752 3938 5808
rect 3698 4256 3754 4312
rect 3146 3440 3202 3496
rect 2870 2896 2926 2952
rect 3790 1944 3846 2000
rect 3882 992 3938 1048
rect 4066 6160 4122 6216
rect 4066 4800 4122 4856
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4158 2488 4214 2544
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4710 5208 4766 5264
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4250 1536 4306 1592
rect 3974 584 4030 640
rect 7470 18808 7526 18864
rect 6458 13232 6514 13288
rect 6734 11328 6790 11384
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 9586 19236 9642 19272
rect 9586 19216 9588 19236
rect 9588 19216 9640 19236
rect 9640 19216 9642 19236
rect 9126 18708 9128 18728
rect 9128 18708 9180 18728
rect 9180 18708 9182 18728
rect 9126 18672 9182 18708
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7930 11736 7986 11792
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7654 7112 7710 7168
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7746 6704 7802 6760
rect 9218 9968 9274 10024
rect 8942 9696 8998 9752
rect 9310 9560 9366 9616
rect 9770 12552 9826 12608
rect 9494 10512 9550 10568
rect 8850 8916 8852 8936
rect 8852 8916 8904 8936
rect 8904 8916 8906 8936
rect 8850 8880 8906 8916
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 10598 12860 10600 12880
rect 10600 12860 10652 12880
rect 10652 12860 10654 12880
rect 10598 12824 10654 12860
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11242 11076 11298 11112
rect 11242 11056 11244 11076
rect 11244 11056 11296 11076
rect 11296 11056 11298 11076
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11978 18672 12034 18728
rect 11978 12844 12034 12880
rect 11978 12824 11980 12844
rect 11980 12824 12032 12844
rect 12032 12824 12034 12844
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 12714 11092 12716 11112
rect 12716 11092 12768 11112
rect 12768 11092 12770 11112
rect 12714 11056 12770 11092
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14370 18672 14426 18728
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14370 12552 14426 12608
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18878 11464 18934 11520
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 3330 176 3386 232
<< metal3 >>
rect 0 22538 480 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 480 22478
rect 1393 22475 1459 22478
rect 0 22130 480 22160
rect 3233 22130 3299 22133
rect 0 22128 3299 22130
rect 0 22072 3238 22128
rect 3294 22072 3299 22128
rect 0 22070 3299 22072
rect 0 22040 480 22070
rect 3233 22067 3299 22070
rect 0 21586 480 21616
rect 2865 21586 2931 21589
rect 0 21584 2931 21586
rect 0 21528 2870 21584
rect 2926 21528 2931 21584
rect 0 21526 2931 21528
rect 0 21496 480 21526
rect 2865 21523 2931 21526
rect 0 21178 480 21208
rect 2773 21178 2839 21181
rect 0 21176 2839 21178
rect 0 21120 2778 21176
rect 2834 21120 2839 21176
rect 0 21118 2839 21120
rect 0 21088 480 21118
rect 2773 21115 2839 21118
rect 0 20634 480 20664
rect 1669 20634 1735 20637
rect 0 20632 1735 20634
rect 0 20576 1674 20632
rect 1730 20576 1735 20632
rect 0 20574 1735 20576
rect 0 20544 480 20574
rect 1669 20571 1735 20574
rect 0 20226 480 20256
rect 3049 20226 3115 20229
rect 0 20224 3115 20226
rect 0 20168 3054 20224
rect 3110 20168 3115 20224
rect 0 20166 3115 20168
rect 0 20136 480 20166
rect 3049 20163 3115 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 2773 19818 2839 19821
rect 0 19816 2839 19818
rect 0 19760 2778 19816
rect 2834 19760 2839 19816
rect 0 19758 2839 19760
rect 0 19728 480 19758
rect 2773 19755 2839 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 2221 19274 2287 19277
rect 0 19272 2287 19274
rect 0 19216 2226 19272
rect 2282 19216 2287 19272
rect 0 19214 2287 19216
rect 0 19184 480 19214
rect 2221 19211 2287 19214
rect 2405 19274 2471 19277
rect 9581 19274 9647 19277
rect 2405 19272 9647 19274
rect 2405 19216 2410 19272
rect 2466 19216 9586 19272
rect 9642 19216 9647 19272
rect 2405 19214 9647 19216
rect 2405 19211 2471 19214
rect 9581 19211 9647 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 2957 18866 3023 18869
rect 0 18864 3023 18866
rect 0 18808 2962 18864
rect 3018 18808 3023 18864
rect 0 18806 3023 18808
rect 0 18776 480 18806
rect 2957 18803 3023 18806
rect 3417 18866 3483 18869
rect 7465 18866 7531 18869
rect 3417 18864 7531 18866
rect 3417 18808 3422 18864
rect 3478 18808 7470 18864
rect 7526 18808 7531 18864
rect 3417 18806 7531 18808
rect 3417 18803 3483 18806
rect 7465 18803 7531 18806
rect 2681 18730 2747 18733
rect 9121 18730 9187 18733
rect 2681 18728 9187 18730
rect 2681 18672 2686 18728
rect 2742 18672 9126 18728
rect 9182 18672 9187 18728
rect 2681 18670 9187 18672
rect 2681 18667 2747 18670
rect 9121 18667 9187 18670
rect 11973 18730 12039 18733
rect 14365 18730 14431 18733
rect 11973 18728 14431 18730
rect 11973 18672 11978 18728
rect 12034 18672 14370 18728
rect 14426 18672 14431 18728
rect 11973 18670 14431 18672
rect 11973 18667 12039 18670
rect 14365 18667 14431 18670
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 480 18262
rect 1945 18259 2011 18262
rect 2313 18322 2379 18325
rect 5165 18322 5231 18325
rect 2313 18320 5231 18322
rect 2313 18264 2318 18320
rect 2374 18264 5170 18320
rect 5226 18264 5231 18320
rect 2313 18262 5231 18264
rect 2313 18259 2379 18262
rect 5165 18259 5231 18262
rect 2037 18186 2103 18189
rect 3601 18186 3667 18189
rect 2037 18184 3667 18186
rect 2037 18128 2042 18184
rect 2098 18128 3606 18184
rect 3662 18128 3667 18184
rect 2037 18126 3667 18128
rect 2037 18123 2103 18126
rect 3601 18123 3667 18126
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 2773 17914 2839 17917
rect 0 17912 2839 17914
rect 0 17856 2778 17912
rect 2834 17856 2839 17912
rect 0 17854 2839 17856
rect 0 17824 480 17854
rect 2773 17851 2839 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 480 17310
rect 1577 17307 1643 17310
rect 0 16962 480 16992
rect 1669 16962 1735 16965
rect 0 16960 1735 16962
rect 0 16904 1674 16960
rect 1730 16904 1735 16960
rect 0 16902 1735 16904
rect 0 16872 480 16902
rect 1669 16899 1735 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 1577 16554 1643 16557
rect 0 16552 1643 16554
rect 0 16496 1582 16552
rect 1638 16496 1643 16552
rect 0 16494 1643 16496
rect 0 16464 480 16494
rect 1577 16491 1643 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 480 15950
rect 1945 15947 2011 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 2773 15602 2839 15605
rect 0 15600 2839 15602
rect 0 15544 2778 15600
rect 2834 15544 2839 15600
rect 0 15542 2839 15544
rect 0 15512 480 15542
rect 2773 15539 2839 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 3141 15058 3207 15061
rect 0 15056 3207 15058
rect 0 15000 3146 15056
rect 3202 15000 3207 15056
rect 0 14998 3207 15000
rect 0 14968 480 14998
rect 3141 14995 3207 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1945 14106 2011 14109
rect 0 14104 2011 14106
rect 0 14048 1950 14104
rect 2006 14048 2011 14104
rect 0 14046 2011 14048
rect 0 14016 480 14046
rect 1945 14043 2011 14046
rect 0 13698 480 13728
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13608 480 13638
rect 1577 13635 1643 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 6453 13290 6519 13293
rect 0 13288 6519 13290
rect 0 13232 6458 13288
rect 6514 13232 6519 13288
rect 0 13230 6519 13232
rect 0 13200 480 13230
rect 6453 13227 6519 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 10593 12882 10659 12885
rect 11973 12882 12039 12885
rect 10593 12880 12039 12882
rect 10593 12824 10598 12880
rect 10654 12824 11978 12880
rect 12034 12824 12039 12880
rect 10593 12822 12039 12824
rect 10593 12819 10659 12822
rect 11973 12819 12039 12822
rect 0 12746 480 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 9765 12610 9831 12613
rect 14365 12610 14431 12613
rect 9765 12608 14431 12610
rect 9765 12552 9770 12608
rect 9826 12552 14370 12608
rect 14426 12552 14431 12608
rect 9765 12550 14431 12552
rect 9765 12547 9831 12550
rect 14365 12547 14431 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 7925 11794 7991 11797
rect 0 11792 7991 11794
rect 0 11736 7930 11792
rect 7986 11736 7991 11792
rect 0 11734 7991 11736
rect 0 11704 480 11734
rect 7925 11731 7991 11734
rect 18873 11522 18939 11525
rect 22320 11522 22800 11552
rect 18873 11520 22800 11522
rect 18873 11464 18878 11520
rect 18934 11464 22800 11520
rect 18873 11462 22800 11464
rect 18873 11459 18939 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 22320 11432 22800 11462
rect 14672 11391 14992 11392
rect 6729 11386 6795 11389
rect 0 11384 6795 11386
rect 0 11328 6734 11384
rect 6790 11328 6795 11384
rect 0 11326 6795 11328
rect 0 11296 480 11326
rect 6729 11323 6795 11326
rect 11237 11114 11303 11117
rect 12709 11114 12775 11117
rect 11237 11112 12775 11114
rect 11237 11056 11242 11112
rect 11298 11056 12714 11112
rect 12770 11056 12775 11112
rect 11237 11054 12775 11056
rect 11237 11051 11303 11054
rect 12709 11051 12775 11054
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3969 10842 4035 10845
rect 0 10840 4035 10842
rect 0 10784 3974 10840
rect 4030 10784 4035 10840
rect 0 10782 4035 10784
rect 0 10752 480 10782
rect 3969 10779 4035 10782
rect 9489 10570 9555 10573
rect 4846 10568 9555 10570
rect 4846 10512 9494 10568
rect 9550 10512 9555 10568
rect 4846 10510 9555 10512
rect 0 10434 480 10464
rect 4846 10434 4906 10510
rect 9489 10507 9555 10510
rect 0 10374 4906 10434
rect 0 10344 480 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10026 480 10056
rect 9213 10026 9279 10029
rect 0 10024 9279 10026
rect 0 9968 9218 10024
rect 9274 9968 9279 10024
rect 0 9966 9279 9968
rect 0 9936 480 9966
rect 9213 9963 9279 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 8937 9754 9003 9757
rect 8937 9752 9506 9754
rect 8937 9696 8942 9752
rect 8998 9696 9506 9752
rect 8937 9694 9506 9696
rect 8937 9691 9003 9694
rect 9305 9618 9371 9621
rect 9446 9618 9506 9694
rect 9305 9616 9506 9618
rect 9305 9560 9310 9616
rect 9366 9560 9506 9616
rect 9305 9558 9506 9560
rect 9305 9555 9371 9558
rect 0 9482 480 9512
rect 3969 9482 4035 9485
rect 0 9480 4035 9482
rect 0 9424 3974 9480
rect 4030 9424 4035 9480
rect 0 9422 4035 9424
rect 0 9392 480 9422
rect 3969 9419 4035 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 480 9014
rect 4061 9011 4127 9014
rect 4245 8938 4311 8941
rect 8845 8938 8911 8941
rect 4245 8936 8911 8938
rect 4245 8880 4250 8936
rect 4306 8880 8850 8936
rect 8906 8880 8911 8936
rect 4245 8878 8911 8880
rect 4245 8875 4311 8878
rect 8845 8875 8911 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 3693 8530 3759 8533
rect 0 8528 3759 8530
rect 0 8472 3698 8528
rect 3754 8472 3759 8528
rect 0 8470 3759 8472
rect 0 8440 480 8470
rect 3693 8467 3759 8470
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 3233 8122 3299 8125
rect 0 8120 3299 8122
rect 0 8064 3238 8120
rect 3294 8064 3299 8120
rect 0 8062 3299 8064
rect 0 8032 480 8062
rect 3233 8059 3299 8062
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3877 7578 3943 7581
rect 0 7576 3943 7578
rect 0 7520 3882 7576
rect 3938 7520 3943 7576
rect 0 7518 3943 7520
rect 0 7488 480 7518
rect 3877 7515 3943 7518
rect 0 7170 480 7200
rect 7649 7170 7715 7173
rect 0 7168 7715 7170
rect 0 7112 7654 7168
rect 7710 7112 7715 7168
rect 0 7110 7715 7112
rect 0 7080 480 7110
rect 7649 7107 7715 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 7741 6762 7807 6765
rect 0 6760 7807 6762
rect 0 6704 7746 6760
rect 7802 6704 7807 6760
rect 0 6702 7807 6704
rect 0 6672 480 6702
rect 7741 6699 7807 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 3877 5810 3943 5813
rect 0 5808 3943 5810
rect 0 5752 3882 5808
rect 3938 5752 3943 5808
rect 0 5750 3943 5752
rect 0 5720 480 5750
rect 3877 5747 3943 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 4705 5266 4771 5269
rect 0 5264 4771 5266
rect 0 5208 4710 5264
rect 4766 5208 4771 5264
rect 0 5206 4771 5208
rect 0 5176 480 5206
rect 4705 5203 4771 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 480 4798
rect 4061 4795 4127 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 3693 4314 3759 4317
rect 0 4312 3759 4314
rect 0 4256 3698 4312
rect 3754 4256 3759 4312
rect 0 4254 3759 4256
rect 0 4224 480 4254
rect 3693 4251 3759 4254
rect 0 3906 480 3936
rect 3049 3906 3115 3909
rect 0 3904 3115 3906
rect 0 3848 3054 3904
rect 3110 3848 3115 3904
rect 0 3846 3115 3848
rect 0 3816 480 3846
rect 3049 3843 3115 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 3141 3498 3207 3501
rect 0 3496 3207 3498
rect 0 3440 3146 3496
rect 3202 3440 3207 3496
rect 0 3438 3207 3440
rect 0 3408 480 3438
rect 3141 3435 3207 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 2865 2954 2931 2957
rect 0 2952 2931 2954
rect 0 2896 2870 2952
rect 2926 2896 2931 2952
rect 0 2894 2931 2896
rect 0 2864 480 2894
rect 2865 2891 2931 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 4153 2546 4219 2549
rect 0 2544 4219 2546
rect 0 2488 4158 2544
rect 4214 2488 4219 2544
rect 0 2486 4219 2488
rect 0 2456 480 2486
rect 4153 2483 4219 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 3785 2002 3851 2005
rect 0 2000 3851 2002
rect 0 1944 3790 2000
rect 3846 1944 3851 2000
rect 0 1942 3851 1944
rect 0 1912 480 1942
rect 3785 1939 3851 1942
rect 0 1594 480 1624
rect 4245 1594 4311 1597
rect 0 1592 4311 1594
rect 0 1536 4250 1592
rect 4306 1536 4311 1592
rect 0 1534 4311 1536
rect 0 1504 480 1534
rect 4245 1531 4311 1534
rect 0 1050 480 1080
rect 3877 1050 3943 1053
rect 0 1048 3943 1050
rect 0 992 3882 1048
rect 3938 992 3943 1048
rect 0 990 3943 992
rect 0 960 480 990
rect 3877 987 3943 990
rect 0 642 480 672
rect 3969 642 4035 645
rect 0 640 4035 642
rect 0 584 3974 640
rect 4030 584 4035 640
rect 0 582 4035 584
rect 0 552 480 582
rect 3969 579 4035 582
rect 0 234 480 264
rect 3325 234 3391 237
rect 0 232 3391 234
rect 0 176 3330 232
rect 3386 176 3391 232
rect 0 174 3391 176
rect 0 144 480 174
rect 3325 171 3391 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1605641404
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1605641404
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1605641404
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1605641404
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1605641404
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1605641404
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1605641404
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1605641404
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1605641404
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1605641404
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1605641404
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1605641404
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1605641404
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1605641404
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1605641404
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1605641404
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1605641404
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1605641404
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1605641404
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1605641404
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1605641404
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1605641404
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1605641404
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1605641404
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1605641404
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1605641404
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1605641404
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1605641404
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1605641404
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1605641404
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1605641404
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1605641404
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1605641404
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1605641404
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1605641404
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1605641404
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1605641404
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1605641404
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1605641404
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1605641404
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1605641404
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1605641404
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1605641404
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1605641404
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1605641404
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1605641404
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1605641404
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1605641404
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1605641404
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1605641404
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1605641404
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1605641404
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp 1605641404
transform 1 0 20240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1605641404
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1605641404
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1605641404
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 7084 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1605641404
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1605641404
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1605641404
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1605641404
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1605641404
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1605641404
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1605641404
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1605641404
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1605641404
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1605641404
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1605641404
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1605641404
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1605641404
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1605641404
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1605641404
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1605641404
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1605641404
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1605641404
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1605641404
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp 1605641404
transform 1 0 20240 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 20516 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1605641404
transform 1 0 20884 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1605641404
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1840 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1605641404
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_14
timestamp 1605641404
transform 1 0 2392 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _066_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1605641404
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_35
timestamp 1605641404
transform 1 0 4324 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5612 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_47
timestamp 1605641404
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1605641404
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_76
timestamp 1605641404
transform 1 0 8096 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1605641404
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1605641404
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1605641404
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1605641404
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1605641404
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1605641404
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1605641404
transform 1 0 20240 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 19688 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1605641404
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1605641404
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1605641404
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2852 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1840 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1605641404
transform 1 0 1748 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 1605641404
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4508 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1605641404
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1605641404
transform 1 0 5980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8004 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6992 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1605641404
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_84
timestamp 1605641404
transform 1 0 8832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1605641404
transform 1 0 9936 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_108
timestamp 1605641404
transform 1 0 11040 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1605641404
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1605641404
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1605641404
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1605641404
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1605641404
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 19320 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1605641404
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_202
timestamp 1605641404
transform 1 0 19688 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_214
timestamp 1605641404
transform 1 0 20792 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1840 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1605641404
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_24
timestamp 1605641404
transform 1 0 3312 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1605641404
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6532 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5060 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_52
timestamp 1605641404
transform 1 0 5888 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_58
timestamp 1605641404
transform 1 0 6440 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8372 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_75
timestamp 1605641404
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1605641404
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1605641404
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1605641404
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1605641404
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1605641404
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1605641404
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1605641404
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1605641404
transform 1 0 18860 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_190
timestamp 1605641404
transform 1 0 18584 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1605641404
transform 1 0 19228 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1605641404
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1605641404
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1605641404
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1748 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 3772 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_11_23
timestamp 1605641404
transform 1 0 3220 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1605641404
transform 1 0 4600 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 5428 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_46
timestamp 1605641404
transform 1 0 5336 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1605641404
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7820 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_89
timestamp 1605641404
transform 1 0 9292 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_101
timestamp 1605641404
transform 1 0 10396 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1605641404
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1605641404
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1605641404
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1605641404
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1605641404
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1605641404
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1605641404
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1605641404
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2484 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1605641404
transform 1 0 2116 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_24
timestamp 1605641404
transform 1 0 3312 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1605641404
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6072 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_44
timestamp 1605641404
transform 1 0 5152 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1605641404
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8372 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1605641404
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_76
timestamp 1605641404
transform 1 0 8096 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1605641404
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1605641404
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1605641404
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1605641404
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1605641404
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1605641404
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1605641404
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1605641404
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1605641404
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1564 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 2484 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1605641404
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 3496 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1605641404
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_35
timestamp 1605641404
transform 1 0 4324 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_21
timestamp 1605641404
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1605641404
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1605641404
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6348 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_48
timestamp 1605641404
transform 1 0 5520 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1605641404
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8556 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_71
timestamp 1605641404
transform 1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_79
timestamp 1605641404
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1605641404
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10212 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 1605641404
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1605641404
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11040 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_108
timestamp 1605641404
transform 1 0 11040 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1605641404
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1605641404
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_124
timestamp 1605641404
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12696 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_132
timestamp 1605641404
transform 1 0 13248 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_144
timestamp 1605641404
transform 1 0 14352 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_142
timestamp 1605641404
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16008 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15364 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_152
timestamp 1605641404
transform 1 0 15088 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1605641404
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 17020 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1605641404
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1605641404
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1605641404
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1605641404
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1605641404
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1605641404
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1605641404
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1605641404
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1748 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1605641404
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3496 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1605641404
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_35
timestamp 1605641404
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1605641404
transform 1 0 5244 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 1605641404
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1605641404
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1605641404
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 8464 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7452 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1605641404
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1605641404
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1605641404
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10028 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 8924 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_88
timestamp 1605641404
transform 1 0 9200 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_96
timestamp 1605641404
transform 1 0 9936 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 12604 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1605641404
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1605641404
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 12880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13340 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1605641404
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16284 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1605641404
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_160
timestamp 1605641404
transform 1 0 15824 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_164
timestamp 1605641404
transform 1 0 16192 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_174
timestamp 1605641404
transform 1 0 17112 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1605641404
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_200
timestamp 1605641404
transform 1 0 19504 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1605641404
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_9
timestamp 1605641404
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_19
timestamp 1605641404
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4508 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1605641404
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5520 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1605641404
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_57
timestamp 1605641404
transform 1 0 6348 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_61
timestamp 1605641404
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1605641404
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_82
timestamp 1605641404
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1605641404
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1605641404
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 1605641404
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_119
timestamp 1605641404
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 1605641404
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1605641404
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1605641404
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17296 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1605641404
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_192
timestamp 1605641404
transform 1 0 18768 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1605641404
transform 1 0 19872 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1605641404
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1605641404
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 2668 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1932 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1605641404
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1605641404
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3772 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_21
timestamp 1605641404
transform 1 0 3036 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1605641404
transform 1 0 5244 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_49
timestamp 1605641404
transform 1 0 5612 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 6992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_67
timestamp 1605641404
transform 1 0 7268 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9752 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1605641404
transform 1 0 8832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1605641404
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1605641404
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1605641404
transform 1 0 13432 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14352 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1605641404
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_137
timestamp 1605641404
transform 1 0 13708 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_143
timestamp 1605641404
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1605641404
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_165
timestamp 1605641404
transform 1 0 16284 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_171
timestamp 1605641404
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1605641404
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_187
timestamp 1605641404
transform 1 0 18308 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18584 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_206
timestamp 1605641404
transform 1 0 20056 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1605641404
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2760 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1605641404
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1605641404
transform 1 0 2576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 3496 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4232 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_24
timestamp 1605641404
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5888 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_50
timestamp 1605641404
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7728 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1605641404
transform 1 0 7360 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1605641404
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_102
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11960 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_114
timestamp 1605641404
transform 1 0 11592 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1605641404
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_145
timestamp 1605641404
transform 1 0 14444 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_149
timestamp 1605641404
transform 1 0 14812 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 17572 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_170
timestamp 1605641404
transform 1 0 16744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_178
timestamp 1605641404
transform 1 0 17480 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_188
timestamp 1605641404
transform 1 0 18400 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_200
timestamp 1605641404
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1605641404
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1605641404
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1932 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1605641404
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_17
timestamp 1605641404
transform 1 0 2668 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1605641404
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2668 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 2300 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3220 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1605641404
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_26
timestamp 1605641404
transform 1 0 3496 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1605641404
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_41
timestamp 1605641404
transform 1 0 4876 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1605641404
transform 1 0 6164 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6256 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5244 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1605641404
transform 1 0 5796 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1605641404
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1605641404
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_73
timestamp 1605641404
transform 1 0 7820 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_72
timestamp 1605641404
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9200 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10672 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10120 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_19_85
timestamp 1605641404
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1605641404
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_96
timestamp 1605641404
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12512 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11500 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_118
timestamp 1605641404
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 14444 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1605641404
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1605641404
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1605641404
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15732 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_148
timestamp 1605641404
transform 1 0 14720 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1605641404
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1605641404
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_173
timestamp 1605641404
transform 1 0 17020 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1605641404
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1605641404
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1605641404
transform 1 0 16744 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1605641404
transform 1 0 17572 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1605641404
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17664 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1605641404
transform 1 0 18860 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1605641404
transform 1 0 19964 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1605641404
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1605641404
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1605641404
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2392 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1605641404
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4508 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_21_30
timestamp 1605641404
transform 1 0 3864 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_36
timestamp 1605641404
transform 1 0 4416 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5520 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 1605641404
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1605641404
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7912 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_71
timestamp 1605641404
transform 1 0 7636 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10212 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_90
timestamp 1605641404
transform 1 0 9384 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_98
timestamp 1605641404
transform 1 0 10120 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12604 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10948 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1605641404
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_116
timestamp 1605641404
transform 1 0 11776 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_134
timestamp 1605641404
transform 1 0 13432 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16008 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1605641404
transform 1 0 14536 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_150
timestamp 1605641404
transform 1 0 14904 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1605641404
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_178
timestamp 1605641404
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1605641404
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1605641404
transform 1 0 18860 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1605641404
transform 1 0 19964 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1605641404
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1932 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1605641404
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1605641404
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4324 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1605641404
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6256 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1605641404
transform 1 0 5796 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_55
timestamp 1605641404
transform 1 0 6164 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1605641404
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_72
timestamp 1605641404
transform 1 0 7728 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1605641404
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10488 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 1605641404
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12328 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1605641404
transform 1 0 11960 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13064 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1605641404
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15456 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_146
timestamp 1605641404
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1605641404
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 17480 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17940 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_172
timestamp 1605641404
transform 1 0 16928 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_181
timestamp 1605641404
transform 1 0 17756 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_199
timestamp 1605641404
transform 1 0 19412 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_211
timestamp 1605641404
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1605641404
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1840 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2576 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1605641404
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1605641404
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4692 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_25
timestamp 1605641404
transform 1 0 3404 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_37
timestamp 1605641404
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_55
timestamp 1605641404
transform 1 0 6164 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8464 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 6992 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_67
timestamp 1605641404
transform 1 0 7268 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1605641404
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_96
timestamp 1605641404
transform 1 0 9936 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_104
timestamp 1605641404
transform 1 0 10672 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1605641404
transform 1 0 10948 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1605641404
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13708 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_126
timestamp 1605641404
transform 1 0 12696 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_133
timestamp 1605641404
transform 1 0 13340 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15916 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_146
timestamp 1605641404
transform 1 0 14536 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_158
timestamp 1605641404
transform 1 0 15640 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 16928 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_170
timestamp 1605641404
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1605641404
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_195
timestamp 1605641404
transform 1 0 19044 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_207
timestamp 1605641404
transform 1 0 20148 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1605641404
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2300 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1605641404
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1605641404
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1605641404
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_35
timestamp 1605641404
transform 1 0 4324 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6532 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 5336 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_44
timestamp 1605641404
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_49
timestamp 1605641404
transform 1 0 5612 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1605641404
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1605641404
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_79
timestamp 1605641404
transform 1 0 8372 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1605641404
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1605641404
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12420 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1605641404
transform 1 0 11224 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1605641404
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13432 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp 1605641404
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15732 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1605641404
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1605641404
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18032 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_175
timestamp 1605641404
transform 1 0 17204 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_183
timestamp 1605641404
transform 1 0 17940 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_200
timestamp 1605641404
transform 1 0 19504 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1605641404
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 2668 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1932 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1605641404
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1605641404
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4600 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1605641404
transform 1 0 3404 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1605641404
transform 1 0 3036 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_34
timestamp 1605641404
transform 1 0 4232 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1605641404
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1605641404
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1605641404
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_78
timestamp 1605641404
transform 1 0 8280 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1605641404
transform 1 0 8924 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9384 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_84
timestamp 1605641404
transform 1 0 8832 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_88
timestamp 1605641404
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1605641404
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1605641404
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1605641404
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14076 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1605641404
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15548 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 15272 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_150
timestamp 1605641404
transform 1 0 14904 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_166
timestamp 1605641404
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1605641404
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1605641404
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1605641404
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1605641404
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_8
timestamp 1605641404
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1605641404
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 1472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1605641404
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1605641404
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_17
timestamp 1605641404
transform 1 0 2668 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2760 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4784 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4508 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1605641404
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1605641404
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_34
timestamp 1605641404
transform 1 0 4232 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1605641404
transform 1 0 6532 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5520 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_46
timestamp 1605641404
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1605641404
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp 1605641404
transform 1 0 6808 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1605641404
transform 1 0 6256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1605641404
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1605641404
transform 1 0 7912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7268 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8740 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 7636 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1605641404
transform 1 0 7176 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_83
timestamp 1605641404
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1605641404
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_77
timestamp 1605641404
transform 1 0 8188 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9752 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1605641404
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1605641404
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_89
timestamp 1605641404
transform 1 0 9292 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_95
timestamp 1605641404
transform 1 0 9844 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12512 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12328 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_110
timestamp 1605641404
transform 1 0 11224 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_105
timestamp 1605641404
transform 1 0 10764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1605641404
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14352 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_131
timestamp 1605641404
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_143
timestamp 1605641404
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_140
timestamp 1605641404
transform 1 0 13984 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1605641404
transform 1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15916 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1605641404
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_154
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_160
timestamp 1605641404
transform 1 0 15824 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_160
timestamp 1605641404
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1605641404
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17756 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16468 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_177
timestamp 1605641404
transform 1 0 17388 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_176
timestamp 1605641404
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1605641404
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19044 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1605641404
transform 1 0 19228 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1605641404
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_204
timestamp 1605641404
transform 1 0 19872 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1605641404
transform 1 0 20332 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1605641404
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_216
timestamp 1605641404
transform 1 0 20976 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 2300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1605641404
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1605641404
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 3404 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1605641404
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1605641404
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 6808 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5612 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_44
timestamp 1605641404
transform 1 0 5152 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_48
timestamp 1605641404
transform 1 0 5520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1605641404
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1605641404
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1605641404
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1605641404
transform 1 0 8740 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9936 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 8832 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1605641404
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1605641404
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_105
timestamp 1605641404
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1605641404
transform 1 0 11224 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_122
timestamp 1605641404
transform 1 0 12328 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_132
timestamp 1605641404
transform 1 0 13248 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_140
timestamp 1605641404
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1605641404
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1605641404
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16928 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_171
timestamp 1605641404
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_188
timestamp 1605641404
transform 1 0 18400 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_200
timestamp 1605641404
transform 1 0 19504 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1605641404
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2668 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1932 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1605641404
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1605641404
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_33
timestamp 1605641404
transform 1 0 4140 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1605641404
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1605641404
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_62
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10304 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1605641404
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_95
timestamp 1605641404
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_99
timestamp 1605641404
transform 1 0 10212 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_116
timestamp 1605641404
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1605641404
transform 1 0 14076 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1605641404
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1605641404
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 15640 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16284 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14628 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_156
timestamp 1605641404
transform 1 0 15456 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_161
timestamp 1605641404
transform 1 0 15916 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1605641404
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_190
timestamp 1605641404
transform 1 0 18584 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_202
timestamp 1605641404
transform 1 0 19688 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_214
timestamp 1605641404
transform 1 0 20792 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1605641404
transform 1 0 2760 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_9
timestamp 1605641404
transform 1 0 1932 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_16
timestamp 1605641404
transform 1 0 2576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1605641404
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1605641404
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1605641404
transform 1 0 6072 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5060 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1605641404
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_57
timestamp 1605641404
transform 1 0 6348 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8372 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 7636 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1605641404
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1605641404
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1605641404
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12512 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11776 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_109
timestamp 1605641404
transform 1 0 11132 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1605641404
transform 1 0 11684 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_122
timestamp 1605641404
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 13524 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_130
timestamp 1605641404
transform 1 0 13064 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_134
timestamp 1605641404
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 15456 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16284 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1605641404
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_162
timestamp 1605641404
transform 1 0 16008 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17756 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17020 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_171
timestamp 1605641404
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_179
timestamp 1605641404
transform 1 0 17572 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_187
timestamp 1605641404
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18492 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_195
timestamp 1605641404
transform 1 0 19044 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1605641404
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1605641404
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 1564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1605641404
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_17
timestamp 1605641404
transform 1 0 2668 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 3036 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_37
timestamp 1605641404
transform 1 0 4508 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5060 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1605641404
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1605641404
transform 1 0 8740 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_78
timestamp 1605641404
transform 1 0 8280 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_82
timestamp 1605641404
transform 1 0 8648 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9200 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1605641404
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1605641404
transform 1 0 10672 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 11500 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_112
timestamp 1605641404
transform 1 0 11408 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1605641404
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1605641404
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 12880 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13616 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_127
timestamp 1605641404
transform 1 0 12788 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_132
timestamp 1605641404
transform 1 0 13248 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1605641404
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16100 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14628 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_156
timestamp 1605641404
transform 1 0 15456 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_162
timestamp 1605641404
transform 1 0 16008 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 17388 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 16836 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1605641404
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1605641404
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1605641404
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 18584 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 19136 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1605641404
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1605641404
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_200
timestamp 1605641404
transform 1 0 19504 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_212
timestamp 1605641404
transform 1 0 20608 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1605641404
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1605641404
transform 1 0 2668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1605641404
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_25
timestamp 1605641404
transform 1 0 3404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1605641404
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_41
timestamp 1605641404
transform 1 0 4876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5336 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1605641404
transform 1 0 5244 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_55
timestamp 1605641404
transform 1 0 6164 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1605641404
transform 1 0 6716 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8648 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_75
timestamp 1605641404
transform 1 0 8004 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_81
timestamp 1605641404
transform 1 0 8556 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1605641404
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_94
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_102
timestamp 1605641404
transform 1 0 10488 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 10764 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_121
timestamp 1605641404
transform 1 0 12236 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 12972 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13800 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_133
timestamp 1605641404
transform 1 0 13340 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_137
timestamp 1605641404
transform 1 0 13708 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1605641404
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 14536 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_152
timestamp 1605641404
transform 1 0 15088 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1605641404
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_166
timestamp 1605641404
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 17112 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_172
timestamp 1605641404
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_178
timestamp 1605641404
transform 1 0 17480 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_191
timestamp 1605641404
transform 1 0 18676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_203
timestamp 1605641404
transform 1 0 19780 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1605641404
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal3 s 22320 11432 22800 11552 6 ccff_head
port 0 nsew default input
rlabel metal2 s 17130 0 17186 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 3882 22320 3938 22800 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 9034 22320 9090 22800 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9494 22320 9550 22800 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9954 22320 10010 22800 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10414 22320 10470 22800 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 10874 22320 10930 22800 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11334 22320 11390 22800 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 11794 22320 11850 22800 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 12254 22320 12310 22800 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 12714 22320 12770 22800 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 4342 22320 4398 22800 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 4802 22320 4858 22800 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 5722 22320 5778 22800 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 6182 22320 6238 22800 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 6642 22320 6698 22800 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 7102 22320 7158 22800 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 7562 22320 7618 22800 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 8114 22320 8170 22800 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 13174 22320 13230 22800 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17866 22320 17922 22800 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 18326 22320 18382 22800 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18786 22320 18842 22800 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 19246 22320 19302 22800 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19706 22320 19762 22800 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 20166 22320 20222 22800 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20626 22320 20682 22800 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 21086 22320 21142 22800 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21546 22320 21602 22800 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 22006 22320 22062 22800 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 14094 22320 14150 22800 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 14554 22320 14610 22800 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 15014 22320 15070 22800 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 15566 22320 15622 22800 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 16026 22320 16082 22800 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 16486 22320 16542 22800 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16946 22320 17002 22800 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 17406 22320 17462 22800 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_13_
port 83 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_15_
port 84 nsew default input
rlabel metal3 s 0 3816 480 3936 6 left_bottom_grid_pin_17_
port 85 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 86 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 87 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_5_
port 88 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_7_
port 89 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_9_
port 90 nsew default input
rlabel metal2 s 5722 0 5778 480 6 prog_clk
port 91 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 92 nsew default input
rlabel metal2 s 662 22320 718 22800 6 top_left_grid_pin_43_
port 93 nsew default input
rlabel metal2 s 1122 22320 1178 22800 6 top_left_grid_pin_44_
port 94 nsew default input
rlabel metal2 s 1582 22320 1638 22800 6 top_left_grid_pin_45_
port 95 nsew default input
rlabel metal2 s 2042 22320 2098 22800 6 top_left_grid_pin_46_
port 96 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 top_left_grid_pin_47_
port 97 nsew default input
rlabel metal2 s 2962 22320 3018 22800 6 top_left_grid_pin_48_
port 98 nsew default input
rlabel metal2 s 3422 22320 3478 22800 6 top_left_grid_pin_49_
port 99 nsew default input
rlabel metal2 s 22466 22320 22522 22800 6 top_right_grid_pin_1_
port 100 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 101 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 102 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
