VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 114.280 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.880 2.400 28.480 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.000 2.400 85.600 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 14.280 115.000 14.880 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 38.760 115.000 39.360 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 41.480 115.000 42.080 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 43.520 115.000 44.120 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 46.240 115.000 46.840 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 48.280 115.000 48.880 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 51.000 115.000 51.600 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 53.720 115.000 54.320 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 55.760 115.000 56.360 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 58.480 115.000 59.080 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 60.520 115.000 61.120 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 17.000 115.000 17.600 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 19.040 115.000 19.640 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 21.760 115.000 22.360 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 23.800 115.000 24.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 26.520 115.000 27.120 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 29.240 115.000 29.840 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 31.280 115.000 31.880 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 34.000 115.000 34.600 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 36.040 115.000 36.640 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 63.240 115.000 63.840 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 87.720 115.000 88.320 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 90.440 115.000 91.040 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 92.480 115.000 93.080 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 95.200 115.000 95.800 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 97.240 115.000 97.840 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 99.960 115.000 100.560 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 102.680 115.000 103.280 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 104.720 115.000 105.320 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 107.440 115.000 108.040 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 109.480 115.000 110.080 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 65.960 115.000 66.560 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 68.000 115.000 68.600 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 70.720 115.000 71.320 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 72.760 115.000 73.360 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 75.480 115.000 76.080 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 78.200 115.000 78.800 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 80.240 115.000 80.840 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 82.960 115.000 83.560 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 85.000 115.000 85.600 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 111.880 4.510 114.280 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 111.880 32.570 114.280 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 111.880 35.330 114.280 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 111.880 38.090 114.280 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 111.880 40.850 114.280 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 111.880 43.610 114.280 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 111.880 46.370 114.280 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 111.880 49.130 114.280 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.610 111.880 51.890 114.280 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 111.880 54.650 114.280 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 111.880 57.410 114.280 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 111.880 7.270 114.280 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 111.880 10.030 114.280 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 111.880 12.790 114.280 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 111.880 15.550 114.280 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 111.880 18.310 114.280 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 111.880 21.070 114.280 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 111.880 23.830 114.280 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 111.880 26.590 114.280 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 111.880 29.350 114.280 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.350 111.880 60.630 114.280 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 111.880 88.690 114.280 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 111.880 91.450 114.280 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 111.880 94.210 114.280 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 111.880 96.970 114.280 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 111.880 99.730 114.280 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 111.880 102.490 114.280 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 111.880 105.250 114.280 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 111.880 108.010 114.280 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 111.880 110.770 114.280 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.250 111.880 113.530 114.280 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 111.880 63.390 114.280 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 111.880 66.150 114.280 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 111.880 68.910 114.280 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 111.880 71.670 114.280 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 111.880 74.430 114.280 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 111.880 77.190 114.280 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 111.880 79.950 114.280 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 111.880 82.710 114.280 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 111.880 85.470 114.280 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 112.200 115.000 112.800 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 11.560 115.000 12.160 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 0.000 115.000 0.600 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 2.040 115.000 2.640 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 4.760 115.000 5.360 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 6.800 115.000 7.400 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 9.520 115.000 10.120 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 111.880 1.750 114.280 ;
    END
  END top_left_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.045 9.920 23.645 102.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.375 9.920 40.975 102.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.075 109.480 102.725 ;
      LAYER met1 ;
        RECT 1.450 5.780 113.550 102.880 ;
      LAYER met2 ;
        RECT 2.030 111.600 3.950 112.685 ;
        RECT 4.790 111.600 6.710 112.685 ;
        RECT 7.550 111.600 9.470 112.685 ;
        RECT 10.310 111.600 12.230 112.685 ;
        RECT 13.070 111.600 14.990 112.685 ;
        RECT 15.830 111.600 17.750 112.685 ;
        RECT 18.590 111.600 20.510 112.685 ;
        RECT 21.350 111.600 23.270 112.685 ;
        RECT 24.110 111.600 26.030 112.685 ;
        RECT 26.870 111.600 28.790 112.685 ;
        RECT 29.630 111.600 32.010 112.685 ;
        RECT 32.850 111.600 34.770 112.685 ;
        RECT 35.610 111.600 37.530 112.685 ;
        RECT 38.370 111.600 40.290 112.685 ;
        RECT 41.130 111.600 43.050 112.685 ;
        RECT 43.890 111.600 45.810 112.685 ;
        RECT 46.650 111.600 48.570 112.685 ;
        RECT 49.410 111.600 51.330 112.685 ;
        RECT 52.170 111.600 54.090 112.685 ;
        RECT 54.930 111.600 56.850 112.685 ;
        RECT 57.690 111.600 60.070 112.685 ;
        RECT 60.910 111.600 62.830 112.685 ;
        RECT 63.670 111.600 65.590 112.685 ;
        RECT 66.430 111.600 68.350 112.685 ;
        RECT 69.190 111.600 71.110 112.685 ;
        RECT 71.950 111.600 73.870 112.685 ;
        RECT 74.710 111.600 76.630 112.685 ;
        RECT 77.470 111.600 79.390 112.685 ;
        RECT 80.230 111.600 82.150 112.685 ;
        RECT 82.990 111.600 84.910 112.685 ;
        RECT 85.750 111.600 88.130 112.685 ;
        RECT 88.970 111.600 90.890 112.685 ;
        RECT 91.730 111.600 93.650 112.685 ;
        RECT 94.490 111.600 96.410 112.685 ;
        RECT 97.250 111.600 99.170 112.685 ;
        RECT 100.010 111.600 101.930 112.685 ;
        RECT 102.770 111.600 104.690 112.685 ;
        RECT 105.530 111.600 107.450 112.685 ;
        RECT 108.290 111.600 110.210 112.685 ;
        RECT 111.050 111.600 112.970 112.685 ;
        RECT 1.480 0.115 113.520 111.600 ;
      LAYER met3 ;
        RECT 2.400 111.800 112.200 112.665 ;
        RECT 2.400 110.480 112.600 111.800 ;
        RECT 2.400 109.080 112.200 110.480 ;
        RECT 2.400 108.440 112.600 109.080 ;
        RECT 2.400 107.040 112.200 108.440 ;
        RECT 2.400 105.720 112.600 107.040 ;
        RECT 2.400 104.320 112.200 105.720 ;
        RECT 2.400 103.680 112.600 104.320 ;
        RECT 2.400 102.280 112.200 103.680 ;
        RECT 2.400 100.960 112.600 102.280 ;
        RECT 2.400 99.560 112.200 100.960 ;
        RECT 2.400 98.240 112.600 99.560 ;
        RECT 2.400 96.840 112.200 98.240 ;
        RECT 2.400 96.200 112.600 96.840 ;
        RECT 2.400 94.800 112.200 96.200 ;
        RECT 2.400 93.480 112.600 94.800 ;
        RECT 2.400 92.080 112.200 93.480 ;
        RECT 2.400 91.440 112.600 92.080 ;
        RECT 2.400 90.040 112.200 91.440 ;
        RECT 2.400 88.720 112.600 90.040 ;
        RECT 2.400 87.320 112.200 88.720 ;
        RECT 2.400 86.000 112.600 87.320 ;
        RECT 2.800 84.600 112.200 86.000 ;
        RECT 2.400 83.960 112.600 84.600 ;
        RECT 2.400 82.560 112.200 83.960 ;
        RECT 2.400 81.240 112.600 82.560 ;
        RECT 2.400 79.840 112.200 81.240 ;
        RECT 2.400 79.200 112.600 79.840 ;
        RECT 2.400 77.800 112.200 79.200 ;
        RECT 2.400 76.480 112.600 77.800 ;
        RECT 2.400 75.080 112.200 76.480 ;
        RECT 2.400 73.760 112.600 75.080 ;
        RECT 2.400 72.360 112.200 73.760 ;
        RECT 2.400 71.720 112.600 72.360 ;
        RECT 2.400 70.320 112.200 71.720 ;
        RECT 2.400 69.000 112.600 70.320 ;
        RECT 2.400 67.600 112.200 69.000 ;
        RECT 2.400 66.960 112.600 67.600 ;
        RECT 2.400 65.560 112.200 66.960 ;
        RECT 2.400 64.240 112.600 65.560 ;
        RECT 2.400 62.840 112.200 64.240 ;
        RECT 2.400 61.520 112.600 62.840 ;
        RECT 2.400 60.120 112.200 61.520 ;
        RECT 2.400 59.480 112.600 60.120 ;
        RECT 2.400 58.080 112.200 59.480 ;
        RECT 2.400 56.760 112.600 58.080 ;
        RECT 2.400 55.360 112.200 56.760 ;
        RECT 2.400 54.720 112.600 55.360 ;
        RECT 2.400 53.320 112.200 54.720 ;
        RECT 2.400 52.000 112.600 53.320 ;
        RECT 2.400 50.600 112.200 52.000 ;
        RECT 2.400 49.280 112.600 50.600 ;
        RECT 2.400 47.880 112.200 49.280 ;
        RECT 2.400 47.240 112.600 47.880 ;
        RECT 2.400 45.840 112.200 47.240 ;
        RECT 2.400 44.520 112.600 45.840 ;
        RECT 2.400 43.120 112.200 44.520 ;
        RECT 2.400 42.480 112.600 43.120 ;
        RECT 2.400 41.080 112.200 42.480 ;
        RECT 2.400 39.760 112.600 41.080 ;
        RECT 2.400 38.360 112.200 39.760 ;
        RECT 2.400 37.040 112.600 38.360 ;
        RECT 2.400 35.640 112.200 37.040 ;
        RECT 2.400 35.000 112.600 35.640 ;
        RECT 2.400 33.600 112.200 35.000 ;
        RECT 2.400 32.280 112.600 33.600 ;
        RECT 2.400 30.880 112.200 32.280 ;
        RECT 2.400 30.240 112.600 30.880 ;
        RECT 2.400 28.880 112.200 30.240 ;
        RECT 2.800 28.840 112.200 28.880 ;
        RECT 2.800 27.520 112.600 28.840 ;
        RECT 2.800 27.480 112.200 27.520 ;
        RECT 2.400 26.120 112.200 27.480 ;
        RECT 2.400 24.800 112.600 26.120 ;
        RECT 2.400 23.400 112.200 24.800 ;
        RECT 2.400 22.760 112.600 23.400 ;
        RECT 2.400 21.360 112.200 22.760 ;
        RECT 2.400 20.040 112.600 21.360 ;
        RECT 2.400 18.640 112.200 20.040 ;
        RECT 2.400 18.000 112.600 18.640 ;
        RECT 2.400 16.600 112.200 18.000 ;
        RECT 2.400 15.280 112.600 16.600 ;
        RECT 2.400 13.880 112.200 15.280 ;
        RECT 2.400 12.560 112.600 13.880 ;
        RECT 2.400 11.160 112.200 12.560 ;
        RECT 2.400 10.520 112.600 11.160 ;
        RECT 2.400 9.120 112.200 10.520 ;
        RECT 2.400 7.800 112.600 9.120 ;
        RECT 2.400 6.400 112.200 7.800 ;
        RECT 2.400 5.760 112.600 6.400 ;
        RECT 2.400 4.360 112.200 5.760 ;
        RECT 2.400 3.040 112.600 4.360 ;
        RECT 2.400 1.640 112.200 3.040 ;
        RECT 2.400 1.000 112.600 1.640 ;
        RECT 2.400 0.135 112.200 1.000 ;
      LAYER met4 ;
        RECT 41.375 9.920 94.465 102.880 ;
  END
END sb_0__0_
END LIBRARY

