magic
tech EFS8A
magscale 1 2
timestamp 1602873394
<< locali >>
rect 22511 24225 22546 24259
rect 17601 23511 17635 23749
rect 12633 23137 12794 23171
rect 16071 23137 16106 23171
rect 22511 23137 22546 23171
rect 23523 23137 23650 23171
rect 12633 22967 12667 23137
rect 16215 21097 16221 21131
rect 16215 21029 16249 21097
rect 16583 20247 16617 20315
rect 16583 20213 16589 20247
rect 18831 17697 18866 17731
rect 20821 17051 20855 17289
rect 12627 15657 12633 15691
rect 12627 15589 12661 15657
rect 5503 14841 5641 14875
rect 22839 13481 22845 13515
rect 22839 13413 22873 13481
rect 21643 11305 21649 11339
rect 21643 11237 21677 11305
rect 17693 10455 17727 10761
rect 19349 8347 19383 8517
rect 12443 8041 12449 8075
rect 12443 7973 12477 8041
rect 14191 5015 14225 5083
rect 14191 4981 14197 5015
rect 18923 4641 18958 4675
rect 15243 3553 15370 3587
rect 24501 3553 24662 3587
rect 24501 3383 24535 3553
<< viali >>
rect 24777 25449 24811 25483
rect 24593 25313 24627 25347
rect 24777 24905 24811 24939
rect 18475 24837 18509 24871
rect 22707 24837 22741 24871
rect 18404 24701 18438 24735
rect 19476 24701 19510 24735
rect 19901 24701 19935 24735
rect 22636 24701 22670 24735
rect 24593 24701 24627 24735
rect 25145 24701 25179 24735
rect 18797 24633 18831 24667
rect 19579 24633 19613 24667
rect 16957 24565 16991 24599
rect 20453 24565 20487 24599
rect 23121 24565 23155 24599
rect 24409 24565 24443 24599
rect 15485 24361 15519 24395
rect 18337 24361 18371 24395
rect 24777 24361 24811 24395
rect 21097 24293 21131 24327
rect 1444 24225 1478 24259
rect 12976 24225 13010 24259
rect 15301 24225 15335 24259
rect 17208 24225 17242 24259
rect 18153 24225 18187 24259
rect 19292 24225 19326 24259
rect 22477 24225 22511 24259
rect 23648 24225 23682 24259
rect 24593 24225 24627 24259
rect 21005 24157 21039 24191
rect 21281 24157 21315 24191
rect 17279 24089 17313 24123
rect 18705 24089 18739 24123
rect 22615 24089 22649 24123
rect 1547 24021 1581 24055
rect 13047 24021 13081 24055
rect 19395 24021 19429 24055
rect 20453 24021 20487 24055
rect 23719 24021 23753 24055
rect 1869 23817 1903 23851
rect 11713 23817 11747 23851
rect 13001 23817 13035 23851
rect 13369 23817 13403 23851
rect 15577 23817 15611 23851
rect 17417 23817 17451 23851
rect 19257 23817 19291 23851
rect 21373 23817 21407 23851
rect 22201 23817 22235 23851
rect 23857 23817 23891 23851
rect 24777 23817 24811 23851
rect 25145 23817 25179 23851
rect 14841 23749 14875 23783
rect 17049 23749 17083 23783
rect 17601 23749 17635 23783
rect 21741 23749 21775 23783
rect 2237 23681 2271 23715
rect 1476 23613 1510 23647
rect 11320 23613 11354 23647
rect 13185 23613 13219 23647
rect 13737 23613 13771 23647
rect 14657 23613 14691 23647
rect 15209 23613 15243 23647
rect 15761 23613 15795 23647
rect 16313 23613 16347 23647
rect 16773 23613 16807 23647
rect 16865 23613 16899 23647
rect 18153 23681 18187 23715
rect 21097 23681 21131 23715
rect 22569 23681 22603 23715
rect 22017 23613 22051 23647
rect 24501 23613 24535 23647
rect 24593 23613 24627 23647
rect 18245 23545 18279 23579
rect 18797 23545 18831 23579
rect 20453 23545 20487 23579
rect 20545 23545 20579 23579
rect 1547 23477 1581 23511
rect 11391 23477 11425 23511
rect 15945 23477 15979 23511
rect 17601 23477 17635 23511
rect 17877 23477 17911 23511
rect 20269 23477 20303 23511
rect 13875 23273 13909 23307
rect 16175 23273 16209 23307
rect 18153 23273 18187 23307
rect 20269 23273 20303 23307
rect 21373 23273 21407 23307
rect 22017 23273 22051 23307
rect 22615 23273 22649 23307
rect 23719 23273 23753 23307
rect 24777 23273 24811 23307
rect 12863 23205 12897 23239
rect 17785 23205 17819 23239
rect 19349 23205 19383 23239
rect 13772 23137 13806 23171
rect 16037 23137 16071 23171
rect 17141 23137 17175 23171
rect 21005 23137 21039 23171
rect 22477 23137 22511 23171
rect 23489 23137 23523 23171
rect 24593 23137 24627 23171
rect 19257 23069 19291 23103
rect 19809 23001 19843 23035
rect 12633 22933 12667 22967
rect 14565 22933 14599 22967
rect 18429 22933 18463 22967
rect 13415 22729 13449 22763
rect 21189 22729 21223 22763
rect 24685 22729 24719 22763
rect 25421 22729 25455 22763
rect 15669 22661 15703 22695
rect 20453 22661 20487 22695
rect 14565 22593 14599 22627
rect 16221 22593 16255 22627
rect 18797 22593 18831 22627
rect 19717 22593 19751 22627
rect 21373 22593 21407 22627
rect 24041 22593 24075 22627
rect 13312 22525 13346 22559
rect 13737 22525 13771 22559
rect 21465 22525 21499 22559
rect 25237 22525 25271 22559
rect 25789 22525 25823 22559
rect 14657 22457 14691 22491
rect 15209 22457 15243 22491
rect 16313 22457 16347 22491
rect 16865 22457 16899 22491
rect 18153 22457 18187 22491
rect 18245 22457 18279 22491
rect 19901 22457 19935 22491
rect 19993 22457 20027 22491
rect 22477 22457 22511 22491
rect 23765 22457 23799 22491
rect 23857 22457 23891 22491
rect 12817 22389 12851 22423
rect 14289 22389 14323 22423
rect 16037 22389 16071 22423
rect 17141 22389 17175 22423
rect 17785 22389 17819 22423
rect 19257 22389 19291 22423
rect 20821 22389 20855 22423
rect 23121 22389 23155 22423
rect 23489 22389 23523 22423
rect 13737 22185 13771 22219
rect 14197 22185 14231 22219
rect 15439 22185 15473 22219
rect 16221 22185 16255 22219
rect 19533 22185 19567 22219
rect 23765 22185 23799 22219
rect 17049 22117 17083 22151
rect 18061 22117 18095 22151
rect 21097 22117 21131 22151
rect 22661 22117 22695 22151
rect 23213 22117 23247 22151
rect 24041 22117 24075 22151
rect 15368 22049 15402 22083
rect 16405 22049 16439 22083
rect 19876 22049 19910 22083
rect 24133 22049 24167 22083
rect 17969 21981 18003 22015
rect 18245 21981 18279 22015
rect 21005 21981 21039 22015
rect 21649 21981 21683 22015
rect 22569 21981 22603 22015
rect 19165 21845 19199 21879
rect 19947 21845 19981 21879
rect 21925 21845 21959 21879
rect 18245 21641 18279 21675
rect 20085 21641 20119 21675
rect 20821 21641 20855 21675
rect 24133 21641 24167 21675
rect 24777 21641 24811 21675
rect 15991 21573 16025 21607
rect 22569 21573 22603 21607
rect 23305 21573 23339 21607
rect 14289 21505 14323 21539
rect 18705 21505 18739 21539
rect 21051 21505 21085 21539
rect 22017 21505 22051 21539
rect 14197 21437 14231 21471
rect 14933 21437 14967 21471
rect 15888 21437 15922 21471
rect 19165 21437 19199 21471
rect 20964 21437 20998 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 16681 21369 16715 21403
rect 19486 21369 19520 21403
rect 22109 21369 22143 21403
rect 15301 21301 15335 21335
rect 16405 21301 16439 21335
rect 19073 21301 19107 21335
rect 20453 21301 20487 21335
rect 21465 21301 21499 21335
rect 21741 21301 21775 21335
rect 22937 21301 22971 21335
rect 16221 21097 16255 21131
rect 16773 21097 16807 21131
rect 19441 21097 19475 21131
rect 20637 21097 20671 21131
rect 21649 21097 21683 21131
rect 22753 21097 22787 21131
rect 25513 21097 25547 21131
rect 13829 21029 13863 21063
rect 14381 21029 14415 21063
rect 18883 21029 18917 21063
rect 1444 20961 1478 20995
rect 11840 20961 11874 20995
rect 21281 20961 21315 20995
rect 23949 20961 23983 20995
rect 25329 20961 25363 20995
rect 13737 20893 13771 20927
rect 15853 20893 15887 20927
rect 18521 20893 18555 20927
rect 1547 20757 1581 20791
rect 11943 20757 11977 20791
rect 12817 20757 12851 20791
rect 13553 20757 13587 20791
rect 18245 20757 18279 20791
rect 19809 20757 19843 20791
rect 24041 20757 24075 20791
rect 1593 20553 1627 20587
rect 5549 20553 5583 20587
rect 11805 20553 11839 20587
rect 13921 20553 13955 20587
rect 15301 20553 15335 20587
rect 17141 20553 17175 20587
rect 20729 20553 20763 20587
rect 21097 20553 21131 20587
rect 22477 20553 22511 20587
rect 24041 20553 24075 20587
rect 14289 20485 14323 20519
rect 15761 20485 15795 20519
rect 16129 20485 16163 20519
rect 12909 20417 12943 20451
rect 18981 20417 19015 20451
rect 19809 20417 19843 20451
rect 23489 20417 23523 20451
rect 24225 20417 24259 20451
rect 5156 20349 5190 20383
rect 14381 20349 14415 20383
rect 16221 20349 16255 20383
rect 17417 20349 17451 20383
rect 18245 20349 18279 20383
rect 18705 20349 18739 20383
rect 21557 20349 21591 20383
rect 12725 20281 12759 20315
rect 13001 20281 13035 20315
rect 13553 20281 13587 20315
rect 14702 20281 14736 20315
rect 20171 20281 20205 20315
rect 21878 20281 21912 20315
rect 24317 20281 24351 20315
rect 24869 20281 24903 20315
rect 5227 20213 5261 20247
rect 16589 20213 16623 20247
rect 17877 20213 17911 20247
rect 19349 20213 19383 20247
rect 19625 20213 19659 20247
rect 21373 20213 21407 20247
rect 23121 20213 23155 20247
rect 25329 20213 25363 20247
rect 14473 20009 14507 20043
rect 15393 20009 15427 20043
rect 21327 20009 21361 20043
rect 25329 20009 25363 20043
rect 18061 19941 18095 19975
rect 19625 19941 19659 19975
rect 21649 19941 21683 19975
rect 22385 19941 22419 19975
rect 23949 19941 23983 19975
rect 24501 19941 24535 19975
rect 13277 19873 13311 19907
rect 15301 19873 15335 19907
rect 15761 19873 15795 19907
rect 16129 19873 16163 19907
rect 17325 19873 17359 19907
rect 17785 19873 17819 19907
rect 18889 19873 18923 19907
rect 19349 19873 19383 19907
rect 21256 19873 21290 19907
rect 15117 19805 15151 19839
rect 22293 19805 22327 19839
rect 22937 19805 22971 19839
rect 23857 19805 23891 19839
rect 13001 19669 13035 19703
rect 13645 19669 13679 19703
rect 16681 19669 16715 19703
rect 18429 19669 18463 19703
rect 18797 19669 18831 19703
rect 23213 19669 23247 19703
rect 16589 19465 16623 19499
rect 20085 19465 20119 19499
rect 25421 19465 25455 19499
rect 22707 19397 22741 19431
rect 14657 19329 14691 19363
rect 23029 19329 23063 19363
rect 24041 19329 24075 19363
rect 24685 19329 24719 19363
rect 13001 19261 13035 19295
rect 15577 19261 15611 19295
rect 15945 19261 15979 19295
rect 16313 19261 16347 19295
rect 17785 19261 17819 19295
rect 18705 19261 18739 19295
rect 19165 19261 19199 19295
rect 19441 19261 19475 19295
rect 20821 19261 20855 19295
rect 22636 19261 22670 19295
rect 25237 19261 25271 19295
rect 25789 19261 25823 19295
rect 12909 19193 12943 19227
rect 13322 19193 13356 19227
rect 15301 19193 15335 19227
rect 16865 19193 16899 19227
rect 20729 19193 20763 19227
rect 21183 19193 21217 19227
rect 23765 19193 23799 19227
rect 23857 19193 23891 19227
rect 13921 19125 13955 19159
rect 15025 19125 15059 19159
rect 17325 19125 17359 19159
rect 18521 19125 18555 19159
rect 19717 19125 19751 19159
rect 21741 19125 21775 19159
rect 22201 19125 22235 19159
rect 23397 19125 23431 19159
rect 13185 18921 13219 18955
rect 15117 18921 15151 18955
rect 16129 18921 16163 18955
rect 20637 18921 20671 18955
rect 21925 18921 21959 18955
rect 23397 18921 23431 18955
rect 23765 18921 23799 18955
rect 24777 18921 24811 18955
rect 13737 18853 13771 18887
rect 22798 18853 22832 18887
rect 15853 18785 15887 18819
rect 16313 18785 16347 18819
rect 16681 18785 16715 18819
rect 18705 18785 18739 18819
rect 19165 18785 19199 18819
rect 21005 18785 21039 18819
rect 21649 18785 21683 18819
rect 24593 18785 24627 18819
rect 13645 18717 13679 18751
rect 13921 18717 13955 18751
rect 19441 18717 19475 18751
rect 22477 18717 22511 18751
rect 15577 18581 15611 18615
rect 24225 18581 24259 18615
rect 3985 18377 4019 18411
rect 13645 18377 13679 18411
rect 19073 18377 19107 18411
rect 20085 18377 20119 18411
rect 22845 18377 22879 18411
rect 24777 18377 24811 18411
rect 17141 18309 17175 18343
rect 15945 18241 15979 18275
rect 16773 18241 16807 18275
rect 18613 18241 18647 18275
rect 21925 18241 21959 18275
rect 3592 18173 3626 18207
rect 15025 18173 15059 18207
rect 15853 18173 15887 18207
rect 16957 18173 16991 18207
rect 17417 18173 17451 18207
rect 18061 18173 18095 18207
rect 18521 18173 18555 18207
rect 24593 18173 24627 18207
rect 19441 18105 19475 18139
rect 20177 18105 20211 18139
rect 20729 18105 20763 18139
rect 21281 18105 21315 18139
rect 21373 18105 21407 18139
rect 3663 18037 3697 18071
rect 14013 18037 14047 18071
rect 14841 18037 14875 18071
rect 15117 18037 15151 18071
rect 16405 18037 16439 18071
rect 17785 18037 17819 18071
rect 21097 18037 21131 18071
rect 22477 18037 22511 18071
rect 24409 18037 24443 18071
rect 25145 18037 25179 18071
rect 18935 17833 18969 17867
rect 15117 17765 15151 17799
rect 21097 17765 21131 17799
rect 21649 17765 21683 17799
rect 22477 17765 22511 17799
rect 1444 17697 1478 17731
rect 16129 17697 16163 17731
rect 18797 17697 18831 17731
rect 19876 17697 19910 17731
rect 22569 17697 22603 17731
rect 24685 17697 24719 17731
rect 17601 17629 17635 17663
rect 21005 17629 21039 17663
rect 24041 17629 24075 17663
rect 1547 17493 1581 17527
rect 15853 17493 15887 17527
rect 16313 17493 16347 17527
rect 18061 17493 18095 17527
rect 19441 17493 19475 17527
rect 19947 17493 19981 17527
rect 1593 17289 1627 17323
rect 2421 17289 2455 17323
rect 15853 17289 15887 17323
rect 16221 17289 16255 17323
rect 20361 17289 20395 17323
rect 20729 17289 20763 17323
rect 20821 17289 20855 17323
rect 22569 17289 22603 17323
rect 23949 17289 23983 17323
rect 16957 17221 16991 17255
rect 16405 17153 16439 17187
rect 2028 17085 2062 17119
rect 12265 17085 12299 17119
rect 12633 17085 12667 17119
rect 14657 17085 14691 17119
rect 15393 17085 15427 17119
rect 19441 17085 19475 17119
rect 24685 17221 24719 17255
rect 21557 17153 21591 17187
rect 24133 17153 24167 17187
rect 25605 17153 25639 17187
rect 15485 17017 15519 17051
rect 16497 17017 16531 17051
rect 19349 17017 19383 17051
rect 19803 17017 19837 17051
rect 20821 17017 20855 17051
rect 21281 17017 21315 17051
rect 21373 17017 21407 17051
rect 24225 17017 24259 17051
rect 2099 16949 2133 16983
rect 13001 16949 13035 16983
rect 18889 16949 18923 16983
rect 21097 16949 21131 16983
rect 23397 16949 23431 16983
rect 16405 16745 16439 16779
rect 19901 16745 19935 16779
rect 20729 16745 20763 16779
rect 21925 16745 21959 16779
rect 24133 16745 24167 16779
rect 13001 16677 13035 16711
rect 13553 16677 13587 16711
rect 15485 16677 15519 16711
rect 17049 16677 17083 16711
rect 18975 16677 19009 16711
rect 21097 16677 21131 16711
rect 21649 16677 21683 16711
rect 23029 16677 23063 16711
rect 24593 16677 24627 16711
rect 11805 16541 11839 16575
rect 12909 16541 12943 16575
rect 15393 16541 15427 16575
rect 16037 16541 16071 16575
rect 16957 16541 16991 16575
rect 18613 16541 18647 16575
rect 21005 16541 21039 16575
rect 22937 16541 22971 16575
rect 23581 16541 23615 16575
rect 24501 16541 24535 16575
rect 24777 16541 24811 16575
rect 17509 16473 17543 16507
rect 19533 16473 19567 16507
rect 18337 16405 18371 16439
rect 12265 16201 12299 16235
rect 12725 16201 12759 16235
rect 14749 16201 14783 16235
rect 15485 16201 15519 16235
rect 16957 16201 16991 16235
rect 19349 16201 19383 16235
rect 21695 16201 21729 16235
rect 24869 16201 24903 16235
rect 25467 16201 25501 16235
rect 22477 16133 22511 16167
rect 13553 16065 13587 16099
rect 15761 16065 15795 16099
rect 16037 16065 16071 16099
rect 19073 16065 19107 16099
rect 20637 16065 20671 16099
rect 20913 16065 20947 16099
rect 21373 16065 21407 16099
rect 22707 16065 22741 16099
rect 23857 16065 23891 16099
rect 18337 15997 18371 16031
rect 18797 15997 18831 16031
rect 19809 15997 19843 16031
rect 20545 15997 20579 16031
rect 21624 15997 21658 16031
rect 22620 15997 22654 16031
rect 25396 15997 25430 16031
rect 12909 15929 12943 15963
rect 13001 15929 13035 15963
rect 15853 15929 15887 15963
rect 23949 15929 23983 15963
rect 24501 15929 24535 15963
rect 13829 15861 13863 15895
rect 15209 15861 15243 15895
rect 17325 15861 17359 15895
rect 17877 15861 17911 15895
rect 22109 15861 22143 15895
rect 23121 15861 23155 15895
rect 23489 15861 23523 15895
rect 25237 15861 25271 15895
rect 25881 15861 25915 15895
rect 12633 15657 12667 15691
rect 13461 15657 13495 15691
rect 14381 15657 14415 15691
rect 16865 15657 16899 15691
rect 17877 15657 17911 15691
rect 23305 15657 23339 15691
rect 25145 15657 25179 15691
rect 15663 15589 15697 15623
rect 22706 15589 22740 15623
rect 23581 15589 23615 15623
rect 24133 15589 24167 15623
rect 13185 15521 13219 15555
rect 14197 15521 14231 15555
rect 16221 15521 16255 15555
rect 17049 15521 17083 15555
rect 18337 15521 18371 15555
rect 18521 15521 18555 15555
rect 24777 15521 24811 15555
rect 12265 15453 12299 15487
rect 15301 15453 15335 15487
rect 18613 15453 18647 15487
rect 19073 15453 19107 15487
rect 22385 15453 22419 15487
rect 17233 15385 17267 15419
rect 16589 15317 16623 15351
rect 19993 15317 20027 15351
rect 21833 15317 21867 15351
rect 24041 15317 24075 15351
rect 12265 15113 12299 15147
rect 15577 15113 15611 15147
rect 15945 15113 15979 15147
rect 19165 15113 19199 15147
rect 22753 15113 22787 15147
rect 24961 15113 24995 15147
rect 11897 14977 11931 15011
rect 12909 14977 12943 15011
rect 17141 14977 17175 15011
rect 19993 14977 20027 15011
rect 20453 14977 20487 15011
rect 5432 14909 5466 14943
rect 5825 14909 5859 14943
rect 14657 14909 14691 14943
rect 16589 14909 16623 14943
rect 21833 14909 21867 14943
rect 24225 14909 24259 14943
rect 5641 14841 5675 14875
rect 12541 14841 12575 14875
rect 12633 14841 12667 14875
rect 14565 14841 14599 14875
rect 14979 14841 15013 14875
rect 16221 14841 16255 14875
rect 18245 14841 18279 14875
rect 18337 14841 18371 14875
rect 18889 14841 18923 14875
rect 19809 14841 19843 14875
rect 20085 14841 20119 14875
rect 21741 14841 21775 14875
rect 22195 14841 22229 14875
rect 23029 14841 23063 14875
rect 24685 14841 24719 14875
rect 13461 14773 13495 14807
rect 14197 14773 14231 14807
rect 17417 14773 17451 14807
rect 17877 14773 17911 14807
rect 25513 14773 25547 14807
rect 12265 14569 12299 14603
rect 17877 14569 17911 14603
rect 19809 14569 19843 14603
rect 22385 14569 22419 14603
rect 12633 14501 12667 14535
rect 18423 14501 18457 14535
rect 20913 14501 20947 14535
rect 23029 14501 23063 14535
rect 24501 14501 24535 14535
rect 24593 14501 24627 14535
rect 11529 14433 11563 14467
rect 14197 14433 14231 14467
rect 15669 14433 15703 14467
rect 16037 14433 16071 14467
rect 16865 14433 16899 14467
rect 21557 14433 21591 14467
rect 11621 14365 11655 14399
rect 12541 14365 12575 14399
rect 12909 14365 12943 14399
rect 18061 14365 18095 14399
rect 22937 14365 22971 14399
rect 23581 14365 23615 14399
rect 24777 14365 24811 14399
rect 17049 14297 17083 14331
rect 14381 14229 14415 14263
rect 14657 14229 14691 14263
rect 16497 14229 16531 14263
rect 18981 14229 19015 14263
rect 24225 14229 24259 14263
rect 10977 14025 11011 14059
rect 11805 14025 11839 14059
rect 13369 14025 13403 14059
rect 14197 14025 14231 14059
rect 17417 14025 17451 14059
rect 17877 14025 17911 14059
rect 18981 14025 19015 14059
rect 22477 14025 22511 14059
rect 23213 14025 23247 14059
rect 24041 14025 24075 14059
rect 25145 14025 25179 14059
rect 20453 13957 20487 13991
rect 24777 13957 24811 13991
rect 15301 13889 15335 13923
rect 17141 13889 17175 13923
rect 19257 13889 19291 13923
rect 22109 13889 22143 13923
rect 24225 13889 24259 13923
rect 25513 13889 25547 13923
rect 12449 13821 12483 13855
rect 14657 13821 14691 13855
rect 14749 13821 14783 13855
rect 15209 13821 15243 13855
rect 16313 13821 16347 13855
rect 16405 13821 16439 13855
rect 16865 13821 16899 13855
rect 18061 13821 18095 13855
rect 21649 13821 21683 13855
rect 21833 13821 21867 13855
rect 12770 13753 12804 13787
rect 18382 13753 18416 13787
rect 19901 13753 19935 13787
rect 19993 13753 20027 13787
rect 24317 13753 24351 13787
rect 12173 13685 12207 13719
rect 13645 13685 13679 13719
rect 15761 13685 15795 13719
rect 19717 13685 19751 13719
rect 20821 13685 20855 13719
rect 21189 13685 21223 13719
rect 22845 13685 22879 13719
rect 12357 13481 12391 13515
rect 15853 13481 15887 13515
rect 18153 13481 18187 13515
rect 22845 13481 22879 13515
rect 23397 13481 23431 13515
rect 14381 13413 14415 13447
rect 17417 13413 17451 13447
rect 18429 13413 18463 13447
rect 19165 13413 19199 13447
rect 21649 13413 21683 13447
rect 24409 13413 24443 13447
rect 12265 13345 12299 13379
rect 12633 13345 12667 13379
rect 13921 13345 13955 13379
rect 14197 13345 14231 13379
rect 15669 13345 15703 13379
rect 16681 13345 16715 13379
rect 17141 13345 17175 13379
rect 20913 13345 20947 13379
rect 21373 13345 21407 13379
rect 19073 13277 19107 13311
rect 19349 13277 19383 13311
rect 19993 13277 20027 13311
rect 22477 13277 22511 13311
rect 24317 13277 24351 13311
rect 24593 13277 24627 13311
rect 13093 13141 13127 13175
rect 13461 13141 13495 13175
rect 14841 13141 14875 13175
rect 16129 13141 16163 13175
rect 16497 13141 16531 13175
rect 21925 13141 21959 13175
rect 12633 12937 12667 12971
rect 14565 12937 14599 12971
rect 15669 12937 15703 12971
rect 16681 12937 16715 12971
rect 17417 12937 17451 12971
rect 19165 12937 19199 12971
rect 22753 12937 22787 12971
rect 12173 12869 12207 12903
rect 16175 12869 16209 12903
rect 16313 12869 16347 12903
rect 19533 12869 19567 12903
rect 11345 12801 11379 12835
rect 13645 12801 13679 12835
rect 13921 12801 13955 12835
rect 16405 12801 16439 12835
rect 21005 12801 21039 12835
rect 21833 12801 21867 12835
rect 24409 12801 24443 12835
rect 24685 12801 24719 12835
rect 12449 12733 12483 12767
rect 12909 12733 12943 12767
rect 15301 12733 15335 12767
rect 16037 12733 16071 12767
rect 18153 12733 18187 12767
rect 20269 12733 20303 12767
rect 20729 12733 20763 12767
rect 23489 12733 23523 12767
rect 23765 12733 23799 12767
rect 13737 12665 13771 12699
rect 20085 12665 20119 12699
rect 21281 12665 21315 12699
rect 22154 12665 22188 12699
rect 11253 12597 11287 12631
rect 13369 12597 13403 12631
rect 15025 12597 15059 12631
rect 17049 12597 17083 12631
rect 17877 12597 17911 12631
rect 18521 12597 18555 12631
rect 21649 12597 21683 12631
rect 23029 12597 23063 12631
rect 25145 12597 25179 12631
rect 14749 12393 14783 12427
rect 15945 12393 15979 12427
rect 16681 12393 16715 12427
rect 17325 12393 17359 12427
rect 18797 12393 18831 12427
rect 25559 12393 25593 12427
rect 12541 12325 12575 12359
rect 13553 12325 13587 12359
rect 15301 12325 15335 12359
rect 16405 12325 16439 12359
rect 21741 12325 21775 12359
rect 22477 12325 22511 12359
rect 11805 12257 11839 12291
rect 12357 12257 12391 12291
rect 17141 12257 17175 12291
rect 17601 12257 17635 12291
rect 18153 12257 18187 12291
rect 18383 12257 18417 12291
rect 21189 12257 21223 12291
rect 21465 12257 21499 12291
rect 24501 12257 24535 12291
rect 25488 12257 25522 12291
rect 13461 12189 13495 12223
rect 13921 12189 13955 12223
rect 15117 12189 15151 12223
rect 15669 12189 15703 12223
rect 18521 12189 18555 12223
rect 20269 12121 20303 12155
rect 12817 12053 12851 12087
rect 13185 12053 13219 12087
rect 15439 12053 15473 12087
rect 15577 12053 15611 12087
rect 18061 12053 18095 12087
rect 18291 12053 18325 12087
rect 19165 12053 19199 12087
rect 20637 12053 20671 12087
rect 24133 12053 24167 12087
rect 11805 11849 11839 11883
rect 14822 11849 14856 11883
rect 16497 11849 16531 11883
rect 16865 11849 16899 11883
rect 18521 11849 18555 11883
rect 19073 11849 19107 11883
rect 20361 11849 20395 11883
rect 21557 11849 21591 11883
rect 24133 11849 24167 11883
rect 25513 11849 25547 11883
rect 13553 11781 13587 11815
rect 14565 11781 14599 11815
rect 14933 11781 14967 11815
rect 18337 11781 18371 11815
rect 19441 11781 19475 11815
rect 11529 11713 11563 11747
rect 14197 11713 14231 11747
rect 15025 11713 15059 11747
rect 16589 11713 16623 11747
rect 18429 11713 18463 11747
rect 19809 11713 19843 11747
rect 24593 11713 24627 11747
rect 10701 11645 10735 11679
rect 10885 11645 10919 11679
rect 12633 11645 12667 11679
rect 15393 11645 15427 11679
rect 16368 11645 16402 11679
rect 18208 11645 18242 11679
rect 20545 11645 20579 11679
rect 21005 11645 21039 11679
rect 12954 11577 12988 11611
rect 14657 11577 14691 11611
rect 16221 11577 16255 11611
rect 17509 11577 17543 11611
rect 18061 11577 18095 11611
rect 21281 11577 21315 11611
rect 22569 11577 22603 11611
rect 24317 11577 24351 11611
rect 24409 11577 24443 11611
rect 12265 11509 12299 11543
rect 15669 11509 15703 11543
rect 16129 11509 16163 11543
rect 17785 11509 17819 11543
rect 23397 11509 23431 11543
rect 11897 11305 11931 11339
rect 13461 11305 13495 11339
rect 13645 11305 13679 11339
rect 14749 11305 14783 11339
rect 15761 11305 15795 11339
rect 21097 11305 21131 11339
rect 21649 11305 21683 11339
rect 22201 11305 22235 11339
rect 24317 11305 24351 11339
rect 12173 11237 12207 11271
rect 15117 11237 15151 11271
rect 16221 11237 16255 11271
rect 19073 11237 19107 11271
rect 23121 11237 23155 11271
rect 23213 11237 23247 11271
rect 24777 11237 24811 11271
rect 1444 11169 1478 11203
rect 13553 11169 13587 11203
rect 14105 11169 14139 11203
rect 15301 11169 15335 11203
rect 16865 11169 16899 11203
rect 18337 11169 18371 11203
rect 12081 11101 12115 11135
rect 12725 11101 12759 11135
rect 16773 11101 16807 11135
rect 18705 11101 18739 11135
rect 21281 11101 21315 11135
rect 23765 11101 23799 11135
rect 24685 11101 24719 11135
rect 24961 11101 24995 11135
rect 18475 11033 18509 11067
rect 1547 10965 1581 10999
rect 15485 10965 15519 10999
rect 16681 10965 16715 10999
rect 17877 10965 17911 10999
rect 18153 10965 18187 10999
rect 18613 10965 18647 10999
rect 20637 10965 20671 10999
rect 1593 10761 1627 10795
rect 13645 10761 13679 10795
rect 15485 10761 15519 10795
rect 17693 10761 17727 10795
rect 18337 10761 18371 10795
rect 18705 10761 18739 10795
rect 23029 10761 23063 10795
rect 24777 10761 24811 10795
rect 10701 10693 10735 10727
rect 12265 10693 12299 10727
rect 15163 10693 15197 10727
rect 15301 10693 15335 10727
rect 17141 10693 17175 10727
rect 15393 10625 15427 10659
rect 10793 10557 10827 10591
rect 11345 10557 11379 10591
rect 11529 10557 11563 10591
rect 12449 10557 12483 10591
rect 14565 10557 14599 10591
rect 15025 10557 15059 10591
rect 16497 10557 16531 10591
rect 16957 10557 16991 10591
rect 11897 10489 11931 10523
rect 12770 10489 12804 10523
rect 14197 10489 14231 10523
rect 17509 10489 17543 10523
rect 18199 10693 18233 10727
rect 22753 10693 22787 10727
rect 25789 10693 25823 10727
rect 18429 10625 18463 10659
rect 24041 10625 24075 10659
rect 25053 10625 25087 10659
rect 20545 10557 20579 10591
rect 20729 10557 20763 10591
rect 21005 10557 21039 10591
rect 21833 10557 21867 10591
rect 25304 10557 25338 10591
rect 18061 10489 18095 10523
rect 22154 10489 22188 10523
rect 23765 10489 23799 10523
rect 23857 10489 23891 10523
rect 13369 10421 13403 10455
rect 14841 10421 14875 10455
rect 16037 10421 16071 10455
rect 16773 10421 16807 10455
rect 17693 10421 17727 10455
rect 17785 10421 17819 10455
rect 19165 10421 19199 10455
rect 19533 10421 19567 10455
rect 19901 10421 19935 10455
rect 21281 10421 21315 10455
rect 21649 10421 21683 10455
rect 23397 10421 23431 10455
rect 25375 10421 25409 10455
rect 10885 10217 10919 10251
rect 12081 10217 12115 10251
rect 12449 10217 12483 10251
rect 13737 10217 13771 10251
rect 14381 10217 14415 10251
rect 14657 10217 14691 10251
rect 15025 10217 15059 10251
rect 16865 10217 16899 10251
rect 17877 10217 17911 10251
rect 20361 10217 20395 10251
rect 22293 10217 22327 10251
rect 23581 10217 23615 10251
rect 24547 10217 24581 10251
rect 12817 10149 12851 10183
rect 19073 10149 19107 10183
rect 20637 10149 20671 10183
rect 21925 10149 21959 10183
rect 23305 10149 23339 10183
rect 24041 10149 24075 10183
rect 14197 10081 14231 10115
rect 15301 10081 15335 10115
rect 15448 10081 15482 10115
rect 17325 10081 17359 10115
rect 18337 10081 18371 10115
rect 20913 10081 20947 10115
rect 21373 10081 21407 10115
rect 23029 10081 23063 10115
rect 24476 10081 24510 10115
rect 25488 10081 25522 10115
rect 12725 10013 12759 10047
rect 13001 10013 13035 10047
rect 15669 10013 15703 10047
rect 18705 10013 18739 10047
rect 21465 10013 21499 10047
rect 17509 9945 17543 9979
rect 18502 9945 18536 9979
rect 15577 9877 15611 9911
rect 15761 9877 15795 9911
rect 16497 9877 16531 9911
rect 18245 9877 18279 9911
rect 18613 9877 18647 9911
rect 19349 9877 19383 9911
rect 25559 9877 25593 9911
rect 14381 9673 14415 9707
rect 14979 9673 15013 9707
rect 16221 9673 16255 9707
rect 16865 9673 16899 9707
rect 19625 9673 19659 9707
rect 20453 9673 20487 9707
rect 21649 9673 21683 9707
rect 22661 9673 22695 9707
rect 24685 9673 24719 9707
rect 25375 9673 25409 9707
rect 26157 9673 26191 9707
rect 13921 9605 13955 9639
rect 15117 9605 15151 9639
rect 16681 9605 16715 9639
rect 18429 9605 18463 9639
rect 13185 9537 13219 9571
rect 13461 9537 13495 9571
rect 14749 9537 14783 9571
rect 15209 9537 15243 9571
rect 16773 9537 16807 9571
rect 17877 9537 17911 9571
rect 18521 9537 18555 9571
rect 21281 9537 21315 9571
rect 25789 9537 25823 9571
rect 12265 9469 12299 9503
rect 13093 9469 13127 9503
rect 14841 9469 14875 9503
rect 16405 9469 16439 9503
rect 16552 9469 16586 9503
rect 18300 9469 18334 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 21189 9469 21223 9503
rect 23489 9469 23523 9503
rect 23765 9469 23799 9503
rect 25304 9469 25338 9503
rect 18153 9401 18187 9435
rect 18889 9401 18923 9435
rect 11897 9333 11931 9367
rect 15485 9333 15519 9367
rect 15945 9333 15979 9367
rect 17417 9333 17451 9367
rect 19165 9333 19199 9367
rect 23949 9333 23983 9367
rect 12081 9129 12115 9163
rect 14105 9129 14139 9163
rect 14381 9129 14415 9163
rect 16497 9129 16531 9163
rect 17233 9129 17267 9163
rect 17509 9129 17543 9163
rect 18797 9129 18831 9163
rect 19993 9129 20027 9163
rect 20729 9129 20763 9163
rect 21189 9129 21223 9163
rect 15301 9061 15335 9095
rect 22293 9061 22327 9095
rect 23765 9061 23799 9095
rect 23857 9061 23891 9095
rect 25237 9061 25271 9095
rect 12265 8993 12299 9027
rect 12541 8993 12575 9027
rect 14197 8993 14231 9027
rect 15448 8993 15482 9027
rect 18061 8993 18095 9027
rect 18337 8993 18371 9027
rect 15669 8925 15703 8959
rect 22201 8925 22235 8959
rect 24409 8925 24443 8959
rect 24685 8925 24719 8959
rect 15761 8857 15795 8891
rect 17877 8857 17911 8891
rect 22753 8857 22787 8891
rect 8677 8789 8711 8823
rect 13001 8789 13035 8823
rect 14933 8789 14967 8823
rect 15577 8789 15611 8823
rect 16865 8789 16899 8823
rect 19257 8789 19291 8823
rect 19717 8789 19751 8823
rect 11253 8585 11287 8619
rect 11897 8585 11931 8619
rect 15761 8585 15795 8619
rect 16129 8585 16163 8619
rect 19901 8585 19935 8619
rect 20269 8585 20303 8619
rect 22201 8585 22235 8619
rect 22477 8585 22511 8619
rect 23489 8585 23523 8619
rect 24961 8585 24995 8619
rect 25559 8585 25593 8619
rect 15393 8517 15427 8551
rect 19349 8517 19383 8551
rect 9045 8449 9079 8483
rect 11345 8449 11379 8483
rect 12541 8449 12575 8483
rect 12909 8449 12943 8483
rect 13829 8449 13863 8483
rect 16497 8449 16531 8483
rect 8677 8381 8711 8415
rect 9229 8381 9263 8415
rect 14289 8381 14323 8415
rect 14565 8381 14599 8415
rect 15577 8381 15611 8415
rect 16589 8381 16623 8415
rect 16773 8381 16807 8415
rect 18705 8381 18739 8415
rect 19533 8449 19567 8483
rect 19993 8449 20027 8483
rect 21281 8449 21315 8483
rect 22845 8449 22879 8483
rect 23949 8449 23983 8483
rect 24593 8449 24627 8483
rect 19772 8381 19806 8415
rect 20637 8381 20671 8415
rect 21189 8381 21223 8415
rect 25488 8381 25522 8415
rect 12633 8313 12667 8347
rect 13553 8313 13587 8347
rect 19165 8313 19199 8347
rect 19349 8313 19383 8347
rect 19624 8313 19658 8347
rect 21643 8313 21677 8347
rect 24041 8313 24075 8347
rect 8585 8245 8619 8279
rect 12173 8245 12207 8279
rect 14105 8245 14139 8279
rect 16865 8245 16899 8279
rect 17509 8245 17543 8279
rect 17785 8245 17819 8279
rect 18337 8245 18371 8279
rect 25973 8245 26007 8279
rect 12449 8041 12483 8075
rect 14381 8041 14415 8075
rect 14749 8041 14783 8075
rect 15117 8041 15151 8075
rect 16405 8041 16439 8075
rect 18245 8041 18279 8075
rect 21373 8041 21407 8075
rect 23949 8041 23983 8075
rect 8769 7973 8803 8007
rect 11253 7973 11287 8007
rect 22246 7973 22280 8007
rect 24225 7973 24259 8007
rect 24317 7973 24351 8007
rect 8217 7905 8251 7939
rect 8401 7905 8435 7939
rect 10609 7905 10643 7939
rect 12081 7905 12115 7939
rect 14197 7905 14231 7939
rect 15301 7905 15335 7939
rect 15761 7905 15795 7939
rect 17601 7905 17635 7939
rect 18613 7905 18647 7939
rect 19349 7905 19383 7939
rect 19717 7905 19751 7939
rect 21925 7905 21959 7939
rect 14105 7837 14139 7871
rect 16037 7837 16071 7871
rect 17969 7837 18003 7871
rect 19993 7837 20027 7871
rect 24593 7837 24627 7871
rect 13001 7701 13035 7735
rect 17509 7701 17543 7735
rect 17766 7701 17800 7735
rect 17877 7701 17911 7735
rect 22845 7701 22879 7735
rect 10609 7497 10643 7531
rect 11805 7497 11839 7531
rect 12173 7497 12207 7531
rect 15025 7497 15059 7531
rect 16957 7497 16991 7531
rect 19349 7497 19383 7531
rect 19625 7497 19659 7531
rect 20453 7497 20487 7531
rect 20821 7497 20855 7531
rect 22385 7497 22419 7531
rect 23489 7497 23523 7531
rect 25467 7497 25501 7531
rect 17601 7429 17635 7463
rect 7941 7361 7975 7395
rect 8493 7361 8527 7395
rect 13001 7361 13035 7395
rect 24501 7361 24535 7395
rect 24777 7361 24811 7395
rect 1444 7293 1478 7327
rect 1869 7293 1903 7327
rect 8677 7293 8711 7327
rect 15485 7293 15519 7327
rect 15945 7293 15979 7327
rect 18153 7293 18187 7327
rect 21005 7293 21039 7327
rect 21465 7293 21499 7327
rect 24041 7293 24075 7327
rect 25396 7293 25430 7327
rect 25881 7293 25915 7327
rect 1547 7225 1581 7259
rect 12725 7225 12759 7259
rect 12817 7225 12851 7259
rect 15301 7225 15335 7259
rect 16221 7225 16255 7259
rect 21741 7225 21775 7259
rect 8309 7157 8343 7191
rect 13645 7157 13679 7191
rect 14289 7157 14323 7191
rect 17233 7157 17267 7191
rect 18337 7157 18371 7191
rect 22017 7157 22051 7191
rect 12173 6953 12207 6987
rect 12909 6953 12943 6987
rect 15577 6953 15611 6987
rect 15853 6953 15887 6987
rect 18797 6953 18831 6987
rect 23857 6953 23891 6987
rect 16450 6885 16484 6919
rect 18198 6885 18232 6919
rect 22706 6885 22740 6919
rect 11897 6817 11931 6851
rect 12357 6817 12391 6851
rect 13737 6817 13771 6851
rect 14105 6817 14139 6851
rect 16129 6817 16163 6851
rect 17877 6817 17911 6851
rect 22385 6817 22419 6851
rect 23305 6817 23339 6851
rect 24225 6817 24259 6851
rect 14197 6749 14231 6783
rect 24133 6749 24167 6783
rect 8493 6613 8527 6647
rect 17049 6613 17083 6647
rect 17693 6613 17727 6647
rect 11989 6409 12023 6443
rect 13185 6409 13219 6443
rect 15853 6409 15887 6443
rect 19441 6409 19475 6443
rect 22385 6409 22419 6443
rect 22707 6409 22741 6443
rect 23029 6409 23063 6443
rect 24041 6409 24075 6443
rect 12633 6341 12667 6375
rect 13553 6341 13587 6375
rect 18705 6341 18739 6375
rect 25145 6341 25179 6375
rect 14013 6273 14047 6307
rect 16497 6273 16531 6307
rect 18153 6273 18187 6307
rect 19073 6273 19107 6307
rect 19625 6273 19659 6307
rect 24501 6273 24535 6307
rect 22109 6205 22143 6239
rect 22604 6205 22638 6239
rect 13829 6137 13863 6171
rect 14334 6137 14368 6171
rect 16129 6137 16163 6171
rect 16589 6137 16623 6171
rect 17141 6137 17175 6171
rect 17509 6137 17543 6171
rect 18245 6137 18279 6171
rect 21557 6137 21591 6171
rect 23397 6137 23431 6171
rect 24225 6137 24259 6171
rect 24317 6137 24351 6171
rect 14933 6069 14967 6103
rect 17785 6069 17819 6103
rect 14657 5865 14691 5899
rect 16773 5865 16807 5899
rect 13829 5797 13863 5831
rect 17877 5797 17911 5831
rect 17969 5797 18003 5831
rect 18521 5797 18555 5831
rect 22706 5797 22740 5831
rect 24409 5797 24443 5831
rect 14381 5729 14415 5763
rect 15393 5729 15427 5763
rect 22385 5729 22419 5763
rect 12633 5661 12667 5695
rect 13737 5661 13771 5695
rect 15301 5661 15335 5695
rect 24317 5661 24351 5695
rect 24593 5661 24627 5695
rect 16497 5593 16531 5627
rect 23305 5525 23339 5559
rect 12955 5321 12989 5355
rect 15117 5321 15151 5355
rect 17509 5321 17543 5355
rect 22385 5321 22419 5355
rect 22753 5321 22787 5355
rect 23489 5321 23523 5355
rect 24961 5321 24995 5355
rect 26065 5321 26099 5355
rect 15393 5253 15427 5287
rect 13829 5185 13863 5219
rect 15945 5185 15979 5219
rect 18429 5185 18463 5219
rect 19073 5185 19107 5219
rect 12884 5117 12918 5151
rect 13369 5117 13403 5151
rect 14749 5117 14783 5151
rect 24041 5117 24075 5151
rect 25580 5117 25614 5151
rect 13645 5049 13679 5083
rect 15669 5049 15703 5083
rect 15761 5049 15795 5083
rect 18153 5049 18187 5083
rect 18245 5049 18279 5083
rect 14197 4981 14231 5015
rect 16589 4981 16623 5015
rect 16957 4981 16991 5015
rect 17785 4981 17819 5015
rect 24409 4981 24443 5015
rect 25651 4981 25685 5015
rect 14657 4777 14691 4811
rect 16313 4777 16347 4811
rect 17785 4777 17819 4811
rect 18337 4777 18371 4811
rect 19027 4777 19061 4811
rect 24041 4777 24075 4811
rect 13829 4709 13863 4743
rect 24501 4709 24535 4743
rect 25053 4709 25087 4743
rect 1476 4641 1510 4675
rect 15393 4641 15427 4675
rect 17417 4641 17451 4675
rect 18889 4641 18923 4675
rect 13737 4573 13771 4607
rect 14381 4573 14415 4607
rect 15301 4573 15335 4607
rect 24409 4573 24443 4607
rect 1547 4505 1581 4539
rect 1593 4233 1627 4267
rect 14013 4233 14047 4267
rect 15853 4233 15887 4267
rect 17417 4233 17451 4267
rect 18981 4233 19015 4267
rect 24133 4233 24167 4267
rect 25237 4233 25271 4267
rect 13737 4097 13771 4131
rect 15209 4097 15243 4131
rect 24685 4097 24719 4131
rect 12265 4029 12299 4063
rect 12541 4029 12575 4063
rect 14933 3961 14967 3995
rect 15025 3961 15059 3995
rect 23489 3961 23523 3995
rect 24317 3961 24351 3995
rect 24409 3961 24443 3995
rect 12909 3893 12943 3927
rect 14749 3893 14783 3927
rect 13001 3689 13035 3723
rect 14933 3689 14967 3723
rect 15439 3689 15473 3723
rect 24225 3689 24259 3723
rect 24731 3689 24765 3723
rect 12443 3621 12477 3655
rect 12081 3553 12115 3587
rect 15209 3553 15243 3587
rect 13369 3349 13403 3383
rect 24501 3349 24535 3383
rect 11805 3145 11839 3179
rect 15393 3145 15427 3179
rect 12173 3009 12207 3043
rect 12817 3009 12851 3043
rect 13277 3009 13311 3043
rect 12909 2873 12943 2907
rect 13737 2873 13771 2907
rect 24685 2805 24719 2839
rect 12449 2601 12483 2635
rect 14335 2601 14369 2635
rect 24731 2601 24765 2635
rect 12817 2533 12851 2567
rect 1476 2465 1510 2499
rect 1869 2465 1903 2499
rect 14264 2465 14298 2499
rect 24660 2465 24694 2499
rect 12725 2397 12759 2431
rect 14749 2397 14783 2431
rect 1547 2329 1581 2363
rect 11989 2329 12023 2363
rect 13277 2329 13311 2363
rect 25145 2261 25179 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 24765 25483 24823 25489
rect 24765 25449 24777 25483
rect 24811 25480 24823 25483
rect 27154 25480 27160 25492
rect 24811 25452 27160 25480
rect 24811 25449 24823 25452
rect 24765 25443 24823 25449
rect 27154 25440 27160 25452
rect 27212 25440 27218 25492
rect 24581 25347 24639 25353
rect 24581 25313 24593 25347
rect 24627 25344 24639 25347
rect 24670 25344 24676 25356
rect 24627 25316 24676 25344
rect 24627 25313 24639 25316
rect 24581 25307 24639 25313
rect 24670 25304 24676 25316
rect 24728 25304 24734 25356
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 24765 24939 24823 24945
rect 24765 24905 24777 24939
rect 24811 24936 24823 24939
rect 25590 24936 25596 24948
rect 24811 24908 25596 24936
rect 24811 24905 24823 24908
rect 24765 24899 24823 24905
rect 25590 24896 25596 24908
rect 25648 24896 25654 24948
rect 18463 24871 18521 24877
rect 18463 24837 18475 24871
rect 18509 24868 18521 24871
rect 18874 24868 18880 24880
rect 18509 24840 18880 24868
rect 18509 24837 18521 24840
rect 18463 24831 18521 24837
rect 18874 24828 18880 24840
rect 18932 24828 18938 24880
rect 22695 24871 22753 24877
rect 22695 24837 22707 24871
rect 22741 24868 22753 24871
rect 25222 24868 25228 24880
rect 22741 24840 25228 24868
rect 22741 24837 22753 24840
rect 22695 24831 22753 24837
rect 25222 24828 25228 24840
rect 25280 24828 25286 24880
rect 18392 24735 18450 24741
rect 18392 24701 18404 24735
rect 18438 24732 18450 24735
rect 19426 24732 19432 24744
rect 19484 24741 19490 24744
rect 19484 24735 19522 24741
rect 18438 24704 18828 24732
rect 19374 24704 19432 24732
rect 18438 24701 18450 24704
rect 18392 24695 18450 24701
rect 18800 24676 18828 24704
rect 19426 24692 19432 24704
rect 19510 24732 19522 24735
rect 19889 24735 19947 24741
rect 19889 24732 19901 24735
rect 19510 24704 19901 24732
rect 19510 24701 19522 24704
rect 19484 24695 19522 24701
rect 19889 24701 19901 24704
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 22624 24735 22682 24741
rect 22624 24701 22636 24735
rect 22670 24732 22682 24735
rect 22670 24704 23152 24732
rect 22670 24701 22682 24704
rect 22624 24695 22682 24701
rect 19484 24692 19490 24695
rect 18782 24664 18788 24676
rect 18743 24636 18788 24664
rect 18782 24624 18788 24636
rect 18840 24624 18846 24676
rect 19567 24667 19625 24673
rect 19567 24633 19579 24667
rect 19613 24664 19625 24667
rect 20346 24664 20352 24676
rect 19613 24636 20352 24664
rect 19613 24633 19625 24636
rect 19567 24627 19625 24633
rect 20346 24624 20352 24636
rect 20404 24624 20410 24676
rect 16942 24596 16948 24608
rect 16903 24568 16948 24596
rect 16942 24556 16948 24568
rect 17000 24556 17006 24608
rect 20441 24599 20499 24605
rect 20441 24565 20453 24599
rect 20487 24596 20499 24599
rect 20990 24596 20996 24608
rect 20487 24568 20996 24596
rect 20487 24565 20499 24568
rect 20441 24559 20499 24565
rect 20990 24556 20996 24568
rect 21048 24556 21054 24608
rect 23124 24605 23152 24704
rect 24210 24692 24216 24744
rect 24268 24732 24274 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24268 24704 24593 24732
rect 24268 24692 24274 24704
rect 24581 24701 24593 24704
rect 24627 24732 24639 24735
rect 25133 24735 25191 24741
rect 25133 24732 25145 24735
rect 24627 24704 25145 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 25133 24701 25145 24704
rect 25179 24701 25191 24735
rect 25133 24695 25191 24701
rect 23109 24599 23167 24605
rect 23109 24565 23121 24599
rect 23155 24596 23167 24599
rect 23198 24596 23204 24608
rect 23155 24568 23204 24596
rect 23155 24565 23167 24568
rect 23109 24559 23167 24565
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 23808 24568 24409 24596
rect 23808 24556 23814 24568
rect 24397 24565 24409 24568
rect 24443 24596 24455 24599
rect 24670 24596 24676 24608
rect 24443 24568 24676 24596
rect 24443 24565 24455 24568
rect 24397 24559 24455 24565
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24361 15531 24395
rect 15473 24355 15531 24361
rect 18325 24395 18383 24401
rect 18325 24361 18337 24395
rect 18371 24392 18383 24395
rect 22462 24392 22468 24404
rect 18371 24364 22468 24392
rect 18371 24361 18383 24364
rect 18325 24355 18383 24361
rect 15488 24324 15516 24355
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 20622 24324 20628 24336
rect 15488 24296 20628 24324
rect 20622 24284 20628 24296
rect 20680 24284 20686 24336
rect 21082 24324 21088 24336
rect 21043 24296 21088 24324
rect 21082 24284 21088 24296
rect 21140 24284 21146 24336
rect 750 24216 756 24268
rect 808 24256 814 24268
rect 1432 24259 1490 24265
rect 1432 24256 1444 24259
rect 808 24228 1444 24256
rect 808 24216 814 24228
rect 1432 24225 1444 24228
rect 1478 24256 1490 24259
rect 1854 24256 1860 24268
rect 1478 24228 1860 24256
rect 1478 24225 1490 24228
rect 1432 24219 1490 24225
rect 1854 24216 1860 24228
rect 1912 24216 1918 24268
rect 12964 24259 13022 24265
rect 12964 24225 12976 24259
rect 13010 24256 13022 24259
rect 13170 24256 13176 24268
rect 13010 24228 13176 24256
rect 13010 24225 13022 24228
rect 12964 24219 13022 24225
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 15286 24256 15292 24268
rect 15247 24228 15292 24256
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 17196 24259 17254 24265
rect 17196 24225 17208 24259
rect 17242 24256 17254 24259
rect 17402 24256 17408 24268
rect 17242 24228 17408 24256
rect 17242 24225 17254 24228
rect 17196 24219 17254 24225
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 18141 24259 18199 24265
rect 18141 24225 18153 24259
rect 18187 24225 18199 24259
rect 18141 24219 18199 24225
rect 17267 24123 17325 24129
rect 17267 24089 17279 24123
rect 17313 24120 17325 24123
rect 18156 24120 18184 24219
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 19150 24256 19156 24268
rect 18656 24228 19156 24256
rect 18656 24216 18662 24228
rect 19150 24216 19156 24228
rect 19208 24256 19214 24268
rect 19280 24259 19338 24265
rect 19280 24256 19292 24259
rect 19208 24228 19292 24256
rect 19208 24216 19214 24228
rect 19280 24225 19292 24228
rect 19326 24225 19338 24259
rect 22462 24256 22468 24268
rect 22423 24228 22468 24256
rect 19280 24219 19338 24225
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 23636 24259 23694 24265
rect 23636 24225 23648 24259
rect 23682 24256 23694 24259
rect 23842 24256 23848 24268
rect 23682 24228 23848 24256
rect 23682 24225 23694 24228
rect 23636 24219 23694 24225
rect 23842 24216 23848 24228
rect 23900 24216 23906 24268
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 25130 24256 25136 24268
rect 24627 24228 25136 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 20990 24188 20996 24200
rect 20951 24160 20996 24188
rect 20990 24148 20996 24160
rect 21048 24148 21054 24200
rect 21266 24188 21272 24200
rect 21227 24160 21272 24188
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 18693 24123 18751 24129
rect 18693 24120 18705 24123
rect 17313 24092 18705 24120
rect 17313 24089 17325 24092
rect 17267 24083 17325 24089
rect 18693 24089 18705 24092
rect 18739 24089 18751 24123
rect 18693 24083 18751 24089
rect 22603 24123 22661 24129
rect 22603 24089 22615 24123
rect 22649 24120 22661 24123
rect 24118 24120 24124 24132
rect 22649 24092 24124 24120
rect 22649 24089 22661 24092
rect 22603 24083 22661 24089
rect 24118 24080 24124 24092
rect 24176 24080 24182 24132
rect 1535 24055 1593 24061
rect 1535 24021 1547 24055
rect 1581 24052 1593 24055
rect 2682 24052 2688 24064
rect 1581 24024 2688 24052
rect 1581 24021 1593 24024
rect 1535 24015 1593 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 13035 24055 13093 24061
rect 13035 24021 13047 24055
rect 13081 24052 13093 24055
rect 13262 24052 13268 24064
rect 13081 24024 13268 24052
rect 13081 24021 13093 24024
rect 13035 24015 13093 24021
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 19242 24012 19248 24064
rect 19300 24052 19306 24064
rect 19383 24055 19441 24061
rect 19383 24052 19395 24055
rect 19300 24024 19395 24052
rect 19300 24012 19306 24024
rect 19383 24021 19395 24024
rect 19429 24021 19441 24055
rect 20438 24052 20444 24064
rect 20399 24024 20444 24052
rect 19383 24015 19441 24021
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 20530 24012 20536 24064
rect 20588 24052 20594 24064
rect 23707 24055 23765 24061
rect 23707 24052 23719 24055
rect 20588 24024 23719 24052
rect 20588 24012 20594 24024
rect 23707 24021 23719 24024
rect 23753 24021 23765 24055
rect 23707 24015 23765 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1854 23848 1860 23860
rect 1815 23820 1860 23848
rect 1854 23808 1860 23820
rect 1912 23808 1918 23860
rect 11698 23848 11704 23860
rect 11659 23820 11704 23848
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 12989 23851 13047 23857
rect 12989 23817 13001 23851
rect 13035 23848 13047 23851
rect 13170 23848 13176 23860
rect 13035 23820 13176 23848
rect 13035 23817 13047 23820
rect 12989 23811 13047 23817
rect 13170 23808 13176 23820
rect 13228 23808 13234 23860
rect 13357 23851 13415 23857
rect 13357 23817 13369 23851
rect 13403 23848 13415 23851
rect 14734 23848 14740 23860
rect 13403 23820 14740 23848
rect 13403 23817 13415 23820
rect 13357 23811 13415 23817
rect 14734 23808 14740 23820
rect 14792 23808 14798 23860
rect 15286 23808 15292 23860
rect 15344 23848 15350 23860
rect 15562 23848 15568 23860
rect 15344 23820 15568 23848
rect 15344 23808 15350 23820
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 17402 23848 17408 23860
rect 17363 23820 17408 23848
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 19150 23808 19156 23860
rect 19208 23848 19214 23860
rect 19245 23851 19303 23857
rect 19245 23848 19257 23851
rect 19208 23820 19257 23848
rect 19208 23808 19214 23820
rect 19245 23817 19257 23820
rect 19291 23817 19303 23851
rect 19245 23811 19303 23817
rect 21082 23808 21088 23860
rect 21140 23848 21146 23860
rect 21358 23848 21364 23860
rect 21140 23820 21364 23848
rect 21140 23808 21146 23820
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23848 22247 23851
rect 23658 23848 23664 23860
rect 22235 23820 23664 23848
rect 22235 23817 22247 23820
rect 22189 23811 22247 23817
rect 23658 23808 23664 23820
rect 23716 23808 23722 23860
rect 23842 23848 23848 23860
rect 23803 23820 23848 23848
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 24946 23848 24952 23860
rect 24811 23820 24952 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 24946 23808 24952 23820
rect 25004 23808 25010 23860
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 14829 23783 14887 23789
rect 14829 23749 14841 23783
rect 14875 23780 14887 23783
rect 15930 23780 15936 23792
rect 14875 23752 15936 23780
rect 14875 23749 14887 23752
rect 14829 23743 14887 23749
rect 15930 23740 15936 23752
rect 15988 23740 15994 23792
rect 17037 23783 17095 23789
rect 17037 23749 17049 23783
rect 17083 23780 17095 23783
rect 17494 23780 17500 23792
rect 17083 23752 17500 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 17494 23740 17500 23752
rect 17552 23740 17558 23792
rect 17589 23783 17647 23789
rect 17589 23749 17601 23783
rect 17635 23780 17647 23783
rect 19334 23780 19340 23792
rect 17635 23752 19340 23780
rect 17635 23749 17647 23752
rect 17589 23743 17647 23749
rect 19334 23740 19340 23752
rect 19392 23740 19398 23792
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 21729 23783 21787 23789
rect 21729 23780 21741 23783
rect 21048 23752 21741 23780
rect 21048 23740 21054 23752
rect 21729 23749 21741 23752
rect 21775 23749 21787 23783
rect 21729 23743 21787 23749
rect 1302 23672 1308 23724
rect 1360 23712 1366 23724
rect 2225 23715 2283 23721
rect 2225 23712 2237 23715
rect 1360 23684 2237 23712
rect 1360 23672 1366 23684
rect 1479 23653 1507 23684
rect 2225 23681 2237 23684
rect 2271 23681 2283 23715
rect 2225 23675 2283 23681
rect 16942 23672 16948 23724
rect 17000 23712 17006 23724
rect 18138 23712 18144 23724
rect 17000 23684 18144 23712
rect 17000 23672 17006 23684
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21266 23712 21272 23724
rect 21131 23684 21272 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21266 23672 21272 23684
rect 21324 23712 21330 23724
rect 22462 23712 22468 23724
rect 21324 23684 22468 23712
rect 21324 23672 21330 23684
rect 22462 23672 22468 23684
rect 22520 23712 22526 23724
rect 22557 23715 22615 23721
rect 22557 23712 22569 23715
rect 22520 23684 22569 23712
rect 22520 23672 22526 23684
rect 22557 23681 22569 23684
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 1464 23647 1522 23653
rect 1464 23613 1476 23647
rect 1510 23613 1522 23647
rect 1464 23607 1522 23613
rect 11308 23647 11366 23653
rect 11308 23613 11320 23647
rect 11354 23644 11366 23647
rect 11698 23644 11704 23656
rect 11354 23616 11704 23644
rect 11354 23613 11366 23616
rect 11308 23607 11366 23613
rect 11698 23604 11704 23616
rect 11756 23604 11762 23656
rect 13173 23647 13231 23653
rect 13173 23613 13185 23647
rect 13219 23644 13231 23647
rect 13538 23644 13544 23656
rect 13219 23616 13544 23644
rect 13219 23613 13231 23616
rect 13173 23607 13231 23613
rect 13538 23604 13544 23616
rect 13596 23644 13602 23656
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 13596 23616 13737 23644
rect 13596 23604 13602 23616
rect 13725 23613 13737 23616
rect 13771 23613 13783 23647
rect 13725 23607 13783 23613
rect 14645 23647 14703 23653
rect 14645 23613 14657 23647
rect 14691 23644 14703 23647
rect 15197 23647 15255 23653
rect 15197 23644 15209 23647
rect 14691 23616 15209 23644
rect 14691 23613 14703 23616
rect 14645 23607 14703 23613
rect 15197 23613 15209 23616
rect 15243 23644 15255 23647
rect 15286 23644 15292 23656
rect 15243 23616 15292 23644
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 15286 23604 15292 23616
rect 15344 23604 15350 23656
rect 15746 23644 15752 23656
rect 15659 23616 15752 23644
rect 15746 23604 15752 23616
rect 15804 23644 15810 23656
rect 16301 23647 16359 23653
rect 16301 23644 16313 23647
rect 15804 23616 16313 23644
rect 15804 23604 15810 23616
rect 16301 23613 16313 23616
rect 16347 23613 16359 23647
rect 16301 23607 16359 23613
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16724 23616 16773 23644
rect 16724 23604 16730 23616
rect 16761 23613 16773 23616
rect 16807 23644 16819 23647
rect 16853 23647 16911 23653
rect 16853 23644 16865 23647
rect 16807 23616 16865 23644
rect 16807 23613 16819 23616
rect 16761 23607 16819 23613
rect 16853 23613 16865 23616
rect 16899 23613 16911 23647
rect 22002 23644 22008 23656
rect 21963 23616 22008 23644
rect 16853 23607 16911 23613
rect 22002 23604 22008 23616
rect 22060 23604 22066 23656
rect 24394 23604 24400 23656
rect 24452 23644 24458 23656
rect 24489 23647 24547 23653
rect 24489 23644 24501 23647
rect 24452 23616 24501 23644
rect 24452 23604 24458 23616
rect 24489 23613 24501 23616
rect 24535 23644 24547 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 24535 23616 24593 23644
rect 24535 23613 24547 23616
rect 24489 23607 24547 23613
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 18233 23579 18291 23585
rect 18233 23545 18245 23579
rect 18279 23545 18291 23579
rect 18782 23576 18788 23588
rect 18743 23548 18788 23576
rect 18233 23539 18291 23545
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1762 23508 1768 23520
rect 1581 23480 1768 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1762 23468 1768 23480
rect 1820 23468 1826 23520
rect 11379 23511 11437 23517
rect 11379 23477 11391 23511
rect 11425 23508 11437 23511
rect 14734 23508 14740 23520
rect 11425 23480 14740 23508
rect 11425 23477 11437 23480
rect 11379 23471 11437 23477
rect 14734 23468 14740 23480
rect 14792 23468 14798 23520
rect 15933 23511 15991 23517
rect 15933 23477 15945 23511
rect 15979 23508 15991 23511
rect 17589 23511 17647 23517
rect 17589 23508 17601 23511
rect 15979 23480 17601 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 17589 23477 17601 23480
rect 17635 23477 17647 23511
rect 17589 23471 17647 23477
rect 17770 23468 17776 23520
rect 17828 23508 17834 23520
rect 17865 23511 17923 23517
rect 17865 23508 17877 23511
rect 17828 23480 17877 23508
rect 17828 23468 17834 23480
rect 17865 23477 17877 23480
rect 17911 23508 17923 23511
rect 18248 23508 18276 23539
rect 18782 23536 18788 23548
rect 18840 23536 18846 23588
rect 20438 23576 20444 23588
rect 20351 23548 20444 23576
rect 20438 23536 20444 23548
rect 20496 23536 20502 23588
rect 20533 23579 20591 23585
rect 20533 23545 20545 23579
rect 20579 23545 20591 23579
rect 20533 23539 20591 23545
rect 17911 23480 18276 23508
rect 20257 23511 20315 23517
rect 17911 23477 17923 23480
rect 17865 23471 17923 23477
rect 20257 23477 20269 23511
rect 20303 23508 20315 23511
rect 20548 23508 20576 23539
rect 20990 23508 20996 23520
rect 20303 23480 20996 23508
rect 20303 23477 20315 23480
rect 20257 23471 20315 23477
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 13863 23307 13921 23313
rect 13863 23273 13875 23307
rect 13909 23304 13921 23307
rect 15562 23304 15568 23316
rect 13909 23276 15568 23304
rect 13909 23273 13921 23276
rect 13863 23267 13921 23273
rect 15562 23264 15568 23276
rect 15620 23264 15626 23316
rect 16163 23307 16221 23313
rect 16163 23273 16175 23307
rect 16209 23304 16221 23307
rect 16666 23304 16672 23316
rect 16209 23276 16672 23304
rect 16209 23273 16221 23276
rect 16163 23267 16221 23273
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 18138 23304 18144 23316
rect 18099 23276 18144 23304
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 20257 23307 20315 23313
rect 20257 23273 20269 23307
rect 20303 23304 20315 23307
rect 20530 23304 20536 23316
rect 20303 23276 20536 23304
rect 20303 23273 20315 23276
rect 20257 23267 20315 23273
rect 12851 23239 12909 23245
rect 12851 23205 12863 23239
rect 12897 23236 12909 23239
rect 15746 23236 15752 23248
rect 12897 23208 15752 23236
rect 12897 23205 12909 23208
rect 12851 23199 12909 23205
rect 15746 23196 15752 23208
rect 15804 23196 15810 23248
rect 17770 23236 17776 23248
rect 17731 23208 17776 23236
rect 17770 23196 17776 23208
rect 17828 23196 17834 23248
rect 19337 23239 19395 23245
rect 19337 23205 19349 23239
rect 19383 23236 19395 23239
rect 19426 23236 19432 23248
rect 19383 23208 19432 23236
rect 19383 23205 19395 23208
rect 19337 23199 19395 23205
rect 19426 23196 19432 23208
rect 19484 23196 19490 23248
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 20272 23236 20300 23267
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 21358 23304 21364 23316
rect 21319 23276 21364 23304
rect 21358 23264 21364 23276
rect 21416 23264 21422 23316
rect 22002 23304 22008 23316
rect 21963 23276 22008 23304
rect 22002 23264 22008 23276
rect 22060 23304 22066 23316
rect 22603 23307 22661 23313
rect 22603 23304 22615 23307
rect 22060 23276 22615 23304
rect 22060 23264 22066 23276
rect 22603 23273 22615 23276
rect 22649 23273 22661 23307
rect 22603 23267 22661 23273
rect 23707 23307 23765 23313
rect 23707 23273 23719 23307
rect 23753 23304 23765 23307
rect 24210 23304 24216 23316
rect 23753 23276 24216 23304
rect 23753 23273 23765 23276
rect 23707 23267 23765 23273
rect 24210 23264 24216 23276
rect 24268 23264 24274 23316
rect 24765 23307 24823 23313
rect 24765 23273 24777 23307
rect 24811 23304 24823 23307
rect 25498 23304 25504 23316
rect 24811 23276 25504 23304
rect 24811 23273 24823 23276
rect 24765 23267 24823 23273
rect 25498 23264 25504 23276
rect 25556 23264 25562 23316
rect 19944 23208 20300 23236
rect 19944 23196 19950 23208
rect 13630 23128 13636 23180
rect 13688 23168 13694 23180
rect 13760 23171 13818 23177
rect 13760 23168 13772 23171
rect 13688 23140 13772 23168
rect 13688 23128 13694 23140
rect 13760 23137 13772 23140
rect 13806 23137 13818 23171
rect 13760 23131 13818 23137
rect 16025 23171 16083 23177
rect 16025 23137 16037 23171
rect 16071 23168 16083 23171
rect 16114 23168 16120 23180
rect 16071 23140 16120 23168
rect 16071 23137 16083 23140
rect 16025 23131 16083 23137
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 17126 23168 17132 23180
rect 17087 23140 17132 23168
rect 17126 23128 17132 23140
rect 17184 23128 17190 23180
rect 20990 23168 20996 23180
rect 20951 23140 20996 23168
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 22462 23168 22468 23180
rect 22423 23140 22468 23168
rect 22462 23128 22468 23140
rect 22520 23128 22526 23180
rect 23106 23128 23112 23180
rect 23164 23168 23170 23180
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 23164 23140 23489 23168
rect 23164 23128 23170 23140
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 24118 23128 24124 23180
rect 24176 23168 24182 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 24176 23140 24593 23168
rect 24176 23128 24182 23140
rect 24581 23137 24593 23140
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 19242 23100 19248 23112
rect 19155 23072 19248 23100
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 19797 23035 19855 23041
rect 19797 23032 19809 23035
rect 19707 23004 19809 23032
rect 19797 23001 19809 23004
rect 19843 23032 19855 23035
rect 20438 23032 20444 23044
rect 19843 23004 20444 23032
rect 19843 23001 19855 23004
rect 19797 22995 19855 23001
rect 20438 22992 20444 23004
rect 20496 22992 20502 23044
rect 12621 22967 12679 22973
rect 12621 22933 12633 22967
rect 12667 22964 12679 22967
rect 12802 22964 12808 22976
rect 12667 22936 12808 22964
rect 12667 22933 12679 22936
rect 12621 22927 12679 22933
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 14550 22964 14556 22976
rect 14511 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 18138 22924 18144 22976
rect 18196 22964 18202 22976
rect 18417 22967 18475 22973
rect 18417 22964 18429 22967
rect 18196 22936 18429 22964
rect 18196 22924 18202 22936
rect 18417 22933 18429 22936
rect 18463 22933 18475 22967
rect 18417 22927 18475 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 13403 22763 13461 22769
rect 13403 22729 13415 22763
rect 13449 22760 13461 22763
rect 13538 22760 13544 22772
rect 13449 22732 13544 22760
rect 13449 22729 13461 22732
rect 13403 22723 13461 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 19484 22732 21189 22760
rect 19484 22720 19490 22732
rect 21177 22729 21189 22732
rect 21223 22760 21235 22763
rect 24670 22760 24676 22772
rect 21223 22732 21496 22760
rect 24631 22732 24676 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 15657 22695 15715 22701
rect 15657 22661 15669 22695
rect 15703 22692 15715 22695
rect 16114 22692 16120 22704
rect 15703 22664 16120 22692
rect 15703 22661 15715 22664
rect 15657 22655 15715 22661
rect 16114 22652 16120 22664
rect 16172 22652 16178 22704
rect 20438 22692 20444 22704
rect 20399 22664 20444 22692
rect 20438 22652 20444 22664
rect 20496 22652 20502 22704
rect 14550 22624 14556 22636
rect 14511 22596 14556 22624
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 14734 22584 14740 22636
rect 14792 22624 14798 22636
rect 16206 22624 16212 22636
rect 14792 22596 16212 22624
rect 14792 22584 14798 22596
rect 16206 22584 16212 22596
rect 16264 22584 16270 22636
rect 18782 22624 18788 22636
rect 18743 22596 18788 22624
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 19978 22624 19984 22636
rect 19751 22596 19984 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 19978 22584 19984 22596
rect 20036 22624 20042 22636
rect 21361 22627 21419 22633
rect 21361 22624 21373 22627
rect 20036 22596 21373 22624
rect 20036 22584 20042 22596
rect 21361 22593 21373 22596
rect 21407 22593 21419 22627
rect 21361 22587 21419 22593
rect 13078 22516 13084 22568
rect 13136 22556 13142 22568
rect 21468 22565 21496 22732
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 25406 22760 25412 22772
rect 25367 22732 25412 22760
rect 25406 22720 25412 22732
rect 25464 22720 25470 22772
rect 23198 22584 23204 22636
rect 23256 22624 23262 22636
rect 24029 22627 24087 22633
rect 24029 22624 24041 22627
rect 23256 22596 24041 22624
rect 23256 22584 23262 22596
rect 24029 22593 24041 22596
rect 24075 22593 24087 22627
rect 24029 22587 24087 22593
rect 13300 22559 13358 22565
rect 13300 22556 13312 22559
rect 13136 22528 13312 22556
rect 13136 22516 13142 22528
rect 13300 22525 13312 22528
rect 13346 22556 13358 22559
rect 13725 22559 13783 22565
rect 13725 22556 13737 22559
rect 13346 22528 13737 22556
rect 13346 22525 13358 22528
rect 13300 22519 13358 22525
rect 13725 22525 13737 22528
rect 13771 22525 13783 22559
rect 13725 22519 13783 22525
rect 21453 22559 21511 22565
rect 21453 22525 21465 22559
rect 21499 22525 21511 22559
rect 25222 22556 25228 22568
rect 25183 22528 25228 22556
rect 21453 22519 21511 22525
rect 25222 22516 25228 22528
rect 25280 22556 25286 22568
rect 25777 22559 25835 22565
rect 25777 22556 25789 22559
rect 25280 22528 25789 22556
rect 25280 22516 25286 22528
rect 25777 22525 25789 22528
rect 25823 22525 25835 22559
rect 25777 22519 25835 22525
rect 14645 22491 14703 22497
rect 14645 22457 14657 22491
rect 14691 22457 14703 22491
rect 14645 22451 14703 22457
rect 15197 22491 15255 22497
rect 15197 22457 15209 22491
rect 15243 22488 15255 22491
rect 15378 22488 15384 22500
rect 15243 22460 15384 22488
rect 15243 22457 15255 22460
rect 15197 22451 15255 22457
rect 12802 22420 12808 22432
rect 12763 22392 12808 22420
rect 12802 22380 12808 22392
rect 12860 22380 12866 22432
rect 14274 22420 14280 22432
rect 14235 22392 14280 22420
rect 14274 22380 14280 22392
rect 14332 22420 14338 22432
rect 14660 22420 14688 22451
rect 15378 22448 15384 22460
rect 15436 22448 15442 22500
rect 16301 22491 16359 22497
rect 16301 22457 16313 22491
rect 16347 22488 16359 22491
rect 16390 22488 16396 22500
rect 16347 22460 16396 22488
rect 16347 22457 16359 22460
rect 16301 22451 16359 22457
rect 14332 22392 14688 22420
rect 16025 22423 16083 22429
rect 14332 22380 14338 22392
rect 16025 22389 16037 22423
rect 16071 22420 16083 22423
rect 16316 22420 16344 22451
rect 16390 22448 16396 22460
rect 16448 22448 16454 22500
rect 16853 22491 16911 22497
rect 16853 22457 16865 22491
rect 16899 22488 16911 22491
rect 18138 22488 18144 22500
rect 16899 22460 18144 22488
rect 16899 22457 16911 22460
rect 16853 22451 16911 22457
rect 18138 22448 18144 22460
rect 18196 22448 18202 22500
rect 18233 22491 18291 22497
rect 18233 22457 18245 22491
rect 18279 22457 18291 22491
rect 19886 22488 19892 22500
rect 19847 22460 19892 22488
rect 18233 22451 18291 22457
rect 17126 22420 17132 22432
rect 16071 22392 16344 22420
rect 17087 22392 17132 22420
rect 16071 22389 16083 22392
rect 16025 22383 16083 22389
rect 17126 22380 17132 22392
rect 17184 22420 17190 22432
rect 17773 22423 17831 22429
rect 17773 22420 17785 22423
rect 17184 22392 17785 22420
rect 17184 22380 17190 22392
rect 17773 22389 17785 22392
rect 17819 22420 17831 22423
rect 18248 22420 18276 22451
rect 19886 22448 19892 22460
rect 19944 22448 19950 22500
rect 19978 22448 19984 22500
rect 20036 22488 20042 22500
rect 20036 22460 20081 22488
rect 20036 22448 20042 22460
rect 20530 22448 20536 22500
rect 20588 22488 20594 22500
rect 22462 22488 22468 22500
rect 20588 22460 22468 22488
rect 20588 22448 20594 22460
rect 22462 22448 22468 22460
rect 22520 22448 22526 22500
rect 23750 22488 23756 22500
rect 23711 22460 23756 22488
rect 23750 22448 23756 22460
rect 23808 22448 23814 22500
rect 23842 22448 23848 22500
rect 23900 22488 23906 22500
rect 23900 22460 23945 22488
rect 23900 22448 23906 22460
rect 17819 22392 18276 22420
rect 19245 22423 19303 22429
rect 17819 22389 17831 22392
rect 17773 22383 17831 22389
rect 19245 22389 19257 22423
rect 19291 22420 19303 22423
rect 19426 22420 19432 22432
rect 19291 22392 19432 22420
rect 19291 22389 19303 22392
rect 19245 22383 19303 22389
rect 19426 22380 19432 22392
rect 19484 22380 19490 22432
rect 20070 22380 20076 22432
rect 20128 22420 20134 22432
rect 20809 22423 20867 22429
rect 20809 22420 20821 22423
rect 20128 22392 20821 22420
rect 20128 22380 20134 22392
rect 20809 22389 20821 22392
rect 20855 22420 20867 22423
rect 20990 22420 20996 22432
rect 20855 22392 20996 22420
rect 20855 22389 20867 22392
rect 20809 22383 20867 22389
rect 20990 22380 20996 22392
rect 21048 22380 21054 22432
rect 23106 22420 23112 22432
rect 23067 22392 23112 22420
rect 23106 22380 23112 22392
rect 23164 22380 23170 22432
rect 23477 22423 23535 22429
rect 23477 22389 23489 22423
rect 23523 22420 23535 22423
rect 23860 22420 23888 22448
rect 23523 22392 23888 22420
rect 23523 22389 23535 22392
rect 23477 22383 23535 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 13630 22176 13636 22228
rect 13688 22216 13694 22228
rect 13725 22219 13783 22225
rect 13725 22216 13737 22219
rect 13688 22188 13737 22216
rect 13688 22176 13694 22188
rect 13725 22185 13737 22188
rect 13771 22185 13783 22219
rect 13725 22179 13783 22185
rect 14185 22219 14243 22225
rect 14185 22185 14197 22219
rect 14231 22216 14243 22219
rect 14550 22216 14556 22228
rect 14231 22188 14556 22216
rect 14231 22185 14243 22188
rect 14185 22179 14243 22185
rect 14550 22176 14556 22188
rect 14608 22176 14614 22228
rect 15286 22176 15292 22228
rect 15344 22216 15350 22228
rect 15427 22219 15485 22225
rect 15427 22216 15439 22219
rect 15344 22188 15439 22216
rect 15344 22176 15350 22188
rect 15427 22185 15439 22188
rect 15473 22185 15485 22219
rect 16206 22216 16212 22228
rect 16167 22188 16212 22216
rect 15427 22179 15485 22185
rect 16206 22176 16212 22188
rect 16264 22176 16270 22228
rect 19518 22216 19524 22228
rect 19479 22188 19524 22216
rect 19518 22176 19524 22188
rect 19576 22176 19582 22228
rect 23750 22216 23756 22228
rect 23711 22188 23756 22216
rect 23750 22176 23756 22188
rect 23808 22176 23814 22228
rect 17037 22151 17095 22157
rect 17037 22117 17049 22151
rect 17083 22148 17095 22151
rect 18049 22151 18107 22157
rect 18049 22148 18061 22151
rect 17083 22120 18061 22148
rect 17083 22117 17095 22120
rect 17037 22111 17095 22117
rect 18049 22117 18061 22120
rect 18095 22148 18107 22151
rect 18230 22148 18236 22160
rect 18095 22120 18236 22148
rect 18095 22117 18107 22120
rect 18049 22111 18107 22117
rect 18230 22108 18236 22120
rect 18288 22108 18294 22160
rect 21082 22148 21088 22160
rect 21043 22120 21088 22148
rect 21082 22108 21088 22120
rect 21140 22108 21146 22160
rect 22646 22148 22652 22160
rect 22607 22120 22652 22148
rect 22646 22108 22652 22120
rect 22704 22108 22710 22160
rect 23198 22148 23204 22160
rect 23159 22120 23204 22148
rect 23198 22108 23204 22120
rect 23256 22108 23262 22160
rect 23842 22108 23848 22160
rect 23900 22148 23906 22160
rect 24029 22151 24087 22157
rect 24029 22148 24041 22151
rect 23900 22120 24041 22148
rect 23900 22108 23906 22120
rect 24029 22117 24041 22120
rect 24075 22117 24087 22151
rect 24029 22111 24087 22117
rect 15356 22083 15414 22089
rect 15356 22049 15368 22083
rect 15402 22080 15414 22083
rect 15470 22080 15476 22092
rect 15402 22052 15476 22080
rect 15402 22049 15414 22052
rect 15356 22043 15414 22049
rect 15470 22040 15476 22052
rect 15528 22040 15534 22092
rect 16390 22080 16396 22092
rect 16351 22052 16396 22080
rect 16390 22040 16396 22052
rect 16448 22040 16454 22092
rect 19864 22083 19922 22089
rect 19864 22049 19876 22083
rect 19910 22080 19922 22083
rect 20806 22080 20812 22092
rect 19910 22052 20812 22080
rect 19910 22049 19922 22052
rect 19864 22043 19922 22049
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 24118 22080 24124 22092
rect 24079 22052 24124 22080
rect 24118 22040 24124 22052
rect 24176 22040 24182 22092
rect 17954 22012 17960 22024
rect 17915 21984 17960 22012
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18138 21972 18144 22024
rect 18196 22012 18202 22024
rect 18233 22015 18291 22021
rect 18233 22012 18245 22015
rect 18196 21984 18245 22012
rect 18196 21972 18202 21984
rect 18233 21981 18245 21984
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 20346 21972 20352 22024
rect 20404 22012 20410 22024
rect 20993 22015 21051 22021
rect 20993 22012 21005 22015
rect 20404 21984 21005 22012
rect 20404 21972 20410 21984
rect 20993 21981 21005 21984
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 22012 21695 22015
rect 22554 22012 22560 22024
rect 21683 21984 22560 22012
rect 21683 21981 21695 21984
rect 21637 21975 21695 21981
rect 22554 21972 22560 21984
rect 22612 21972 22618 22024
rect 19150 21876 19156 21888
rect 19111 21848 19156 21876
rect 19150 21836 19156 21848
rect 19208 21836 19214 21888
rect 19935 21879 19993 21885
rect 19935 21845 19947 21879
rect 19981 21876 19993 21879
rect 21913 21879 21971 21885
rect 21913 21876 21925 21879
rect 19981 21848 21925 21876
rect 19981 21845 19993 21848
rect 19935 21839 19993 21845
rect 21913 21845 21925 21848
rect 21959 21876 21971 21879
rect 22002 21876 22008 21888
rect 21959 21848 22008 21876
rect 21959 21845 21971 21848
rect 21913 21839 21971 21845
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22738 21836 22744 21888
rect 22796 21876 22802 21888
rect 23750 21876 23756 21888
rect 22796 21848 23756 21876
rect 22796 21836 22802 21848
rect 23750 21836 23756 21848
rect 23808 21836 23814 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 18230 21672 18236 21684
rect 18191 21644 18236 21672
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 20070 21672 20076 21684
rect 20031 21644 20076 21672
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 20809 21675 20867 21681
rect 20809 21641 20821 21675
rect 20855 21672 20867 21675
rect 21082 21672 21088 21684
rect 20855 21644 21088 21672
rect 20855 21641 20867 21644
rect 20809 21635 20867 21641
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 22646 21632 22652 21684
rect 22704 21672 22710 21684
rect 24118 21672 24124 21684
rect 22704 21644 24124 21672
rect 22704 21632 22710 21644
rect 24118 21632 24124 21644
rect 24176 21632 24182 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 15979 21607 16037 21613
rect 15979 21573 15991 21607
rect 16025 21604 16037 21607
rect 19702 21604 19708 21616
rect 16025 21576 19708 21604
rect 16025 21573 16037 21576
rect 15979 21567 16037 21573
rect 19702 21564 19708 21576
rect 19760 21564 19766 21616
rect 22554 21604 22560 21616
rect 22515 21576 22560 21604
rect 22554 21564 22560 21576
rect 22612 21604 22618 21616
rect 23293 21607 23351 21613
rect 23293 21604 23305 21607
rect 22612 21576 23305 21604
rect 22612 21564 22618 21576
rect 23293 21573 23305 21576
rect 23339 21573 23351 21607
rect 23293 21567 23351 21573
rect 14274 21536 14280 21548
rect 14235 21508 14280 21536
rect 14274 21496 14280 21508
rect 14332 21496 14338 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 18012 21508 18705 21536
rect 18012 21496 18018 21508
rect 18693 21505 18705 21508
rect 18739 21536 18751 21539
rect 21039 21539 21097 21545
rect 21039 21536 21051 21539
rect 18739 21508 21051 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 21039 21505 21051 21508
rect 21085 21505 21097 21539
rect 22002 21536 22008 21548
rect 21963 21508 22008 21536
rect 21039 21499 21097 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 14185 21471 14243 21477
rect 14185 21437 14197 21471
rect 14231 21468 14243 21471
rect 14921 21471 14979 21477
rect 14921 21468 14933 21471
rect 14231 21440 14933 21468
rect 14231 21437 14243 21440
rect 14185 21431 14243 21437
rect 14921 21437 14933 21440
rect 14967 21468 14979 21471
rect 15286 21468 15292 21480
rect 14967 21440 15292 21468
rect 14967 21437 14979 21440
rect 14921 21431 14979 21437
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 15876 21471 15934 21477
rect 15876 21437 15888 21471
rect 15922 21437 15934 21471
rect 15876 21431 15934 21437
rect 14366 21360 14372 21412
rect 14424 21400 14430 21412
rect 15378 21400 15384 21412
rect 14424 21372 15384 21400
rect 14424 21360 14430 21372
rect 15378 21360 15384 21372
rect 15436 21400 15442 21412
rect 15891 21400 15919 21431
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 19150 21468 19156 21480
rect 18104 21440 19156 21468
rect 18104 21428 18110 21440
rect 19150 21428 19156 21440
rect 19208 21428 19214 21480
rect 20952 21471 21010 21477
rect 20952 21437 20964 21471
rect 20998 21468 21010 21471
rect 20998 21440 21496 21468
rect 20998 21437 21010 21440
rect 20952 21431 21010 21437
rect 16669 21403 16727 21409
rect 16669 21400 16681 21403
rect 15436 21372 16681 21400
rect 15436 21360 15442 21372
rect 16669 21369 16681 21372
rect 16715 21369 16727 21403
rect 19474 21403 19532 21409
rect 19474 21400 19486 21403
rect 16669 21363 16727 21369
rect 19352 21372 19486 21400
rect 19352 21344 19380 21372
rect 19474 21369 19486 21372
rect 19520 21369 19532 21403
rect 19474 21363 19532 21369
rect 21468 21344 21496 21440
rect 24210 21428 24216 21480
rect 24268 21468 24274 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 24268 21440 24593 21468
rect 24268 21428 24274 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24627 21440 25145 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 22097 21403 22155 21409
rect 22097 21369 22109 21403
rect 22143 21369 22155 21403
rect 22097 21363 22155 21369
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 15289 21335 15347 21341
rect 15289 21332 15301 21335
rect 14516 21304 15301 21332
rect 14516 21292 14522 21304
rect 15289 21301 15301 21304
rect 15335 21332 15347 21335
rect 15470 21332 15476 21344
rect 15335 21304 15476 21332
rect 15335 21301 15347 21304
rect 15289 21295 15347 21301
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16390 21332 16396 21344
rect 16351 21304 16396 21332
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 19061 21335 19119 21341
rect 19061 21301 19073 21335
rect 19107 21332 19119 21335
rect 19334 21332 19340 21344
rect 19107 21304 19340 21332
rect 19107 21301 19119 21304
rect 19061 21295 19119 21301
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 20441 21335 20499 21341
rect 20441 21301 20453 21335
rect 20487 21332 20499 21335
rect 20806 21332 20812 21344
rect 20487 21304 20812 21332
rect 20487 21301 20499 21304
rect 20441 21295 20499 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 21450 21332 21456 21344
rect 21411 21304 21456 21332
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 21726 21332 21732 21344
rect 21687 21304 21732 21332
rect 21726 21292 21732 21304
rect 21784 21332 21790 21344
rect 22112 21332 22140 21363
rect 21784 21304 22140 21332
rect 21784 21292 21790 21304
rect 22462 21292 22468 21344
rect 22520 21332 22526 21344
rect 22646 21332 22652 21344
rect 22520 21304 22652 21332
rect 22520 21292 22526 21304
rect 22646 21292 22652 21304
rect 22704 21332 22710 21344
rect 22925 21335 22983 21341
rect 22925 21332 22937 21335
rect 22704 21304 22937 21332
rect 22704 21292 22710 21304
rect 22925 21301 22937 21304
rect 22971 21301 22983 21335
rect 22925 21295 22983 21301
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23658 21332 23664 21344
rect 23072 21304 23664 21332
rect 23072 21292 23078 21304
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 16114 21088 16120 21140
rect 16172 21128 16178 21140
rect 16209 21131 16267 21137
rect 16209 21128 16221 21131
rect 16172 21100 16221 21128
rect 16172 21088 16178 21100
rect 16209 21097 16221 21100
rect 16255 21097 16267 21131
rect 16209 21091 16267 21097
rect 16390 21088 16396 21140
rect 16448 21128 16454 21140
rect 16761 21131 16819 21137
rect 16761 21128 16773 21131
rect 16448 21100 16773 21128
rect 16448 21088 16454 21100
rect 16761 21097 16773 21100
rect 16807 21097 16819 21131
rect 19426 21128 19432 21140
rect 19387 21100 19432 21128
rect 16761 21091 16819 21097
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 20346 21088 20352 21140
rect 20404 21128 20410 21140
rect 20625 21131 20683 21137
rect 20625 21128 20637 21131
rect 20404 21100 20637 21128
rect 20404 21088 20410 21100
rect 20625 21097 20637 21100
rect 20671 21097 20683 21131
rect 20625 21091 20683 21097
rect 21637 21131 21695 21137
rect 21637 21097 21649 21131
rect 21683 21128 21695 21131
rect 21726 21128 21732 21140
rect 21683 21100 21732 21128
rect 21683 21097 21695 21100
rect 21637 21091 21695 21097
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 22738 21128 22744 21140
rect 22699 21100 22744 21128
rect 22738 21088 22744 21100
rect 22796 21088 22802 21140
rect 25498 21128 25504 21140
rect 25459 21100 25504 21128
rect 25498 21088 25504 21100
rect 25556 21088 25562 21140
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 14366 21060 14372 21072
rect 13872 21032 13917 21060
rect 14327 21032 14372 21060
rect 13872 21020 13878 21032
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 18871 21063 18929 21069
rect 18871 21029 18883 21063
rect 18917 21060 18929 21063
rect 19334 21060 19340 21072
rect 18917 21032 19340 21060
rect 18917 21029 18929 21032
rect 18871 21023 18929 21029
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 1118 20952 1124 21004
rect 1176 20992 1182 21004
rect 1432 20995 1490 21001
rect 1432 20992 1444 20995
rect 1176 20964 1444 20992
rect 1176 20952 1182 20964
rect 1432 20961 1444 20964
rect 1478 20961 1490 20995
rect 1432 20955 1490 20961
rect 10042 20952 10048 21004
rect 10100 20992 10106 21004
rect 11790 20992 11796 21004
rect 11848 21001 11854 21004
rect 11848 20995 11886 21001
rect 10100 20964 11796 20992
rect 10100 20952 10106 20964
rect 11790 20952 11796 20964
rect 11874 20961 11886 20995
rect 11848 20955 11886 20961
rect 11848 20952 11854 20955
rect 21082 20952 21088 21004
rect 21140 20992 21146 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 21140 20964 21281 20992
rect 21140 20952 21146 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 23934 20992 23940 21004
rect 23895 20964 23940 20992
rect 21269 20955 21327 20961
rect 23934 20952 23940 20964
rect 23992 20952 23998 21004
rect 25130 20952 25136 21004
rect 25188 20992 25194 21004
rect 25317 20995 25375 21001
rect 25317 20992 25329 20995
rect 25188 20964 25329 20992
rect 25188 20952 25194 20964
rect 25317 20961 25329 20964
rect 25363 20961 25375 20995
rect 25317 20955 25375 20961
rect 13725 20927 13783 20933
rect 13725 20893 13737 20927
rect 13771 20893 13783 20927
rect 13725 20887 13783 20893
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20924 15899 20927
rect 16574 20924 16580 20936
rect 15887 20896 16580 20924
rect 15887 20893 15899 20896
rect 15841 20887 15899 20893
rect 13740 20800 13768 20887
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18598 20924 18604 20936
rect 18555 20896 18604 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 18598 20884 18604 20896
rect 18656 20884 18662 20936
rect 24026 20884 24032 20936
rect 24084 20924 24090 20936
rect 27614 20924 27620 20936
rect 24084 20896 27620 20924
rect 24084 20884 24090 20896
rect 27614 20884 27620 20896
rect 27672 20884 27678 20936
rect 1535 20791 1593 20797
rect 1535 20757 1547 20791
rect 1581 20788 1593 20791
rect 3234 20788 3240 20800
rect 1581 20760 3240 20788
rect 1581 20757 1593 20760
rect 1535 20751 1593 20757
rect 3234 20748 3240 20760
rect 3292 20748 3298 20800
rect 11931 20791 11989 20797
rect 11931 20757 11943 20791
rect 11977 20788 11989 20791
rect 12805 20791 12863 20797
rect 12805 20788 12817 20791
rect 11977 20760 12817 20788
rect 11977 20757 11989 20760
rect 11931 20751 11989 20757
rect 12805 20757 12817 20760
rect 12851 20788 12863 20791
rect 12894 20788 12900 20800
rect 12851 20760 12900 20788
rect 12851 20757 12863 20760
rect 12805 20751 12863 20757
rect 12894 20748 12900 20760
rect 12952 20748 12958 20800
rect 13541 20791 13599 20797
rect 13541 20757 13553 20791
rect 13587 20788 13599 20791
rect 13722 20788 13728 20800
rect 13587 20760 13728 20788
rect 13587 20757 13599 20760
rect 13541 20751 13599 20757
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 18233 20791 18291 20797
rect 18233 20788 18245 20791
rect 17460 20760 18245 20788
rect 17460 20748 17466 20760
rect 18233 20757 18245 20760
rect 18279 20788 18291 20791
rect 18690 20788 18696 20800
rect 18279 20760 18696 20788
rect 18279 20757 18291 20760
rect 18233 20751 18291 20757
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19794 20788 19800 20800
rect 19755 20760 19800 20788
rect 19794 20748 19800 20760
rect 19852 20748 19858 20800
rect 24026 20788 24032 20800
rect 23987 20760 24032 20788
rect 24026 20748 24032 20760
rect 24084 20748 24090 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1118 20544 1124 20596
rect 1176 20584 1182 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 1176 20556 1593 20584
rect 1176 20544 1182 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 5534 20584 5540 20596
rect 5495 20556 5540 20584
rect 1581 20547 1639 20553
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 11790 20584 11796 20596
rect 11751 20556 11796 20584
rect 11790 20544 11796 20556
rect 11848 20544 11854 20596
rect 13814 20544 13820 20596
rect 13872 20584 13878 20596
rect 13909 20587 13967 20593
rect 13909 20584 13921 20587
rect 13872 20556 13921 20584
rect 13872 20544 13878 20556
rect 13909 20553 13921 20556
rect 13955 20584 13967 20587
rect 15286 20584 15292 20596
rect 13955 20556 15292 20584
rect 13955 20553 13967 20556
rect 13909 20547 13967 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 17126 20584 17132 20596
rect 17087 20556 17132 20584
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 20717 20587 20775 20593
rect 20717 20553 20729 20587
rect 20763 20584 20775 20587
rect 21082 20584 21088 20596
rect 20763 20556 21088 20584
rect 20763 20553 20775 20556
rect 20717 20547 20775 20553
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 22462 20584 22468 20596
rect 22423 20556 22468 20584
rect 22462 20544 22468 20556
rect 22520 20544 22526 20596
rect 24026 20584 24032 20596
rect 23987 20556 24032 20584
rect 24026 20544 24032 20556
rect 24084 20544 24090 20596
rect 14277 20519 14335 20525
rect 14277 20485 14289 20519
rect 14323 20516 14335 20519
rect 15749 20519 15807 20525
rect 15749 20516 15761 20519
rect 14323 20488 15761 20516
rect 14323 20485 14335 20488
rect 14277 20479 14335 20485
rect 12894 20448 12900 20460
rect 12855 20420 12900 20448
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 5144 20383 5202 20389
rect 5144 20349 5156 20383
rect 5190 20380 5202 20383
rect 5534 20380 5540 20392
rect 5190 20352 5540 20380
rect 5190 20349 5202 20352
rect 5144 20343 5202 20349
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 14366 20380 14372 20392
rect 14327 20352 14372 20380
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 12713 20315 12771 20321
rect 12713 20281 12725 20315
rect 12759 20312 12771 20315
rect 12986 20312 12992 20324
rect 12759 20284 12992 20312
rect 12759 20281 12771 20284
rect 12713 20275 12771 20281
rect 12986 20272 12992 20284
rect 13044 20272 13050 20324
rect 13541 20315 13599 20321
rect 13541 20281 13553 20315
rect 13587 20312 13599 20315
rect 13722 20312 13728 20324
rect 13587 20284 13728 20312
rect 13587 20281 13599 20284
rect 13541 20275 13599 20281
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 14705 20321 14733 20488
rect 15749 20485 15761 20488
rect 15795 20516 15807 20519
rect 16114 20516 16120 20528
rect 15795 20488 16120 20516
rect 15795 20485 15807 20488
rect 15749 20479 15807 20485
rect 16114 20476 16120 20488
rect 16172 20516 16178 20528
rect 16482 20516 16488 20528
rect 16172 20488 16488 20516
rect 16172 20476 16178 20488
rect 16482 20476 16488 20488
rect 16540 20516 16546 20528
rect 19334 20516 19340 20528
rect 16540 20488 19340 20516
rect 16540 20476 16546 20488
rect 19334 20476 19340 20488
rect 19392 20476 19398 20528
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20448 19027 20451
rect 19794 20448 19800 20460
rect 19015 20420 19800 20448
rect 19015 20417 19027 20420
rect 18969 20411 19027 20417
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 23477 20451 23535 20457
rect 23477 20417 23489 20451
rect 23523 20448 23535 20451
rect 24213 20451 24271 20457
rect 24213 20448 24225 20451
rect 23523 20420 24225 20448
rect 23523 20417 23535 20420
rect 23477 20411 23535 20417
rect 24213 20417 24225 20420
rect 24259 20448 24271 20451
rect 25314 20448 25320 20460
rect 24259 20420 25320 20448
rect 24259 20417 24271 20420
rect 24213 20411 24271 20417
rect 25314 20408 25320 20420
rect 25372 20408 25378 20460
rect 16114 20340 16120 20392
rect 16172 20380 16178 20392
rect 16209 20383 16267 20389
rect 16209 20380 16221 20383
rect 16172 20352 16221 20380
rect 16172 20340 16178 20352
rect 16209 20349 16221 20352
rect 16255 20380 16267 20383
rect 17405 20383 17463 20389
rect 17405 20380 17417 20383
rect 16255 20352 17417 20380
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 17405 20349 17417 20352
rect 17451 20349 17463 20383
rect 18233 20383 18291 20389
rect 18233 20380 18245 20383
rect 17405 20343 17463 20349
rect 17880 20352 18245 20380
rect 14690 20315 14748 20321
rect 14690 20281 14702 20315
rect 14736 20281 14748 20315
rect 14690 20275 14748 20281
rect 5215 20247 5273 20253
rect 5215 20213 5227 20247
rect 5261 20244 5273 20247
rect 9674 20244 9680 20256
rect 5261 20216 9680 20244
rect 5261 20213 5273 20216
rect 5215 20207 5273 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 12894 20204 12900 20256
rect 12952 20244 12958 20256
rect 14705 20244 14733 20275
rect 17880 20256 17908 20352
rect 18233 20349 18245 20352
rect 18279 20349 18291 20383
rect 18690 20380 18696 20392
rect 18651 20352 18696 20380
rect 18233 20343 18291 20349
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 21542 20380 21548 20392
rect 21503 20352 21548 20380
rect 21542 20340 21548 20352
rect 21600 20340 21606 20392
rect 20159 20315 20217 20321
rect 20159 20281 20171 20315
rect 20205 20281 20217 20315
rect 21866 20315 21924 20321
rect 21866 20312 21878 20315
rect 20159 20275 20217 20281
rect 21376 20284 21878 20312
rect 12952 20216 14733 20244
rect 12952 20204 12958 20216
rect 16482 20204 16488 20256
rect 16540 20244 16546 20256
rect 16577 20247 16635 20253
rect 16577 20244 16589 20247
rect 16540 20216 16589 20244
rect 16540 20204 16546 20216
rect 16577 20213 16589 20216
rect 16623 20213 16635 20247
rect 17862 20244 17868 20256
rect 17823 20216 17868 20244
rect 16577 20207 16635 20213
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 19334 20244 19340 20256
rect 19295 20216 19340 20244
rect 19334 20204 19340 20216
rect 19392 20244 19398 20256
rect 19613 20247 19671 20253
rect 19613 20244 19625 20247
rect 19392 20216 19625 20244
rect 19392 20204 19398 20216
rect 19613 20213 19625 20216
rect 19659 20244 19671 20247
rect 20174 20244 20202 20275
rect 21376 20253 21404 20284
rect 21866 20281 21878 20284
rect 21912 20281 21924 20315
rect 23934 20312 23940 20324
rect 21866 20275 21924 20281
rect 23446 20284 23940 20312
rect 21361 20247 21419 20253
rect 21361 20244 21373 20247
rect 19659 20216 21373 20244
rect 19659 20213 19671 20216
rect 19613 20207 19671 20213
rect 21361 20213 21373 20216
rect 21407 20213 21419 20247
rect 21361 20207 21419 20213
rect 23109 20247 23167 20253
rect 23109 20213 23121 20247
rect 23155 20244 23167 20247
rect 23290 20244 23296 20256
rect 23155 20216 23296 20244
rect 23155 20213 23167 20216
rect 23109 20207 23167 20213
rect 23290 20204 23296 20216
rect 23348 20244 23354 20256
rect 23446 20244 23474 20284
rect 23934 20272 23940 20284
rect 23992 20272 23998 20324
rect 24305 20315 24363 20321
rect 24305 20281 24317 20315
rect 24351 20281 24363 20315
rect 24305 20275 24363 20281
rect 23348 20216 23474 20244
rect 23348 20204 23354 20216
rect 24026 20204 24032 20256
rect 24084 20244 24090 20256
rect 24320 20244 24348 20275
rect 24486 20272 24492 20324
rect 24544 20312 24550 20324
rect 24857 20315 24915 20321
rect 24857 20312 24869 20315
rect 24544 20284 24869 20312
rect 24544 20272 24550 20284
rect 24857 20281 24869 20284
rect 24903 20281 24915 20315
rect 24857 20275 24915 20281
rect 24084 20216 24348 20244
rect 24084 20204 24090 20216
rect 25130 20204 25136 20256
rect 25188 20244 25194 20256
rect 25317 20247 25375 20253
rect 25317 20244 25329 20247
rect 25188 20216 25329 20244
rect 25188 20204 25194 20216
rect 25317 20213 25329 20216
rect 25363 20213 25375 20247
rect 25317 20207 25375 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 14461 20043 14519 20049
rect 14461 20040 14473 20043
rect 14424 20012 14473 20040
rect 14424 20000 14430 20012
rect 14461 20009 14473 20012
rect 14507 20040 14519 20043
rect 15381 20043 15439 20049
rect 15381 20040 15393 20043
rect 14507 20012 15393 20040
rect 14507 20009 14519 20012
rect 14461 20003 14519 20009
rect 15381 20009 15393 20012
rect 15427 20009 15439 20043
rect 15381 20003 15439 20009
rect 21315 20043 21373 20049
rect 21315 20009 21327 20043
rect 21361 20040 21373 20043
rect 25130 20040 25136 20052
rect 21361 20012 25136 20040
rect 21361 20009 21373 20012
rect 21315 20003 21373 20009
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 25314 20040 25320 20052
rect 25275 20012 25320 20040
rect 25314 20000 25320 20012
rect 25372 20000 25378 20052
rect 18046 19972 18052 19984
rect 18007 19944 18052 19972
rect 18046 19932 18052 19944
rect 18104 19932 18110 19984
rect 18690 19932 18696 19984
rect 18748 19972 18754 19984
rect 19613 19975 19671 19981
rect 18748 19944 19380 19972
rect 18748 19932 18754 19944
rect 12986 19864 12992 19916
rect 13044 19904 13050 19916
rect 13170 19904 13176 19916
rect 13044 19876 13176 19904
rect 13044 19864 13050 19876
rect 13170 19864 13176 19876
rect 13228 19904 13234 19916
rect 13265 19907 13323 19913
rect 13265 19904 13277 19907
rect 13228 19876 13277 19904
rect 13228 19864 13234 19876
rect 13265 19873 13277 19876
rect 13311 19873 13323 19907
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 13265 19867 13323 19873
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19873 15807 19907
rect 15749 19867 15807 19873
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19836 15163 19839
rect 15764 19836 15792 19867
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 15896 19876 16129 19904
rect 15896 19864 15902 19876
rect 16117 19873 16129 19876
rect 16163 19904 16175 19907
rect 17313 19907 17371 19913
rect 17313 19904 17325 19907
rect 16163 19876 17325 19904
rect 16163 19873 16175 19876
rect 16117 19867 16175 19873
rect 17313 19873 17325 19876
rect 17359 19873 17371 19907
rect 17770 19904 17776 19916
rect 17731 19876 17776 19904
rect 17313 19867 17371 19873
rect 15930 19836 15936 19848
rect 15151 19808 15936 19836
rect 15151 19805 15163 19808
rect 15105 19799 15163 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 17328 19836 17356 19867
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 19352 19913 19380 19944
rect 19613 19941 19625 19975
rect 19659 19972 19671 19975
rect 21542 19972 21548 19984
rect 19659 19944 21548 19972
rect 19659 19941 19671 19944
rect 19613 19935 19671 19941
rect 21542 19932 21548 19944
rect 21600 19972 21606 19984
rect 21637 19975 21695 19981
rect 21637 19972 21649 19975
rect 21600 19944 21649 19972
rect 21600 19932 21606 19944
rect 21637 19941 21649 19944
rect 21683 19941 21695 19975
rect 22370 19972 22376 19984
rect 22331 19944 22376 19972
rect 21637 19935 21695 19941
rect 22370 19932 22376 19944
rect 22428 19932 22434 19984
rect 23934 19972 23940 19984
rect 23895 19944 23940 19972
rect 23934 19932 23940 19944
rect 23992 19932 23998 19984
rect 24486 19972 24492 19984
rect 24447 19944 24492 19972
rect 24486 19932 24492 19944
rect 24544 19932 24550 19984
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 19337 19907 19395 19913
rect 19337 19873 19349 19907
rect 19383 19904 19395 19907
rect 20070 19904 20076 19916
rect 19383 19876 20076 19904
rect 19383 19873 19395 19876
rect 19337 19867 19395 19873
rect 18892 19836 18920 19867
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 21244 19907 21302 19913
rect 21244 19873 21256 19907
rect 21290 19904 21302 19907
rect 21910 19904 21916 19916
rect 21290 19876 21916 19904
rect 21290 19873 21302 19876
rect 21244 19867 21302 19873
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 22278 19836 22284 19848
rect 17328 19808 18920 19836
rect 22239 19808 22284 19836
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 22925 19839 22983 19845
rect 22925 19805 22937 19839
rect 22971 19836 22983 19839
rect 23845 19839 23903 19845
rect 23845 19836 23857 19839
rect 22971 19808 23857 19836
rect 22971 19805 22983 19808
rect 22925 19799 22983 19805
rect 23845 19805 23857 19808
rect 23891 19836 23903 19839
rect 24026 19836 24032 19848
rect 23891 19808 24032 19836
rect 23891 19805 23903 19808
rect 23845 19799 23903 19805
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 23106 19728 23112 19780
rect 23164 19768 23170 19780
rect 23658 19768 23664 19780
rect 23164 19740 23664 19768
rect 23164 19728 23170 19740
rect 23658 19728 23664 19740
rect 23716 19728 23722 19780
rect 24486 19768 24492 19780
rect 23860 19740 24492 19768
rect 12986 19700 12992 19712
rect 12947 19672 12992 19700
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 13630 19700 13636 19712
rect 13591 19672 13636 19700
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 16669 19703 16727 19709
rect 16669 19700 16681 19703
rect 16632 19672 16681 19700
rect 16632 19660 16638 19672
rect 16669 19669 16681 19672
rect 16715 19669 16727 19703
rect 16669 19663 16727 19669
rect 18417 19703 18475 19709
rect 18417 19669 18429 19703
rect 18463 19700 18475 19703
rect 18598 19700 18604 19712
rect 18463 19672 18604 19700
rect 18463 19669 18475 19672
rect 18417 19663 18475 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 18785 19703 18843 19709
rect 18785 19669 18797 19703
rect 18831 19700 18843 19703
rect 19150 19700 19156 19712
rect 18831 19672 19156 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 23198 19700 23204 19712
rect 23159 19672 23204 19700
rect 23198 19660 23204 19672
rect 23256 19700 23262 19712
rect 23860 19700 23888 19740
rect 24486 19728 24492 19740
rect 24544 19728 24550 19780
rect 23256 19672 23888 19700
rect 23256 19660 23262 19672
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 16574 19456 16580 19508
rect 16632 19496 16638 19508
rect 20070 19496 20076 19508
rect 16632 19468 16677 19496
rect 20031 19468 20076 19496
rect 16632 19456 16638 19468
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 25406 19496 25412 19508
rect 25367 19468 25412 19496
rect 25406 19456 25412 19468
rect 25464 19456 25470 19508
rect 22695 19431 22753 19437
rect 22695 19397 22707 19431
rect 22741 19428 22753 19431
rect 24210 19428 24216 19440
rect 22741 19400 24216 19428
rect 22741 19397 22753 19400
rect 22695 19391 22753 19397
rect 24210 19388 24216 19400
rect 24268 19388 24274 19440
rect 14645 19363 14703 19369
rect 14645 19329 14657 19363
rect 14691 19360 14703 19363
rect 14691 19332 16344 19360
rect 14691 19329 14703 19332
rect 14645 19323 14703 19329
rect 12986 19292 12992 19304
rect 12947 19264 12992 19292
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 15562 19292 15568 19304
rect 15523 19264 15568 19292
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 15930 19292 15936 19304
rect 15891 19264 15936 19292
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 16316 19301 16344 19332
rect 22278 19320 22284 19372
rect 22336 19360 22342 19372
rect 23017 19363 23075 19369
rect 23017 19360 23029 19363
rect 22336 19332 23029 19360
rect 22336 19320 22342 19332
rect 23017 19329 23029 19332
rect 23063 19329 23075 19363
rect 24026 19360 24032 19372
rect 23987 19332 24032 19360
rect 23017 19323 23075 19329
rect 24026 19320 24032 19332
rect 24084 19360 24090 19372
rect 24673 19363 24731 19369
rect 24673 19360 24685 19363
rect 24084 19332 24685 19360
rect 24084 19320 24090 19332
rect 24673 19329 24685 19332
rect 24719 19329 24731 19363
rect 24673 19323 24731 19329
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19292 16359 19295
rect 17770 19292 17776 19304
rect 16347 19264 17356 19292
rect 17683 19264 17776 19292
rect 16347 19261 16359 19264
rect 16301 19255 16359 19261
rect 12618 19184 12624 19236
rect 12676 19224 12682 19236
rect 12894 19224 12900 19236
rect 12676 19196 12900 19224
rect 12676 19184 12682 19196
rect 12894 19184 12900 19196
rect 12952 19224 12958 19236
rect 13310 19227 13368 19233
rect 13310 19224 13322 19227
rect 12952 19196 13322 19224
rect 12952 19184 12958 19196
rect 13310 19193 13322 19196
rect 13356 19193 13368 19227
rect 13310 19187 13368 19193
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 15286 19224 15292 19236
rect 14884 19196 15292 19224
rect 14884 19184 14890 19196
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 15948 19224 15976 19252
rect 16853 19227 16911 19233
rect 16853 19224 16865 19227
rect 15948 19196 16865 19224
rect 16853 19193 16865 19196
rect 16899 19193 16911 19227
rect 17328 19224 17356 19264
rect 17770 19252 17776 19264
rect 17828 19292 17834 19304
rect 18506 19292 18512 19304
rect 17828 19264 18512 19292
rect 17828 19252 17834 19264
rect 18506 19252 18512 19264
rect 18564 19252 18570 19304
rect 18693 19295 18751 19301
rect 18693 19261 18705 19295
rect 18739 19261 18751 19295
rect 19150 19292 19156 19304
rect 19111 19264 19156 19292
rect 18693 19255 18751 19261
rect 17862 19224 17868 19236
rect 17328 19196 17868 19224
rect 16853 19187 16911 19193
rect 17862 19184 17868 19196
rect 17920 19224 17926 19236
rect 18708 19224 18736 19255
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19429 19295 19487 19301
rect 19429 19261 19441 19295
rect 19475 19292 19487 19295
rect 20622 19292 20628 19304
rect 19475 19264 20628 19292
rect 19475 19261 19487 19264
rect 19429 19255 19487 19261
rect 20622 19252 20628 19264
rect 20680 19292 20686 19304
rect 20809 19295 20867 19301
rect 20809 19292 20821 19295
rect 20680 19264 20821 19292
rect 20680 19252 20686 19264
rect 20809 19261 20821 19264
rect 20855 19261 20867 19295
rect 20809 19255 20867 19261
rect 22624 19295 22682 19301
rect 22624 19261 22636 19295
rect 22670 19292 22682 19295
rect 23198 19292 23204 19304
rect 22670 19264 23204 19292
rect 22670 19261 22682 19264
rect 22624 19255 22682 19261
rect 23198 19252 23204 19264
rect 23256 19252 23262 19304
rect 25222 19292 25228 19304
rect 25183 19264 25228 19292
rect 25222 19252 25228 19264
rect 25280 19292 25286 19304
rect 25777 19295 25835 19301
rect 25777 19292 25789 19295
rect 25280 19264 25789 19292
rect 25280 19252 25286 19264
rect 25777 19261 25789 19264
rect 25823 19261 25835 19295
rect 25777 19255 25835 19261
rect 17920 19196 18092 19224
rect 17920 19184 17926 19196
rect 18064 19168 18092 19196
rect 18524 19196 18736 19224
rect 13170 19116 13176 19168
rect 13228 19156 13234 19168
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 13228 19128 13921 19156
rect 13228 19116 13234 19128
rect 13909 19125 13921 19128
rect 13955 19125 13967 19159
rect 13909 19119 13967 19125
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19156 15071 19159
rect 15838 19156 15844 19168
rect 15059 19128 15844 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15838 19116 15844 19128
rect 15896 19156 15902 19168
rect 17313 19159 17371 19165
rect 17313 19156 17325 19159
rect 15896 19128 17325 19156
rect 15896 19116 15902 19128
rect 17313 19125 17325 19128
rect 17359 19125 17371 19159
rect 17313 19119 17371 19125
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 18524 19165 18552 19196
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 20717 19227 20775 19233
rect 20717 19224 20729 19227
rect 19392 19196 20729 19224
rect 19392 19184 19398 19196
rect 20717 19193 20729 19196
rect 20763 19224 20775 19227
rect 21171 19227 21229 19233
rect 21171 19224 21183 19227
rect 20763 19196 21183 19224
rect 20763 19193 20775 19196
rect 20717 19187 20775 19193
rect 21171 19193 21183 19196
rect 21217 19224 21229 19227
rect 22094 19224 22100 19236
rect 21217 19196 22100 19224
rect 21217 19193 21229 19196
rect 21171 19187 21229 19193
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 23750 19224 23756 19236
rect 23711 19196 23756 19224
rect 23750 19184 23756 19196
rect 23808 19184 23814 19236
rect 23845 19227 23903 19233
rect 23845 19193 23857 19227
rect 23891 19193 23903 19227
rect 23845 19187 23903 19193
rect 18509 19159 18567 19165
rect 18509 19156 18521 19159
rect 18104 19128 18521 19156
rect 18104 19116 18110 19128
rect 18509 19125 18521 19128
rect 18555 19125 18567 19159
rect 18509 19119 18567 19125
rect 18690 19116 18696 19168
rect 18748 19156 18754 19168
rect 19705 19159 19763 19165
rect 19705 19156 19717 19159
rect 18748 19128 19717 19156
rect 18748 19116 18754 19128
rect 19705 19125 19717 19128
rect 19751 19125 19763 19159
rect 19705 19119 19763 19125
rect 20990 19116 20996 19168
rect 21048 19156 21054 19168
rect 21729 19159 21787 19165
rect 21729 19156 21741 19159
rect 21048 19128 21741 19156
rect 21048 19116 21054 19128
rect 21729 19125 21741 19128
rect 21775 19156 21787 19159
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21775 19128 22201 19156
rect 21775 19125 21787 19128
rect 21729 19119 21787 19125
rect 22189 19125 22201 19128
rect 22235 19156 22247 19159
rect 22370 19156 22376 19168
rect 22235 19128 22376 19156
rect 22235 19125 22247 19128
rect 22189 19119 22247 19125
rect 22370 19116 22376 19128
rect 22428 19116 22434 19168
rect 23382 19156 23388 19168
rect 23343 19128 23388 19156
rect 23382 19116 23388 19128
rect 23440 19156 23446 19168
rect 23860 19156 23888 19187
rect 23440 19128 23888 19156
rect 23440 19116 23446 19128
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 13170 18952 13176 18964
rect 13131 18924 13176 18952
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 15105 18955 15163 18961
rect 15105 18921 15117 18955
rect 15151 18952 15163 18955
rect 15930 18952 15936 18964
rect 15151 18924 15936 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 16114 18952 16120 18964
rect 16075 18924 16120 18952
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 20622 18952 20628 18964
rect 20583 18924 20628 18952
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 21910 18952 21916 18964
rect 21871 18924 21916 18952
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 23290 18912 23296 18964
rect 23348 18952 23354 18964
rect 23385 18955 23443 18961
rect 23385 18952 23397 18955
rect 23348 18924 23397 18952
rect 23348 18912 23354 18924
rect 23385 18921 23397 18924
rect 23431 18952 23443 18955
rect 23753 18955 23811 18961
rect 23753 18952 23765 18955
rect 23431 18924 23765 18952
rect 23431 18921 23443 18924
rect 23385 18915 23443 18921
rect 23753 18921 23765 18924
rect 23799 18921 23811 18955
rect 23753 18915 23811 18921
rect 24765 18955 24823 18961
rect 24765 18921 24777 18955
rect 24811 18952 24823 18955
rect 24854 18952 24860 18964
rect 24811 18924 24860 18952
rect 24811 18921 24823 18924
rect 24765 18915 24823 18921
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 13630 18844 13636 18896
rect 13688 18884 13694 18896
rect 13725 18887 13783 18893
rect 13725 18884 13737 18887
rect 13688 18856 13737 18884
rect 13688 18844 13694 18856
rect 13725 18853 13737 18856
rect 13771 18853 13783 18887
rect 13725 18847 13783 18853
rect 15562 18776 15568 18828
rect 15620 18816 15626 18828
rect 15841 18819 15899 18825
rect 15841 18816 15853 18819
rect 15620 18788 15853 18816
rect 15620 18776 15626 18788
rect 15841 18785 15853 18788
rect 15887 18785 15899 18819
rect 15948 18816 15976 18912
rect 22278 18844 22284 18896
rect 22336 18884 22342 18896
rect 22786 18887 22844 18893
rect 22786 18884 22798 18887
rect 22336 18856 22798 18884
rect 22336 18844 22342 18856
rect 22786 18853 22798 18856
rect 22832 18853 22844 18887
rect 22786 18847 22844 18853
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15948 18788 16313 18816
rect 15841 18779 15899 18785
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18816 16727 18819
rect 18690 18816 18696 18828
rect 16715 18788 18696 18816
rect 16715 18785 16727 18788
rect 16669 18779 16727 18785
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 13648 18612 13676 18711
rect 13722 18708 13728 18760
rect 13780 18748 13786 18760
rect 13909 18751 13967 18757
rect 13909 18748 13921 18751
rect 13780 18720 13921 18748
rect 13780 18708 13786 18720
rect 13909 18717 13921 18720
rect 13955 18717 13967 18751
rect 16684 18748 16712 18779
rect 18690 18776 18696 18788
rect 18748 18776 18754 18828
rect 19150 18816 19156 18828
rect 19111 18788 19156 18816
rect 19150 18776 19156 18788
rect 19208 18776 19214 18828
rect 20990 18816 20996 18828
rect 20951 18788 20996 18816
rect 20990 18776 20996 18788
rect 21048 18776 21054 18828
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 23382 18816 23388 18828
rect 21683 18788 23388 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 23382 18776 23388 18788
rect 23440 18776 23446 18828
rect 24210 18776 24216 18828
rect 24268 18816 24274 18828
rect 24581 18819 24639 18825
rect 24581 18816 24593 18819
rect 24268 18788 24593 18816
rect 24268 18776 24274 18788
rect 24581 18785 24593 18788
rect 24627 18785 24639 18819
rect 24581 18779 24639 18785
rect 13909 18711 13967 18717
rect 16218 18720 16712 18748
rect 19429 18751 19487 18757
rect 15838 18640 15844 18692
rect 15896 18680 15902 18692
rect 16218 18680 16246 18720
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 22465 18751 22523 18757
rect 22465 18748 22477 18751
rect 19475 18720 22477 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 22465 18717 22477 18720
rect 22511 18748 22523 18751
rect 22830 18748 22836 18760
rect 22511 18720 22836 18748
rect 22511 18717 22523 18720
rect 22465 18711 22523 18717
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 15896 18652 16246 18680
rect 15896 18640 15902 18652
rect 13998 18612 14004 18624
rect 13648 18584 14004 18612
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 15562 18612 15568 18624
rect 15523 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 23750 18572 23756 18624
rect 23808 18612 23814 18624
rect 24213 18615 24271 18621
rect 24213 18612 24225 18615
rect 23808 18584 24225 18612
rect 23808 18572 23814 18584
rect 24213 18581 24225 18584
rect 24259 18612 24271 18615
rect 25038 18612 25044 18624
rect 24259 18584 25044 18612
rect 24259 18581 24271 18584
rect 24213 18575 24271 18581
rect 25038 18572 25044 18584
rect 25096 18572 25102 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 3786 18368 3792 18420
rect 3844 18408 3850 18420
rect 3973 18411 4031 18417
rect 3973 18408 3985 18411
rect 3844 18380 3985 18408
rect 3844 18368 3850 18380
rect 3973 18377 3985 18380
rect 4019 18377 4031 18411
rect 13630 18408 13636 18420
rect 13591 18380 13636 18408
rect 3973 18371 4031 18377
rect 13630 18368 13636 18380
rect 13688 18368 13694 18420
rect 18690 18368 18696 18420
rect 18748 18408 18754 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 18748 18380 19073 18408
rect 18748 18368 18754 18380
rect 19061 18377 19073 18380
rect 19107 18377 19119 18411
rect 19061 18371 19119 18377
rect 20073 18411 20131 18417
rect 20073 18377 20085 18411
rect 20119 18408 20131 18411
rect 20990 18408 20996 18420
rect 20119 18380 20996 18408
rect 20119 18377 20131 18380
rect 20073 18371 20131 18377
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 22830 18408 22836 18420
rect 22791 18380 22836 18408
rect 22830 18368 22836 18380
rect 22888 18368 22894 18420
rect 24762 18408 24768 18420
rect 24723 18380 24768 18408
rect 24762 18368 24768 18380
rect 24820 18368 24826 18420
rect 17129 18343 17187 18349
rect 17129 18309 17141 18343
rect 17175 18309 17187 18343
rect 17129 18303 17187 18309
rect 15930 18272 15936 18284
rect 15891 18244 15936 18272
rect 15930 18232 15936 18244
rect 15988 18272 15994 18284
rect 16761 18275 16819 18281
rect 16761 18272 16773 18275
rect 15988 18244 16773 18272
rect 15988 18232 15994 18244
rect 16761 18241 16773 18244
rect 16807 18272 16819 18275
rect 17144 18272 17172 18303
rect 18598 18272 18604 18284
rect 16807 18244 17172 18272
rect 18559 18244 18604 18272
rect 16807 18241 16819 18244
rect 16761 18235 16819 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 21910 18272 21916 18284
rect 21871 18244 21916 18272
rect 21910 18232 21916 18244
rect 21968 18232 21974 18284
rect 3580 18207 3638 18213
rect 3580 18173 3592 18207
rect 3626 18204 3638 18207
rect 3786 18204 3792 18216
rect 3626 18176 3792 18204
rect 3626 18173 3638 18176
rect 3580 18167 3638 18173
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15013 18207 15071 18213
rect 15013 18204 15025 18207
rect 14884 18176 15025 18204
rect 14884 18164 14890 18176
rect 15013 18173 15025 18176
rect 15059 18173 15071 18207
rect 15013 18167 15071 18173
rect 15841 18207 15899 18213
rect 15841 18173 15853 18207
rect 15887 18173 15899 18207
rect 15841 18167 15899 18173
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18204 17003 18207
rect 17034 18204 17040 18216
rect 16991 18176 17040 18204
rect 16991 18173 17003 18176
rect 16945 18167 17003 18173
rect 12986 18096 12992 18148
rect 13044 18136 13050 18148
rect 13044 18108 15010 18136
rect 13044 18096 13050 18108
rect 3651 18071 3709 18077
rect 3651 18037 3663 18071
rect 3697 18068 3709 18071
rect 3878 18068 3884 18080
rect 3697 18040 3884 18068
rect 3697 18037 3709 18040
rect 3651 18031 3709 18037
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 13998 18068 14004 18080
rect 13959 18040 14004 18068
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 14826 18068 14832 18080
rect 14787 18040 14832 18068
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 14982 18068 15010 18108
rect 15194 18096 15200 18148
rect 15252 18136 15258 18148
rect 15856 18136 15884 18167
rect 17034 18164 17040 18176
rect 17092 18204 17098 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 17092 18176 17417 18204
rect 17092 18164 17098 18176
rect 17405 18173 17417 18176
rect 17451 18173 17463 18207
rect 18046 18204 18052 18216
rect 17405 18167 17463 18173
rect 17788 18176 18052 18204
rect 17788 18136 17816 18176
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 18506 18204 18512 18216
rect 18467 18176 18512 18204
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 24581 18207 24639 18213
rect 24581 18173 24593 18207
rect 24627 18204 24639 18207
rect 24627 18176 24900 18204
rect 24627 18173 24639 18176
rect 24581 18167 24639 18173
rect 15252 18108 17816 18136
rect 15252 18096 15258 18108
rect 17788 18080 17816 18108
rect 18782 18096 18788 18148
rect 18840 18136 18846 18148
rect 19150 18136 19156 18148
rect 18840 18108 19156 18136
rect 18840 18096 18846 18108
rect 19150 18096 19156 18108
rect 19208 18136 19214 18148
rect 19429 18139 19487 18145
rect 19429 18136 19441 18139
rect 19208 18108 19441 18136
rect 19208 18096 19214 18108
rect 19429 18105 19441 18108
rect 19475 18105 19487 18139
rect 19429 18099 19487 18105
rect 20165 18139 20223 18145
rect 20165 18105 20177 18139
rect 20211 18136 20223 18139
rect 20717 18139 20775 18145
rect 20717 18136 20729 18139
rect 20211 18108 20729 18136
rect 20211 18105 20223 18108
rect 20165 18099 20223 18105
rect 20717 18105 20729 18108
rect 20763 18136 20775 18139
rect 21269 18139 21327 18145
rect 21269 18136 21281 18139
rect 20763 18108 21281 18136
rect 20763 18105 20775 18108
rect 20717 18099 20775 18105
rect 21269 18105 21281 18108
rect 21315 18105 21327 18139
rect 21269 18099 21327 18105
rect 21361 18139 21419 18145
rect 21361 18105 21373 18139
rect 21407 18136 21419 18139
rect 22002 18136 22008 18148
rect 21407 18108 22008 18136
rect 21407 18105 21419 18108
rect 21361 18099 21419 18105
rect 15105 18071 15163 18077
rect 15105 18068 15117 18071
rect 14982 18040 15117 18068
rect 15105 18037 15117 18040
rect 15151 18037 15163 18071
rect 15105 18031 15163 18037
rect 15562 18028 15568 18080
rect 15620 18068 15626 18080
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 15620 18040 16405 18068
rect 15620 18028 15626 18040
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 17770 18068 17776 18080
rect 17731 18040 17776 18068
rect 16393 18031 16451 18037
rect 17770 18028 17776 18040
rect 17828 18028 17834 18080
rect 21085 18071 21143 18077
rect 21085 18037 21097 18071
rect 21131 18068 21143 18071
rect 21376 18068 21404 18099
rect 22002 18096 22008 18108
rect 22060 18096 22066 18148
rect 24872 18080 24900 18176
rect 21131 18040 21404 18068
rect 21131 18037 21143 18040
rect 21085 18031 21143 18037
rect 22278 18028 22284 18080
rect 22336 18068 22342 18080
rect 22465 18071 22523 18077
rect 22465 18068 22477 18071
rect 22336 18040 22477 18068
rect 22336 18028 22342 18040
rect 22465 18037 22477 18040
rect 22511 18037 22523 18071
rect 22465 18031 22523 18037
rect 24210 18028 24216 18080
rect 24268 18068 24274 18080
rect 24397 18071 24455 18077
rect 24397 18068 24409 18071
rect 24268 18040 24409 18068
rect 24268 18028 24274 18040
rect 24397 18037 24409 18040
rect 24443 18037 24455 18071
rect 24397 18031 24455 18037
rect 24854 18028 24860 18080
rect 24912 18068 24918 18080
rect 25133 18071 25191 18077
rect 25133 18068 25145 18071
rect 24912 18040 25145 18068
rect 24912 18028 24918 18040
rect 25133 18037 25145 18040
rect 25179 18037 25191 18071
rect 25133 18031 25191 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 13998 17824 14004 17876
rect 14056 17864 14062 17876
rect 18923 17867 18981 17873
rect 18923 17864 18935 17867
rect 14056 17836 18935 17864
rect 14056 17824 14062 17836
rect 18923 17833 18935 17836
rect 18969 17833 18981 17867
rect 18923 17827 18981 17833
rect 21100 17836 22600 17864
rect 15105 17799 15163 17805
rect 15105 17765 15117 17799
rect 15151 17796 15163 17799
rect 15194 17796 15200 17808
rect 15151 17768 15200 17796
rect 15151 17765 15163 17768
rect 15105 17759 15163 17765
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 20714 17756 20720 17808
rect 20772 17796 20778 17808
rect 21100 17805 21128 17836
rect 21085 17799 21143 17805
rect 21085 17796 21097 17799
rect 20772 17768 21097 17796
rect 20772 17756 20778 17768
rect 21085 17765 21097 17768
rect 21131 17765 21143 17799
rect 21085 17759 21143 17765
rect 21637 17799 21695 17805
rect 21637 17765 21649 17799
rect 21683 17796 21695 17799
rect 21910 17796 21916 17808
rect 21683 17768 21916 17796
rect 21683 17765 21695 17768
rect 21637 17759 21695 17765
rect 21910 17756 21916 17768
rect 21968 17756 21974 17808
rect 22002 17756 22008 17808
rect 22060 17796 22066 17808
rect 22465 17799 22523 17805
rect 22465 17796 22477 17799
rect 22060 17768 22477 17796
rect 22060 17756 22066 17768
rect 22465 17765 22477 17768
rect 22511 17765 22523 17799
rect 22465 17759 22523 17765
rect 22572 17740 22600 17836
rect 1118 17688 1124 17740
rect 1176 17728 1182 17740
rect 1432 17731 1490 17737
rect 1432 17728 1444 17731
rect 1176 17700 1444 17728
rect 1176 17688 1182 17700
rect 1432 17697 1444 17700
rect 1478 17697 1490 17731
rect 16114 17728 16120 17740
rect 16075 17700 16120 17728
rect 1432 17691 1490 17697
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 18874 17728 18880 17740
rect 18831 17700 18880 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 18874 17688 18880 17700
rect 18932 17688 18938 17740
rect 19864 17731 19922 17737
rect 19864 17697 19876 17731
rect 19910 17728 19922 17731
rect 19978 17728 19984 17740
rect 19910 17700 19984 17728
rect 19910 17697 19922 17700
rect 19864 17691 19922 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 22554 17728 22560 17740
rect 22515 17700 22560 17728
rect 22554 17688 22560 17700
rect 22612 17688 22618 17740
rect 24673 17731 24731 17737
rect 24673 17697 24685 17731
rect 24719 17728 24731 17731
rect 24946 17728 24952 17740
rect 24719 17700 24952 17728
rect 24719 17697 24731 17700
rect 24673 17691 24731 17697
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 17586 17660 17592 17672
rect 17547 17632 17592 17660
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 20990 17660 20996 17672
rect 20951 17632 20996 17660
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 24026 17660 24032 17672
rect 23987 17632 24032 17660
rect 24026 17620 24032 17632
rect 24084 17620 24090 17672
rect 25222 17592 25228 17604
rect 21881 17564 25228 17592
rect 1535 17527 1593 17533
rect 1535 17493 1547 17527
rect 1581 17524 1593 17527
rect 8938 17524 8944 17536
rect 1581 17496 8944 17524
rect 1581 17493 1593 17496
rect 1535 17487 1593 17493
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 15838 17524 15844 17536
rect 15799 17496 15844 17524
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 16298 17524 16304 17536
rect 16259 17496 16304 17524
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 18049 17527 18107 17533
rect 18049 17524 18061 17527
rect 16540 17496 18061 17524
rect 16540 17484 16546 17496
rect 18049 17493 18061 17496
rect 18095 17524 18107 17527
rect 18506 17524 18512 17536
rect 18095 17496 18512 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 19426 17524 19432 17536
rect 19387 17496 19432 17524
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 19935 17527 19993 17533
rect 19935 17493 19947 17527
rect 19981 17524 19993 17527
rect 21881 17524 21909 17564
rect 25222 17552 25228 17564
rect 25280 17552 25286 17604
rect 19981 17496 21909 17524
rect 19981 17493 19993 17496
rect 19935 17487 19993 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1118 17280 1124 17332
rect 1176 17320 1182 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1176 17292 1593 17320
rect 1176 17280 1182 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 2406 17320 2412 17332
rect 2367 17292 2412 17320
rect 1581 17283 1639 17289
rect 2406 17280 2412 17292
rect 2464 17280 2470 17332
rect 15841 17323 15899 17329
rect 15841 17289 15853 17323
rect 15887 17320 15899 17323
rect 16114 17320 16120 17332
rect 15887 17292 16120 17320
rect 15887 17289 15899 17292
rect 15841 17283 15899 17289
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16298 17320 16304 17332
rect 16255 17292 16304 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 20349 17323 20407 17329
rect 20349 17289 20361 17323
rect 20395 17320 20407 17323
rect 20714 17320 20720 17332
rect 20395 17292 20720 17320
rect 20395 17289 20407 17292
rect 20349 17283 20407 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17320 20867 17323
rect 22278 17320 22284 17332
rect 20855 17292 22284 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 22278 17280 22284 17292
rect 22336 17280 22342 17332
rect 22554 17320 22560 17332
rect 22515 17292 22560 17320
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 23937 17323 23995 17329
rect 23937 17289 23949 17323
rect 23983 17320 23995 17323
rect 24026 17320 24032 17332
rect 23983 17292 24032 17320
rect 23983 17289 23995 17292
rect 23937 17283 23995 17289
rect 24026 17280 24032 17292
rect 24084 17280 24090 17332
rect 16945 17255 17003 17261
rect 16945 17221 16957 17255
rect 16991 17252 17003 17255
rect 17494 17252 17500 17264
rect 16991 17224 17500 17252
rect 16991 17221 17003 17224
rect 16945 17215 17003 17221
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 19978 17212 19984 17264
rect 20036 17252 20042 17264
rect 24673 17255 24731 17261
rect 24673 17252 24685 17255
rect 20036 17224 24685 17252
rect 20036 17212 20042 17224
rect 24673 17221 24685 17224
rect 24719 17252 24731 17255
rect 24762 17252 24768 17264
rect 24719 17224 24768 17252
rect 24719 17221 24731 17224
rect 24673 17215 24731 17221
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 16390 17184 16396 17196
rect 16303 17156 16396 17184
rect 16390 17144 16396 17156
rect 16448 17184 16454 17196
rect 17586 17184 17592 17196
rect 16448 17156 17592 17184
rect 16448 17144 16454 17156
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 21048 17156 21557 17184
rect 21048 17144 21054 17156
rect 21545 17153 21557 17156
rect 21591 17184 21603 17187
rect 21634 17184 21640 17196
rect 21591 17156 21640 17184
rect 21591 17153 21603 17156
rect 21545 17147 21603 17153
rect 21634 17144 21640 17156
rect 21692 17144 21698 17196
rect 24118 17184 24124 17196
rect 24031 17156 24124 17184
rect 24118 17144 24124 17156
rect 24176 17184 24182 17196
rect 25593 17187 25651 17193
rect 25593 17184 25605 17187
rect 24176 17156 25605 17184
rect 24176 17144 24182 17156
rect 25593 17153 25605 17156
rect 25639 17153 25651 17187
rect 25593 17147 25651 17153
rect 2016 17119 2074 17125
rect 2016 17085 2028 17119
rect 2062 17116 2074 17119
rect 2406 17116 2412 17128
rect 2062 17088 2412 17116
rect 2062 17085 2074 17088
rect 2016 17079 2074 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 12253 17119 12311 17125
rect 12253 17085 12265 17119
rect 12299 17116 12311 17119
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12299 17088 12633 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12621 17085 12633 17088
rect 12667 17116 12679 17119
rect 12894 17116 12900 17128
rect 12667 17088 12900 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 14645 17119 14703 17125
rect 14645 17085 14657 17119
rect 14691 17116 14703 17119
rect 15378 17116 15384 17128
rect 14691 17088 15384 17116
rect 14691 17085 14703 17088
rect 14645 17079 14703 17085
rect 15378 17076 15384 17088
rect 15436 17076 15442 17128
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19426 17116 19432 17128
rect 19116 17088 19432 17116
rect 19116 17076 19122 17088
rect 19426 17076 19432 17088
rect 19484 17076 19490 17128
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 23014 17116 23020 17128
rect 22612 17088 23020 17116
rect 22612 17076 22618 17088
rect 23014 17076 23020 17088
rect 23072 17076 23078 17128
rect 15470 17048 15476 17060
rect 15431 17020 15476 17048
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 16485 17051 16543 17057
rect 16485 17017 16497 17051
rect 16531 17017 16543 17051
rect 19334 17048 19340 17060
rect 19247 17020 19340 17048
rect 16485 17011 16543 17017
rect 1946 16940 1952 16992
rect 2004 16980 2010 16992
rect 2087 16983 2145 16989
rect 2087 16980 2099 16983
rect 2004 16952 2099 16980
rect 2004 16940 2010 16952
rect 2087 16949 2099 16952
rect 2133 16949 2145 16983
rect 12986 16980 12992 16992
rect 12947 16952 12992 16980
rect 2087 16943 2145 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 16500 16980 16528 17011
rect 19334 17008 19340 17020
rect 19392 17048 19398 17060
rect 19791 17051 19849 17057
rect 19791 17048 19803 17051
rect 19392 17020 19803 17048
rect 19392 17008 19398 17020
rect 19791 17017 19803 17020
rect 19837 17048 19849 17051
rect 20809 17051 20867 17057
rect 20809 17048 20821 17051
rect 19837 17020 20821 17048
rect 19837 17017 19849 17020
rect 19791 17011 19849 17017
rect 20809 17017 20821 17020
rect 20855 17017 20867 17051
rect 21266 17048 21272 17060
rect 21227 17020 21272 17048
rect 20809 17011 20867 17017
rect 21266 17008 21272 17020
rect 21324 17008 21330 17060
rect 21361 17051 21419 17057
rect 21361 17017 21373 17051
rect 21407 17017 21419 17051
rect 21361 17011 21419 17017
rect 24213 17051 24271 17057
rect 24213 17017 24225 17051
rect 24259 17017 24271 17051
rect 24213 17011 24271 17017
rect 18874 16980 18880 16992
rect 16356 16952 16528 16980
rect 18835 16952 18880 16980
rect 16356 16940 16362 16952
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 20530 16940 20536 16992
rect 20588 16980 20594 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20588 16952 21097 16980
rect 20588 16940 20594 16952
rect 21085 16949 21097 16952
rect 21131 16980 21143 16983
rect 21376 16980 21404 17011
rect 23382 16980 23388 16992
rect 21131 16952 21404 16980
rect 23343 16952 23388 16980
rect 21131 16949 21143 16952
rect 21085 16943 21143 16949
rect 23382 16940 23388 16952
rect 23440 16940 23446 16992
rect 24026 16940 24032 16992
rect 24084 16980 24090 16992
rect 24228 16980 24256 17011
rect 24084 16952 24256 16980
rect 24084 16940 24090 16952
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 16390 16776 16396 16788
rect 16351 16748 16396 16776
rect 16390 16736 16396 16748
rect 16448 16736 16454 16788
rect 19889 16779 19947 16785
rect 19889 16745 19901 16779
rect 19935 16776 19947 16779
rect 19978 16776 19984 16788
rect 19935 16748 19984 16776
rect 19935 16745 19947 16748
rect 19889 16739 19947 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 20990 16776 20996 16788
rect 20763 16748 20996 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 20990 16736 20996 16748
rect 21048 16736 21054 16788
rect 21266 16736 21272 16788
rect 21324 16776 21330 16788
rect 21913 16779 21971 16785
rect 21913 16776 21925 16779
rect 21324 16748 21925 16776
rect 21324 16736 21330 16748
rect 21913 16745 21925 16748
rect 21959 16745 21971 16779
rect 24118 16776 24124 16788
rect 24079 16748 24124 16776
rect 21913 16739 21971 16745
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 12986 16708 12992 16720
rect 12947 16680 12992 16708
rect 12986 16668 12992 16680
rect 13044 16668 13050 16720
rect 13538 16708 13544 16720
rect 13499 16680 13544 16708
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 15378 16668 15384 16720
rect 15436 16708 15442 16720
rect 15473 16711 15531 16717
rect 15473 16708 15485 16711
rect 15436 16680 15485 16708
rect 15436 16668 15442 16680
rect 15473 16677 15485 16680
rect 15519 16677 15531 16711
rect 15473 16671 15531 16677
rect 16114 16668 16120 16720
rect 16172 16708 16178 16720
rect 16942 16708 16948 16720
rect 16172 16680 16948 16708
rect 16172 16668 16178 16680
rect 16942 16668 16948 16680
rect 17000 16708 17006 16720
rect 17037 16711 17095 16717
rect 17037 16708 17049 16711
rect 17000 16680 17049 16708
rect 17000 16668 17006 16680
rect 17037 16677 17049 16680
rect 17083 16677 17095 16711
rect 17037 16671 17095 16677
rect 18963 16711 19021 16717
rect 18963 16677 18975 16711
rect 19009 16708 19021 16711
rect 19334 16708 19340 16720
rect 19009 16680 19340 16708
rect 19009 16677 19021 16680
rect 18963 16671 19021 16677
rect 19334 16668 19340 16680
rect 19392 16668 19398 16720
rect 21082 16708 21088 16720
rect 21043 16680 21088 16708
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 21634 16708 21640 16720
rect 21595 16680 21640 16708
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 22462 16668 22468 16720
rect 22520 16708 22526 16720
rect 23017 16711 23075 16717
rect 23017 16708 23029 16711
rect 22520 16680 23029 16708
rect 22520 16668 22526 16680
rect 23017 16677 23029 16680
rect 23063 16677 23075 16711
rect 23017 16671 23075 16677
rect 23382 16668 23388 16720
rect 23440 16708 23446 16720
rect 24581 16711 24639 16717
rect 24581 16708 24593 16711
rect 23440 16680 24593 16708
rect 23440 16668 23446 16680
rect 24581 16677 24593 16680
rect 24627 16708 24639 16711
rect 24946 16708 24952 16720
rect 24627 16680 24952 16708
rect 24627 16677 24639 16680
rect 24581 16671 24639 16677
rect 24946 16668 24952 16680
rect 25004 16668 25010 16720
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16572 11851 16575
rect 12250 16572 12256 16584
rect 11839 16544 12256 16572
rect 11839 16541 11851 16544
rect 11793 16535 11851 16541
rect 12250 16532 12256 16544
rect 12308 16572 12314 16584
rect 12897 16575 12955 16581
rect 12897 16572 12909 16575
rect 12308 16544 12909 16572
rect 12308 16532 12314 16544
rect 12897 16541 12909 16544
rect 12943 16541 12955 16575
rect 12897 16535 12955 16541
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 14792 16544 15393 16572
rect 14792 16532 14798 16544
rect 15381 16541 15393 16544
rect 15427 16541 15439 16575
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 15381 16535 15439 16541
rect 16022 16532 16028 16544
rect 16080 16572 16086 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16080 16544 16957 16572
rect 16080 16532 16086 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 18598 16572 18604 16584
rect 18559 16544 18604 16572
rect 16945 16535 17003 16541
rect 18598 16532 18604 16544
rect 18656 16532 18662 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16572 21051 16575
rect 21358 16572 21364 16584
rect 21039 16544 21364 16572
rect 21039 16541 21051 16544
rect 20993 16535 21051 16541
rect 21358 16532 21364 16544
rect 21416 16532 21422 16584
rect 22922 16572 22928 16584
rect 22883 16544 22928 16572
rect 22922 16532 22928 16544
rect 22980 16532 22986 16584
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 24489 16575 24547 16581
rect 24489 16572 24501 16575
rect 23615 16544 24501 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 24489 16541 24501 16544
rect 24535 16541 24547 16575
rect 24762 16572 24768 16584
rect 24723 16544 24768 16572
rect 24489 16535 24547 16541
rect 17494 16504 17500 16516
rect 17455 16476 17500 16504
rect 17494 16464 17500 16476
rect 17552 16464 17558 16516
rect 19521 16507 19579 16513
rect 19521 16473 19533 16507
rect 19567 16504 19579 16507
rect 20530 16504 20536 16516
rect 19567 16476 20536 16504
rect 19567 16473 19579 16476
rect 19521 16467 19579 16473
rect 20530 16464 20536 16476
rect 20588 16464 20594 16516
rect 24504 16504 24532 16535
rect 24762 16532 24768 16544
rect 24820 16532 24826 16584
rect 24670 16504 24676 16516
rect 24504 16476 24676 16504
rect 24670 16464 24676 16476
rect 24728 16464 24734 16516
rect 15838 16396 15844 16448
rect 15896 16436 15902 16448
rect 18322 16436 18328 16448
rect 15896 16408 18328 16436
rect 15896 16396 15902 16408
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 12250 16232 12256 16244
rect 12211 16204 12256 16232
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 12986 16232 12992 16244
rect 12759 16204 12992 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 14734 16232 14740 16244
rect 14695 16204 14740 16232
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 15470 16232 15476 16244
rect 15431 16204 15476 16232
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 16942 16232 16948 16244
rect 16903 16204 16948 16232
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 19334 16232 19340 16244
rect 19295 16204 19340 16232
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 21683 16235 21741 16241
rect 21683 16201 21695 16235
rect 21729 16232 21741 16235
rect 24210 16232 24216 16244
rect 21729 16204 24216 16232
rect 21729 16201 21741 16204
rect 21683 16195 21741 16201
rect 24210 16192 24216 16204
rect 24268 16192 24274 16244
rect 24857 16235 24915 16241
rect 24857 16201 24869 16235
rect 24903 16232 24915 16235
rect 24946 16232 24952 16244
rect 24903 16204 24952 16232
rect 24903 16201 24915 16204
rect 24857 16195 24915 16201
rect 24946 16192 24952 16204
rect 25004 16192 25010 16244
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 25455 16235 25513 16241
rect 25455 16232 25467 16235
rect 25096 16204 25467 16232
rect 25096 16192 25102 16204
rect 25455 16201 25467 16204
rect 25501 16201 25513 16235
rect 25455 16195 25513 16201
rect 22462 16164 22468 16176
rect 15764 16136 17356 16164
rect 22423 16136 22468 16164
rect 13538 16096 13544 16108
rect 13499 16068 13544 16096
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 15764 16105 15792 16136
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 16022 16096 16028 16108
rect 15983 16068 16028 16096
rect 15749 16059 15807 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 12894 15960 12900 15972
rect 12855 15932 12900 15960
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 12986 15920 12992 15972
rect 13044 15960 13050 15972
rect 15841 15963 15899 15969
rect 13044 15932 13089 15960
rect 13044 15920 13050 15932
rect 15841 15929 15853 15963
rect 15887 15929 15899 15963
rect 15841 15923 15899 15929
rect 13004 15892 13032 15920
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13004 15864 13829 15892
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15378 15892 15384 15904
rect 15243 15864 15384 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 15470 15852 15476 15904
rect 15528 15892 15534 15904
rect 15856 15892 15884 15923
rect 17328 15901 17356 16136
rect 22462 16124 22468 16136
rect 22520 16124 22526 16176
rect 19058 16096 19064 16108
rect 19019 16068 19064 16096
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16096 20683 16099
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20671 16068 20913 16096
rect 20671 16065 20683 16068
rect 20625 16059 20683 16065
rect 20901 16065 20913 16068
rect 20947 16096 20959 16099
rect 21082 16096 21088 16108
rect 20947 16068 21088 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 21358 16096 21364 16108
rect 21271 16068 21364 16096
rect 21358 16056 21364 16068
rect 21416 16096 21422 16108
rect 22695 16099 22753 16105
rect 22695 16096 22707 16099
rect 21416 16068 22707 16096
rect 21416 16056 21422 16068
rect 22695 16065 22707 16068
rect 22741 16065 22753 16099
rect 22695 16059 22753 16065
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16096 23903 16099
rect 25222 16096 25228 16108
rect 23891 16068 25228 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 25222 16056 25228 16068
rect 25280 16056 25286 16108
rect 18322 16028 18328 16040
rect 18283 16000 18328 16028
rect 18322 15988 18328 16000
rect 18380 15988 18386 16040
rect 18785 16031 18843 16037
rect 18785 16028 18797 16031
rect 18524 16000 18797 16028
rect 18524 15904 18552 16000
rect 18785 15997 18797 16000
rect 18831 15997 18843 16031
rect 18785 15991 18843 15997
rect 19797 16031 19855 16037
rect 19797 15997 19809 16031
rect 19843 16028 19855 16031
rect 20530 16028 20536 16040
rect 19843 16000 20536 16028
rect 19843 15997 19855 16000
rect 19797 15991 19855 15997
rect 20530 15988 20536 16000
rect 20588 15988 20594 16040
rect 21612 16031 21670 16037
rect 21612 15997 21624 16031
rect 21658 16028 21670 16031
rect 22608 16031 22666 16037
rect 21658 16000 22140 16028
rect 21658 15997 21670 16000
rect 21612 15991 21670 15997
rect 15528 15864 15884 15892
rect 17313 15895 17371 15901
rect 15528 15852 15534 15864
rect 17313 15861 17325 15895
rect 17359 15892 17371 15895
rect 17678 15892 17684 15904
rect 17359 15864 17684 15892
rect 17359 15861 17371 15864
rect 17313 15855 17371 15861
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 17865 15895 17923 15901
rect 17865 15861 17877 15895
rect 17911 15892 17923 15895
rect 18506 15892 18512 15904
rect 17911 15864 18512 15892
rect 17911 15861 17923 15864
rect 17865 15855 17923 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 22112 15901 22140 16000
rect 22608 15997 22620 16031
rect 22654 16028 22666 16031
rect 25384 16031 25442 16037
rect 22654 16000 23152 16028
rect 22654 15997 22666 16000
rect 22608 15991 22666 15997
rect 23124 15904 23152 16000
rect 25384 15997 25396 16031
rect 25430 16028 25442 16031
rect 25430 16000 25912 16028
rect 25430 15997 25442 16000
rect 25384 15991 25442 15997
rect 23934 15920 23940 15972
rect 23992 15960 23998 15972
rect 24486 15960 24492 15972
rect 23992 15932 24037 15960
rect 24447 15932 24492 15960
rect 23992 15920 23998 15932
rect 24486 15920 24492 15932
rect 24544 15920 24550 15972
rect 22097 15895 22155 15901
rect 22097 15861 22109 15895
rect 22143 15892 22155 15895
rect 22186 15892 22192 15904
rect 22143 15864 22192 15892
rect 22143 15861 22155 15864
rect 22097 15855 22155 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23106 15892 23112 15904
rect 23067 15864 23112 15892
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 23477 15895 23535 15901
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 23952 15892 23980 15920
rect 25884 15904 25912 16000
rect 25222 15892 25228 15904
rect 23523 15864 23980 15892
rect 25183 15864 25228 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 25222 15852 25228 15864
rect 25280 15852 25286 15904
rect 25866 15892 25872 15904
rect 25827 15864 25872 15892
rect 25866 15852 25872 15864
rect 25924 15852 25930 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 12618 15688 12624 15700
rect 12579 15660 12624 15688
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12952 15660 13461 15688
rect 12952 15648 12958 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 13449 15651 13507 15657
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15688 14427 15691
rect 15838 15688 15844 15700
rect 14415 15660 15844 15688
rect 14415 15657 14427 15660
rect 14369 15651 14427 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 16022 15648 16028 15700
rect 16080 15688 16086 15700
rect 16853 15691 16911 15697
rect 16853 15688 16865 15691
rect 16080 15660 16865 15688
rect 16080 15648 16086 15660
rect 16853 15657 16865 15660
rect 16899 15657 16911 15691
rect 17862 15688 17868 15700
rect 17823 15660 17868 15688
rect 16853 15651 16911 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 23293 15691 23351 15697
rect 23293 15657 23305 15691
rect 23339 15688 23351 15691
rect 23382 15688 23388 15700
rect 23339 15660 23388 15688
rect 23339 15657 23351 15660
rect 23293 15651 23351 15657
rect 23382 15648 23388 15660
rect 23440 15648 23446 15700
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 25133 15691 25191 15697
rect 25133 15688 25145 15691
rect 24544 15660 25145 15688
rect 24544 15648 24550 15660
rect 25133 15657 25145 15660
rect 25179 15657 25191 15691
rect 25133 15651 25191 15657
rect 15651 15623 15709 15629
rect 15651 15589 15663 15623
rect 15697 15620 15709 15623
rect 15930 15620 15936 15632
rect 15697 15592 15936 15620
rect 15697 15589 15709 15592
rect 15651 15583 15709 15589
rect 15930 15580 15936 15592
rect 15988 15580 15994 15632
rect 22278 15580 22284 15632
rect 22336 15620 22342 15632
rect 22694 15623 22752 15629
rect 22694 15620 22706 15623
rect 22336 15592 22706 15620
rect 22336 15580 22342 15592
rect 22694 15589 22706 15592
rect 22740 15589 22752 15623
rect 22694 15583 22752 15589
rect 22922 15580 22928 15632
rect 22980 15620 22986 15632
rect 23569 15623 23627 15629
rect 23569 15620 23581 15623
rect 22980 15592 23581 15620
rect 22980 15580 22986 15592
rect 23569 15589 23581 15592
rect 23615 15589 23627 15623
rect 23569 15583 23627 15589
rect 23934 15580 23940 15632
rect 23992 15620 23998 15632
rect 24121 15623 24179 15629
rect 24121 15620 24133 15623
rect 23992 15592 24133 15620
rect 23992 15580 23998 15592
rect 24121 15589 24133 15592
rect 24167 15589 24179 15623
rect 24121 15583 24179 15589
rect 12986 15512 12992 15564
rect 13044 15552 13050 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 13044 15524 13185 15552
rect 13044 15512 13050 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 13173 15515 13231 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 16172 15524 16221 15552
rect 16172 15512 16178 15524
rect 16209 15521 16221 15524
rect 16255 15521 16267 15555
rect 16209 15515 16267 15521
rect 16942 15512 16948 15564
rect 17000 15552 17006 15564
rect 17037 15555 17095 15561
rect 17037 15552 17049 15555
rect 17000 15524 17049 15552
rect 17000 15512 17006 15524
rect 17037 15521 17049 15524
rect 17083 15521 17095 15555
rect 18322 15552 18328 15564
rect 18283 15524 18328 15552
rect 17037 15515 17095 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 18506 15552 18512 15564
rect 18467 15524 18512 15552
rect 18506 15512 18512 15524
rect 18564 15512 18570 15564
rect 24762 15552 24768 15564
rect 24723 15524 24768 15552
rect 24762 15512 24768 15524
rect 24820 15512 24826 15564
rect 12250 15484 12256 15496
rect 12211 15456 12256 15484
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 15286 15484 15292 15496
rect 15247 15456 15292 15484
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 18598 15484 18604 15496
rect 18559 15456 18604 15484
rect 18598 15444 18604 15456
rect 18656 15484 18662 15496
rect 19061 15487 19119 15493
rect 19061 15484 19073 15487
rect 18656 15456 19073 15484
rect 18656 15444 18662 15456
rect 19061 15453 19073 15456
rect 19107 15453 19119 15487
rect 22370 15484 22376 15496
rect 22331 15456 22376 15484
rect 19061 15447 19119 15453
rect 22370 15444 22376 15456
rect 22428 15444 22434 15496
rect 17221 15419 17279 15425
rect 17221 15385 17233 15419
rect 17267 15416 17279 15419
rect 17770 15416 17776 15428
rect 17267 15388 17776 15416
rect 17267 15385 17279 15388
rect 17221 15379 17279 15385
rect 17770 15376 17776 15388
rect 17828 15416 17834 15428
rect 18322 15416 18328 15428
rect 17828 15388 18328 15416
rect 17828 15376 17834 15388
rect 18322 15376 18328 15388
rect 18380 15376 18386 15428
rect 16574 15348 16580 15360
rect 16535 15320 16580 15348
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 19978 15348 19984 15360
rect 19939 15320 19984 15348
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 21634 15308 21640 15360
rect 21692 15348 21698 15360
rect 21821 15351 21879 15357
rect 21821 15348 21833 15351
rect 21692 15320 21833 15348
rect 21692 15308 21698 15320
rect 21821 15317 21833 15320
rect 21867 15317 21879 15351
rect 21821 15311 21879 15317
rect 24029 15351 24087 15357
rect 24029 15317 24041 15351
rect 24075 15348 24087 15351
rect 24210 15348 24216 15360
rect 24075 15320 24216 15348
rect 24075 15317 24087 15320
rect 24029 15311 24087 15317
rect 24210 15308 24216 15320
rect 24268 15308 24274 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 12158 15104 12164 15156
rect 12216 15144 12222 15156
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 12216 15116 12265 15144
rect 12216 15104 12222 15116
rect 12253 15113 12265 15116
rect 12299 15144 12311 15147
rect 12618 15144 12624 15156
rect 12299 15116 12624 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 15565 15147 15623 15153
rect 15565 15144 15577 15147
rect 15436 15116 15577 15144
rect 15436 15104 15442 15116
rect 15565 15113 15577 15116
rect 15611 15113 15623 15147
rect 15930 15144 15936 15156
rect 15843 15116 15936 15144
rect 15565 15107 15623 15113
rect 15930 15104 15936 15116
rect 15988 15144 15994 15156
rect 18138 15144 18144 15156
rect 15988 15116 18144 15144
rect 15988 15104 15994 15116
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 18322 15104 18328 15156
rect 18380 15144 18386 15156
rect 19153 15147 19211 15153
rect 19153 15144 19165 15147
rect 18380 15116 19165 15144
rect 18380 15104 18386 15116
rect 19153 15113 19165 15116
rect 19199 15113 19211 15147
rect 19153 15107 19211 15113
rect 22462 15104 22468 15156
rect 22520 15144 22526 15156
rect 22741 15147 22799 15153
rect 22741 15144 22753 15147
rect 22520 15116 22753 15144
rect 22520 15104 22526 15116
rect 22741 15113 22753 15116
rect 22787 15144 22799 15147
rect 24762 15144 24768 15156
rect 22787 15116 24768 15144
rect 22787 15113 22799 15116
rect 22741 15107 22799 15113
rect 24762 15104 24768 15116
rect 24820 15144 24826 15156
rect 24949 15147 25007 15153
rect 24949 15144 24961 15147
rect 24820 15116 24961 15144
rect 24820 15104 24826 15116
rect 24949 15113 24961 15116
rect 24995 15113 25007 15147
rect 24949 15107 25007 15113
rect 11514 14968 11520 15020
rect 11572 15008 11578 15020
rect 11885 15011 11943 15017
rect 11885 15008 11897 15011
rect 11572 14980 11897 15008
rect 11572 14968 11578 14980
rect 11885 14977 11897 14980
rect 11931 15008 11943 15011
rect 12618 15008 12624 15020
rect 11931 14980 12624 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 12894 15008 12900 15020
rect 12855 14980 12900 15008
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 18874 15008 18880 15020
rect 17175 14980 18880 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20438 15008 20444 15020
rect 20399 14980 20444 15008
rect 20438 14968 20444 14980
rect 20496 14968 20502 15020
rect 5442 14949 5448 14952
rect 5420 14943 5448 14949
rect 5420 14940 5432 14943
rect 5355 14912 5432 14940
rect 5420 14909 5432 14912
rect 5500 14940 5506 14952
rect 5813 14943 5871 14949
rect 5813 14940 5825 14943
rect 5500 14912 5825 14940
rect 5420 14903 5448 14909
rect 5442 14900 5448 14903
rect 5500 14900 5506 14912
rect 5813 14909 5825 14912
rect 5859 14909 5871 14943
rect 14642 14940 14648 14952
rect 14603 14912 14648 14940
rect 5813 14903 5871 14909
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 15930 14940 15936 14952
rect 14982 14912 15936 14940
rect 5629 14875 5687 14881
rect 5629 14841 5641 14875
rect 5675 14872 5687 14875
rect 12529 14875 12587 14881
rect 12529 14872 12541 14875
rect 5675 14844 12541 14872
rect 5675 14841 5687 14844
rect 5629 14835 5687 14841
rect 12529 14841 12541 14844
rect 12575 14841 12587 14875
rect 12529 14835 12587 14841
rect 12544 14804 12572 14835
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 14982 14881 15010 14912
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 16574 14940 16580 14952
rect 16535 14912 16580 14940
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 17862 14900 17868 14952
rect 17920 14940 17926 14952
rect 17920 14912 18092 14940
rect 17920 14900 17926 14912
rect 14553 14875 14611 14881
rect 12676 14844 12721 14872
rect 12676 14832 12682 14844
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 14967 14875 15025 14881
rect 14967 14872 14979 14875
rect 14599 14844 14979 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 14967 14841 14979 14844
rect 15013 14841 15025 14875
rect 14967 14835 15025 14841
rect 15286 14832 15292 14884
rect 15344 14872 15350 14884
rect 16209 14875 16267 14881
rect 16209 14872 16221 14875
rect 15344 14844 16221 14872
rect 15344 14832 15350 14844
rect 16209 14841 16221 14844
rect 16255 14841 16267 14875
rect 18064 14872 18092 14912
rect 21634 14900 21640 14952
rect 21692 14940 21698 14952
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21692 14912 21833 14940
rect 21692 14900 21698 14912
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 24210 14940 24216 14952
rect 24171 14912 24216 14940
rect 21821 14903 21879 14909
rect 24210 14900 24216 14912
rect 24268 14900 24274 14952
rect 18233 14875 18291 14881
rect 18233 14872 18245 14875
rect 18064 14844 18245 14872
rect 16209 14835 16267 14841
rect 18233 14841 18245 14844
rect 18279 14841 18291 14875
rect 18233 14835 18291 14841
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 18877 14875 18935 14881
rect 18380 14844 18425 14872
rect 18380 14832 18386 14844
rect 18877 14841 18889 14875
rect 18923 14872 18935 14875
rect 19058 14872 19064 14884
rect 18923 14844 19064 14872
rect 18923 14841 18935 14844
rect 18877 14835 18935 14841
rect 19058 14832 19064 14844
rect 19116 14832 19122 14884
rect 19797 14875 19855 14881
rect 19797 14841 19809 14875
rect 19843 14872 19855 14875
rect 20070 14872 20076 14884
rect 19843 14844 20076 14872
rect 19843 14841 19855 14844
rect 19797 14835 19855 14841
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 21729 14875 21787 14881
rect 21729 14841 21741 14875
rect 21775 14872 21787 14875
rect 22183 14875 22241 14881
rect 22183 14872 22195 14875
rect 21775 14844 22195 14872
rect 21775 14841 21787 14844
rect 21729 14835 21787 14841
rect 22183 14841 22195 14844
rect 22229 14872 22241 14875
rect 22278 14872 22284 14884
rect 22229 14844 22284 14872
rect 22229 14841 22241 14844
rect 22183 14835 22241 14841
rect 22278 14832 22284 14844
rect 22336 14872 22342 14884
rect 23017 14875 23075 14881
rect 23017 14872 23029 14875
rect 22336 14844 23029 14872
rect 22336 14832 22342 14844
rect 23017 14841 23029 14844
rect 23063 14841 23075 14875
rect 24670 14872 24676 14884
rect 24631 14844 24676 14872
rect 23017 14835 23075 14841
rect 24670 14832 24676 14844
rect 24728 14832 24734 14884
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 12544 14776 13461 14804
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 14182 14804 14188 14816
rect 14143 14776 14188 14804
rect 13449 14767 13507 14773
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 16942 14804 16948 14816
rect 15712 14776 16948 14804
rect 15712 14764 15718 14776
rect 16942 14764 16948 14776
rect 17000 14804 17006 14816
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17000 14776 17417 14804
rect 17000 14764 17006 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 17405 14767 17463 14773
rect 17865 14807 17923 14813
rect 17865 14773 17877 14807
rect 17911 14804 17923 14807
rect 18506 14804 18512 14816
rect 17911 14776 18512 14804
rect 17911 14773 17923 14776
rect 17865 14767 17923 14773
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 25501 14807 25559 14813
rect 25501 14804 25513 14807
rect 24544 14776 25513 14804
rect 24544 14764 24550 14776
rect 25501 14773 25513 14776
rect 25547 14773 25559 14807
rect 25501 14767 25559 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 12250 14600 12256 14612
rect 12211 14572 12256 14600
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 16632 14572 17877 14600
rect 16632 14560 16638 14572
rect 17865 14569 17877 14572
rect 17911 14600 17923 14603
rect 18230 14600 18236 14612
rect 17911 14572 18236 14600
rect 17911 14569 17923 14572
rect 17865 14563 17923 14569
rect 18230 14560 18236 14572
rect 18288 14560 18294 14612
rect 19797 14603 19855 14609
rect 19797 14569 19809 14603
rect 19843 14600 19855 14603
rect 19978 14600 19984 14612
rect 19843 14572 19984 14600
rect 19843 14569 19855 14572
rect 19797 14563 19855 14569
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 22370 14600 22376 14612
rect 22331 14572 22376 14600
rect 22370 14560 22376 14572
rect 22428 14560 22434 14612
rect 12621 14535 12679 14541
rect 12621 14532 12633 14535
rect 11808 14504 12633 14532
rect 11514 14464 11520 14476
rect 11475 14436 11520 14464
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11808 14408 11836 14504
rect 12621 14501 12633 14504
rect 12667 14501 12679 14535
rect 12621 14495 12679 14501
rect 14200 14504 16068 14532
rect 14200 14476 14228 14504
rect 14182 14464 14188 14476
rect 14095 14436 14188 14464
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 15654 14464 15660 14476
rect 15615 14436 15660 14464
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 16040 14473 16068 14504
rect 18138 14492 18144 14544
rect 18196 14532 18202 14544
rect 18411 14535 18469 14541
rect 18411 14532 18423 14535
rect 18196 14504 18423 14532
rect 18196 14492 18202 14504
rect 18411 14501 18423 14504
rect 18457 14532 18469 14535
rect 19334 14532 19340 14544
rect 18457 14504 19340 14532
rect 18457 14501 18469 14504
rect 18411 14495 18469 14501
rect 19334 14492 19340 14504
rect 19392 14492 19398 14544
rect 20070 14492 20076 14544
rect 20128 14532 20134 14544
rect 20901 14535 20959 14541
rect 20901 14532 20913 14535
rect 20128 14504 20913 14532
rect 20128 14492 20134 14504
rect 20901 14501 20913 14504
rect 20947 14501 20959 14535
rect 20901 14495 20959 14501
rect 22922 14492 22928 14544
rect 22980 14532 22986 14544
rect 23017 14535 23075 14541
rect 23017 14532 23029 14535
rect 22980 14504 23029 14532
rect 22980 14492 22986 14504
rect 23017 14501 23029 14504
rect 23063 14501 23075 14535
rect 23017 14495 23075 14501
rect 24026 14492 24032 14544
rect 24084 14532 24090 14544
rect 24486 14532 24492 14544
rect 24084 14504 24492 14532
rect 24084 14492 24090 14504
rect 24486 14492 24492 14504
rect 24544 14492 24550 14544
rect 24581 14535 24639 14541
rect 24581 14501 24593 14535
rect 24627 14532 24639 14535
rect 24670 14532 24676 14544
rect 24627 14504 24676 14532
rect 24627 14501 24639 14504
rect 24581 14495 24639 14501
rect 24670 14492 24676 14504
rect 24728 14492 24734 14544
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16071 14436 16865 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16853 14433 16865 14436
rect 16899 14464 16911 14467
rect 17402 14464 17408 14476
rect 16899 14436 17408 14464
rect 16899 14433 16911 14436
rect 16853 14427 16911 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 21542 14464 21548 14476
rect 21503 14436 21548 14464
rect 21542 14424 21548 14436
rect 21600 14424 21606 14476
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 11790 14396 11796 14408
rect 11655 14368 11796 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 12894 14396 12900 14408
rect 12575 14368 12801 14396
rect 12855 14368 12900 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 12773 14328 12801 14368
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 18049 14399 18107 14405
rect 18049 14396 18061 14399
rect 17184 14368 18061 14396
rect 17184 14356 17190 14368
rect 18049 14365 18061 14368
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 22925 14399 22983 14405
rect 22925 14396 22937 14399
rect 22796 14368 22937 14396
rect 22796 14356 22802 14368
rect 22925 14365 22937 14368
rect 22971 14365 22983 14399
rect 23566 14396 23572 14408
rect 23527 14368 23572 14396
rect 22925 14359 22983 14365
rect 23566 14356 23572 14368
rect 23624 14356 23630 14408
rect 23658 14356 23664 14408
rect 23716 14396 23722 14408
rect 24762 14396 24768 14408
rect 23716 14368 24768 14396
rect 23716 14356 23722 14368
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 13538 14328 13544 14340
rect 12773 14300 13544 14328
rect 13538 14288 13544 14300
rect 13596 14288 13602 14340
rect 16390 14288 16396 14340
rect 16448 14328 16454 14340
rect 17037 14331 17095 14337
rect 17037 14328 17049 14331
rect 16448 14300 17049 14328
rect 16448 14288 16454 14300
rect 17037 14297 17049 14300
rect 17083 14297 17095 14331
rect 17037 14291 17095 14297
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 14642 14260 14648 14272
rect 14603 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 16482 14260 16488 14272
rect 16443 14232 16488 14260
rect 16482 14220 16488 14232
rect 16540 14220 16546 14272
rect 18969 14263 19027 14269
rect 18969 14229 18981 14263
rect 19015 14260 19027 14263
rect 19518 14260 19524 14272
rect 19015 14232 19524 14260
rect 19015 14229 19027 14232
rect 18969 14223 19027 14229
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 24210 14260 24216 14272
rect 24171 14232 24216 14260
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 10965 14059 11023 14065
rect 10965 14025 10977 14059
rect 11011 14056 11023 14059
rect 11514 14056 11520 14068
rect 11011 14028 11520 14056
rect 11011 14025 11023 14028
rect 10965 14019 11023 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 12676 14028 13369 14056
rect 12676 14016 12682 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 14182 14056 14188 14068
rect 14143 14028 14188 14056
rect 13357 14019 13415 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17865 14059 17923 14065
rect 17865 14025 17877 14059
rect 17911 14056 17923 14059
rect 18138 14056 18144 14068
rect 17911 14028 18144 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 18969 14059 19027 14065
rect 18969 14056 18981 14059
rect 18288 14028 18981 14056
rect 18288 14016 18294 14028
rect 18969 14025 18981 14028
rect 19015 14025 19027 14059
rect 18969 14019 19027 14025
rect 21542 14016 21548 14068
rect 21600 14056 21606 14068
rect 22465 14059 22523 14065
rect 22465 14056 22477 14059
rect 21600 14028 22477 14056
rect 21600 14016 21606 14028
rect 22465 14025 22477 14028
rect 22511 14025 22523 14059
rect 22465 14019 22523 14025
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 23201 14059 23259 14065
rect 23201 14056 23213 14059
rect 22796 14028 23213 14056
rect 22796 14016 22802 14028
rect 23201 14025 23213 14028
rect 23247 14025 23259 14059
rect 24026 14056 24032 14068
rect 23987 14028 24032 14056
rect 23201 14019 23259 14025
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 24670 14016 24676 14068
rect 24728 14056 24734 14068
rect 25133 14059 25191 14065
rect 25133 14056 25145 14059
rect 24728 14028 25145 14056
rect 24728 14016 24734 14028
rect 25133 14025 25145 14028
rect 25179 14025 25191 14059
rect 25133 14019 25191 14025
rect 20438 13988 20444 14000
rect 20399 13960 20444 13988
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 22370 13988 22376 14000
rect 22112 13960 22376 13988
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 15286 13920 15292 13932
rect 12308 13892 14412 13920
rect 15247 13892 15292 13920
rect 12308 13880 12314 13892
rect 14384 13864 14412 13892
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 17126 13920 17132 13932
rect 17087 13892 17132 13920
rect 17126 13880 17132 13892
rect 17184 13920 17190 13932
rect 22112 13929 22140 13960
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 24762 13988 24768 14000
rect 24723 13960 24768 13988
rect 24762 13948 24768 13960
rect 24820 13948 24826 14000
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 17184 13892 19257 13920
rect 17184 13880 17190 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 19245 13883 19303 13889
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 23566 13880 23572 13932
rect 23624 13920 23630 13932
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 23624 13892 24225 13920
rect 23624 13880 23630 13892
rect 24213 13889 24225 13892
rect 24259 13920 24271 13923
rect 24578 13920 24584 13932
rect 24259 13892 24584 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 24578 13880 24584 13892
rect 24636 13920 24642 13932
rect 25501 13923 25559 13929
rect 25501 13920 25513 13923
rect 24636 13892 25513 13920
rect 24636 13880 24642 13892
rect 25501 13889 25513 13892
rect 25547 13889 25559 13923
rect 25501 13883 25559 13889
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12526 13852 12532 13864
rect 12483 13824 12532 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14424 13824 14657 13852
rect 14424 13812 14430 13824
rect 14645 13821 14657 13824
rect 14691 13852 14703 13855
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14691 13824 14749 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 14737 13815 14795 13821
rect 14826 13812 14832 13864
rect 14884 13852 14890 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 14884 13824 15209 13852
rect 14884 13812 14890 13824
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16390 13852 16396 13864
rect 16347 13824 16396 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 16850 13852 16856 13864
rect 16540 13824 16856 13852
rect 16540 13812 16546 13824
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13821 21695 13855
rect 21818 13852 21824 13864
rect 21779 13824 21824 13852
rect 21637 13815 21695 13821
rect 12758 13787 12816 13793
rect 12758 13784 12770 13787
rect 12176 13756 12770 13784
rect 12176 13728 12204 13756
rect 12758 13753 12770 13756
rect 12804 13753 12816 13787
rect 12758 13747 12816 13753
rect 18138 13744 18144 13796
rect 18196 13784 18202 13796
rect 18370 13787 18428 13793
rect 18370 13784 18382 13787
rect 18196 13756 18382 13784
rect 18196 13744 18202 13756
rect 18370 13753 18382 13756
rect 18416 13753 18428 13787
rect 18370 13747 18428 13753
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 19334 13784 19340 13796
rect 19116 13756 19340 13784
rect 19116 13744 19122 13756
rect 19334 13744 19340 13756
rect 19392 13784 19398 13796
rect 19889 13787 19947 13793
rect 19889 13784 19901 13787
rect 19392 13756 19901 13784
rect 19392 13744 19398 13756
rect 19889 13753 19901 13756
rect 19935 13753 19947 13787
rect 19889 13747 19947 13753
rect 19981 13787 20039 13793
rect 19981 13753 19993 13787
rect 20027 13784 20039 13787
rect 21542 13784 21548 13796
rect 20027 13756 21548 13784
rect 20027 13753 20039 13756
rect 19981 13747 20039 13753
rect 12158 13716 12164 13728
rect 12119 13688 12164 13716
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13596 13688 13645 13716
rect 13596 13676 13602 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13633 13679 13691 13685
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15712 13688 15761 13716
rect 15712 13676 15718 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 19705 13719 19763 13725
rect 19705 13716 19717 13719
rect 19576 13688 19717 13716
rect 19576 13676 19582 13688
rect 19705 13685 19717 13688
rect 19751 13716 19763 13719
rect 19996 13716 20024 13747
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 19751 13688 20024 13716
rect 19751 13685 19763 13688
rect 19705 13679 19763 13685
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 20680 13688 20821 13716
rect 20680 13676 20686 13688
rect 20809 13685 20821 13688
rect 20855 13685 20867 13719
rect 21174 13716 21180 13728
rect 21135 13688 21180 13716
rect 20809 13679 20867 13685
rect 21174 13676 21180 13688
rect 21232 13716 21238 13728
rect 21652 13716 21680 13815
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 24302 13784 24308 13796
rect 24263 13756 24308 13784
rect 24302 13744 24308 13756
rect 24360 13744 24366 13796
rect 22830 13716 22836 13728
rect 21232 13688 21680 13716
rect 22791 13688 22836 13716
rect 21232 13676 21238 13688
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 12342 13512 12348 13524
rect 12303 13484 12348 13512
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 15841 13515 15899 13521
rect 15841 13481 15853 13515
rect 15887 13512 15899 13515
rect 18138 13512 18144 13524
rect 15887 13484 16712 13512
rect 18099 13484 18144 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 14369 13447 14427 13453
rect 14369 13413 14381 13447
rect 14415 13444 14427 13447
rect 14642 13444 14648 13456
rect 14415 13416 14648 13444
rect 14415 13413 14427 13416
rect 14369 13407 14427 13413
rect 14642 13404 14648 13416
rect 14700 13404 14706 13456
rect 16684 13388 16712 13484
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 22738 13472 22744 13524
rect 22796 13512 22802 13524
rect 22833 13515 22891 13521
rect 22833 13512 22845 13515
rect 22796 13484 22845 13512
rect 22796 13472 22802 13484
rect 22833 13481 22845 13484
rect 22879 13481 22891 13515
rect 22833 13475 22891 13481
rect 23385 13515 23443 13521
rect 23385 13481 23397 13515
rect 23431 13512 23443 13515
rect 24302 13512 24308 13524
rect 23431 13484 24308 13512
rect 23431 13481 23443 13484
rect 23385 13475 23443 13481
rect 24302 13472 24308 13484
rect 24360 13472 24366 13524
rect 17405 13447 17463 13453
rect 17405 13413 17417 13447
rect 17451 13444 17463 13447
rect 18046 13444 18052 13456
rect 17451 13416 18052 13444
rect 17451 13413 17463 13416
rect 17405 13407 17463 13413
rect 18046 13404 18052 13416
rect 18104 13444 18110 13456
rect 18417 13447 18475 13453
rect 18417 13444 18429 13447
rect 18104 13416 18429 13444
rect 18104 13404 18110 13416
rect 18417 13413 18429 13416
rect 18463 13413 18475 13447
rect 18417 13407 18475 13413
rect 18874 13404 18880 13456
rect 18932 13444 18938 13456
rect 19153 13447 19211 13453
rect 19153 13444 19165 13447
rect 18932 13416 19165 13444
rect 18932 13404 18938 13416
rect 19153 13413 19165 13416
rect 19199 13413 19211 13447
rect 21634 13444 21640 13456
rect 21595 13416 21640 13444
rect 19153 13407 19211 13413
rect 21634 13404 21640 13416
rect 21692 13404 21698 13456
rect 24397 13447 24455 13453
rect 24397 13413 24409 13447
rect 24443 13444 24455 13447
rect 24670 13444 24676 13456
rect 24443 13416 24676 13444
rect 24443 13413 24455 13416
rect 24397 13407 24455 13413
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 12250 13376 12256 13388
rect 12211 13348 12256 13376
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 12618 13376 12624 13388
rect 12579 13348 12624 13376
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 13906 13376 13912 13388
rect 13867 13348 13912 13376
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 14826 13376 14832 13388
rect 14231 13348 14832 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16666 13376 16672 13388
rect 16579 13348 16672 13376
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17129 13379 17187 13385
rect 17129 13376 17141 13379
rect 16908 13348 17141 13376
rect 16908 13336 16914 13348
rect 17129 13345 17141 13348
rect 17175 13345 17187 13379
rect 17129 13339 17187 13345
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20404 13348 20913 13376
rect 20404 13336 20410 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 21361 13379 21419 13385
rect 21361 13345 21373 13379
rect 21407 13376 21419 13379
rect 21818 13376 21824 13388
rect 21407 13348 21824 13376
rect 21407 13345 21419 13348
rect 21361 13339 21419 13345
rect 19058 13308 19064 13320
rect 19019 13280 19064 13308
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19334 13308 19340 13320
rect 19295 13280 19340 13308
rect 19334 13268 19340 13280
rect 19392 13308 19398 13320
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19392 13280 19993 13308
rect 19392 13268 19398 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 20622 13268 20628 13320
rect 20680 13308 20686 13320
rect 21376 13308 21404 13339
rect 21818 13336 21824 13348
rect 21876 13336 21882 13388
rect 22462 13308 22468 13320
rect 20680 13280 21404 13308
rect 22423 13280 22468 13308
rect 20680 13268 20686 13280
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 24305 13311 24363 13317
rect 24305 13277 24317 13311
rect 24351 13277 24363 13311
rect 24578 13308 24584 13320
rect 24539 13280 24584 13308
rect 24305 13271 24363 13277
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 21174 13240 21180 13252
rect 16448 13212 21180 13240
rect 16448 13200 16454 13212
rect 21174 13200 21180 13212
rect 21232 13200 21238 13252
rect 24320 13240 24348 13271
rect 24578 13268 24584 13280
rect 24636 13268 24642 13320
rect 25130 13240 25136 13252
rect 24320 13212 25136 13240
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 12584 13144 13093 13172
rect 12584 13132 12590 13144
rect 13081 13141 13093 13144
rect 13127 13141 13139 13175
rect 13446 13172 13452 13184
rect 13407 13144 13452 13172
rect 13081 13135 13139 13141
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 14826 13172 14832 13184
rect 14787 13144 14832 13172
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 16114 13172 16120 13184
rect 16075 13144 16120 13172
rect 16114 13132 16120 13144
rect 16172 13132 16178 13184
rect 16482 13172 16488 13184
rect 16443 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 21910 13172 21916 13184
rect 21871 13144 21916 13172
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 11848 12940 12633 12968
rect 11848 12928 11854 12940
rect 12621 12937 12633 12940
rect 12667 12968 12679 12971
rect 13906 12968 13912 12980
rect 12667 12940 13912 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 13906 12928 13912 12940
rect 13964 12968 13970 12980
rect 14553 12971 14611 12977
rect 14553 12968 14565 12971
rect 13964 12940 14565 12968
rect 13964 12928 13970 12940
rect 14553 12937 14565 12940
rect 14599 12937 14611 12971
rect 15654 12968 15660 12980
rect 15615 12940 15660 12968
rect 14553 12931 14611 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12968 16727 12971
rect 16850 12968 16856 12980
rect 16715 12940 16856 12968
rect 16715 12937 16727 12940
rect 16669 12931 16727 12937
rect 16850 12928 16856 12940
rect 16908 12968 16914 12980
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 16908 12940 17417 12968
rect 16908 12928 16914 12940
rect 17405 12937 17417 12940
rect 17451 12937 17463 12971
rect 17405 12931 17463 12937
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 19153 12971 19211 12977
rect 19153 12968 19165 12971
rect 18932 12940 19165 12968
rect 18932 12928 18938 12940
rect 19153 12937 19165 12940
rect 19199 12937 19211 12971
rect 19153 12931 19211 12937
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 22830 12968 22836 12980
rect 22787 12940 22836 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 12161 12903 12219 12909
rect 12161 12869 12173 12903
rect 12207 12900 12219 12903
rect 12250 12900 12256 12912
rect 12207 12872 12256 12900
rect 12207 12869 12219 12872
rect 12161 12863 12219 12869
rect 12250 12860 12256 12872
rect 12308 12860 12314 12912
rect 12802 12860 12808 12912
rect 12860 12900 12866 12912
rect 12860 12872 13952 12900
rect 12860 12860 12866 12872
rect 13924 12844 13952 12872
rect 16114 12860 16120 12912
rect 16172 12909 16178 12912
rect 16172 12903 16221 12909
rect 16172 12869 16175 12903
rect 16209 12869 16221 12903
rect 16172 12863 16221 12869
rect 16301 12903 16359 12909
rect 16301 12869 16313 12903
rect 16347 12900 16359 12903
rect 16482 12900 16488 12912
rect 16347 12872 16488 12900
rect 16347 12869 16359 12872
rect 16301 12863 16359 12869
rect 16172 12860 16178 12863
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 19058 12860 19064 12912
rect 19116 12900 19122 12912
rect 19521 12903 19579 12909
rect 19521 12900 19533 12903
rect 19116 12872 19533 12900
rect 19116 12860 19122 12872
rect 19521 12869 19533 12872
rect 19567 12900 19579 12903
rect 25406 12900 25412 12912
rect 19567 12872 25412 12900
rect 19567 12869 19579 12872
rect 19521 12863 19579 12869
rect 25406 12860 25412 12872
rect 25464 12860 25470 12912
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 13446 12832 13452 12844
rect 11379 12804 13452 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 13446 12792 13452 12804
rect 13504 12832 13510 12844
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13504 12804 13645 12832
rect 13504 12792 13510 12804
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13906 12832 13912 12844
rect 13819 12804 13912 12832
rect 13633 12795 13691 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 16393 12835 16451 12841
rect 16393 12801 16405 12835
rect 16439 12832 16451 12835
rect 16574 12832 16580 12844
rect 16439 12804 16580 12832
rect 16439 12801 16451 12804
rect 16393 12795 16451 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 21039 12804 21833 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 21821 12801 21833 12804
rect 21867 12832 21879 12835
rect 21910 12832 21916 12844
rect 21867 12804 21916 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24670 12832 24676 12844
rect 24443 12804 24676 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24670 12792 24676 12804
rect 24728 12792 24734 12844
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12032 12736 12449 12764
rect 12032 12724 12038 12736
rect 12437 12733 12449 12736
rect 12483 12764 12495 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12483 12736 12909 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 13354 12764 13360 12776
rect 12943 12736 13360 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 14734 12724 14740 12776
rect 14792 12764 14798 12776
rect 15289 12767 15347 12773
rect 15289 12764 15301 12767
rect 14792 12736 15301 12764
rect 14792 12724 14798 12736
rect 15289 12733 15301 12736
rect 15335 12764 15347 12767
rect 16025 12767 16083 12773
rect 16025 12764 16037 12767
rect 15335 12736 16037 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 16025 12733 16037 12736
rect 16071 12733 16083 12767
rect 16025 12727 16083 12733
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18141 12767 18199 12773
rect 18141 12764 18153 12767
rect 18012 12736 18153 12764
rect 18012 12724 18018 12736
rect 18141 12733 18153 12736
rect 18187 12733 18199 12767
rect 20257 12767 20315 12773
rect 20257 12764 20269 12767
rect 18141 12727 18199 12733
rect 20088 12736 20269 12764
rect 13725 12699 13783 12705
rect 13725 12665 13737 12699
rect 13771 12665 13783 12699
rect 13725 12659 13783 12665
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11882 12628 11888 12640
rect 11287 12600 11888 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 13354 12628 13360 12640
rect 13315 12600 13360 12628
rect 13354 12588 13360 12600
rect 13412 12628 13418 12640
rect 13740 12628 13768 12659
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 20088 12705 20116 12736
rect 20257 12733 20269 12736
rect 20303 12764 20315 12767
rect 20346 12764 20352 12776
rect 20303 12736 20352 12764
rect 20303 12733 20315 12736
rect 20257 12727 20315 12733
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 20714 12764 20720 12776
rect 20675 12736 20720 12764
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 22830 12724 22836 12776
rect 22888 12764 22894 12776
rect 23477 12767 23535 12773
rect 23477 12764 23489 12767
rect 22888 12736 23489 12764
rect 22888 12724 22894 12736
rect 23477 12733 23489 12736
rect 23523 12764 23535 12767
rect 23753 12767 23811 12773
rect 23753 12764 23765 12767
rect 23523 12736 23765 12764
rect 23523 12733 23535 12736
rect 23477 12727 23535 12733
rect 23753 12733 23765 12736
rect 23799 12733 23811 12767
rect 23753 12727 23811 12733
rect 20073 12699 20131 12705
rect 20073 12696 20085 12699
rect 16724 12668 20085 12696
rect 16724 12656 16730 12668
rect 20073 12665 20085 12668
rect 20119 12665 20131 12699
rect 20364 12696 20392 12724
rect 21269 12699 21327 12705
rect 21269 12696 21281 12699
rect 20364 12668 21281 12696
rect 20073 12659 20131 12665
rect 21269 12665 21281 12668
rect 21315 12665 21327 12699
rect 21269 12659 21327 12665
rect 22142 12699 22200 12705
rect 22142 12665 22154 12699
rect 22188 12665 22200 12699
rect 22142 12659 22200 12665
rect 15010 12628 15016 12640
rect 13412 12600 13768 12628
rect 14971 12600 15016 12628
rect 13412 12588 13418 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 17037 12631 17095 12637
rect 17037 12628 17049 12631
rect 16632 12600 17049 12628
rect 16632 12588 16638 12600
rect 17037 12597 17049 12600
rect 17083 12597 17095 12631
rect 17037 12591 17095 12597
rect 17865 12631 17923 12637
rect 17865 12597 17877 12631
rect 17911 12628 17923 12631
rect 17954 12628 17960 12640
rect 17911 12600 17960 12628
rect 17911 12597 17923 12600
rect 17865 12591 17923 12597
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 18509 12631 18567 12637
rect 18509 12597 18521 12631
rect 18555 12628 18567 12631
rect 18598 12628 18604 12640
rect 18555 12600 18604 12628
rect 18555 12597 18567 12600
rect 18509 12591 18567 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 21634 12628 21640 12640
rect 21595 12600 21640 12628
rect 21634 12588 21640 12600
rect 21692 12628 21698 12640
rect 22157 12628 22185 12659
rect 22738 12628 22744 12640
rect 21692 12600 22744 12628
rect 21692 12588 21698 12600
rect 22738 12588 22744 12600
rect 22796 12628 22802 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 22796 12600 23029 12628
rect 22796 12588 22802 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 25130 12628 25136 12640
rect 25091 12600 25136 12628
rect 23017 12591 23075 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 14734 12424 14740 12436
rect 14695 12396 14740 12424
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 15010 12384 15016 12436
rect 15068 12424 15074 12436
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 15068 12396 15945 12424
rect 15068 12384 15074 12396
rect 15933 12393 15945 12396
rect 15979 12393 15991 12427
rect 16666 12424 16672 12436
rect 16627 12396 16672 12424
rect 15933 12387 15991 12393
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17313 12427 17371 12433
rect 17313 12393 17325 12427
rect 17359 12393 17371 12427
rect 17313 12387 17371 12393
rect 12526 12356 12532 12368
rect 12487 12328 12532 12356
rect 12526 12316 12532 12328
rect 12584 12316 12590 12368
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 13541 12359 13599 12365
rect 13541 12356 13553 12359
rect 13504 12328 13553 12356
rect 13504 12316 13510 12328
rect 13541 12325 13553 12328
rect 13587 12325 13599 12359
rect 13541 12319 13599 12325
rect 15289 12359 15347 12365
rect 15289 12325 15301 12359
rect 15335 12356 15347 12359
rect 15562 12356 15568 12368
rect 15335 12328 15568 12356
rect 15335 12325 15347 12328
rect 15289 12319 15347 12325
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16393 12359 16451 12365
rect 16393 12325 16405 12359
rect 16439 12356 16451 12359
rect 16482 12356 16488 12368
rect 16439 12328 16488 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 16482 12316 16488 12328
rect 16540 12356 16546 12368
rect 17328 12356 17356 12387
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 18785 12427 18843 12433
rect 18785 12424 18797 12427
rect 17552 12396 18797 12424
rect 17552 12384 17558 12396
rect 18785 12393 18797 12396
rect 18831 12393 18843 12427
rect 18785 12387 18843 12393
rect 25222 12384 25228 12436
rect 25280 12424 25286 12436
rect 25547 12427 25605 12433
rect 25547 12424 25559 12427
rect 25280 12396 25559 12424
rect 25280 12384 25286 12396
rect 25547 12393 25559 12396
rect 25593 12393 25605 12427
rect 25547 12387 25605 12393
rect 18690 12356 18696 12368
rect 16540 12328 18696 12356
rect 16540 12316 16546 12328
rect 18690 12316 18696 12328
rect 18748 12316 18754 12368
rect 21729 12359 21787 12365
rect 21729 12325 21741 12359
rect 21775 12356 21787 12359
rect 22462 12356 22468 12368
rect 21775 12328 22468 12356
rect 21775 12325 21787 12328
rect 21729 12319 21787 12325
rect 22462 12316 22468 12328
rect 22520 12316 22526 12368
rect 27614 12356 27620 12368
rect 25491 12328 27620 12356
rect 25491 12300 25519 12328
rect 27614 12316 27620 12328
rect 27672 12316 27678 12368
rect 11790 12288 11796 12300
rect 11751 12260 11796 12288
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 12345 12291 12403 12297
rect 12345 12288 12357 12291
rect 11940 12260 12357 12288
rect 11940 12248 11946 12260
rect 12345 12257 12357 12260
rect 12391 12288 12403 12291
rect 12618 12288 12624 12300
rect 12391 12260 12624 12288
rect 12391 12257 12403 12260
rect 12345 12251 12403 12257
rect 12618 12248 12624 12260
rect 12676 12288 12682 12300
rect 13078 12288 13084 12300
rect 12676 12260 13084 12288
rect 12676 12248 12682 12260
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 16724 12260 17141 12288
rect 16724 12248 16730 12260
rect 17129 12257 17141 12260
rect 17175 12288 17187 12291
rect 17589 12291 17647 12297
rect 17589 12288 17601 12291
rect 17175 12260 17601 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17589 12257 17601 12260
rect 17635 12257 17647 12291
rect 18138 12288 18144 12300
rect 18099 12260 18144 12288
rect 17589 12251 17647 12257
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13188 12192 13461 12220
rect 12802 12084 12808 12096
rect 12763 12056 12808 12084
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13188 12093 13216 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13906 12220 13912 12232
rect 13867 12192 13912 12220
rect 13449 12183 13507 12189
rect 13906 12180 13912 12192
rect 13964 12180 13970 12232
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12220 15163 12223
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15151 12192 15669 12220
rect 15151 12189 15163 12192
rect 15105 12183 15163 12189
rect 15657 12189 15669 12192
rect 15703 12220 15715 12223
rect 16574 12220 16580 12232
rect 15703 12192 16580 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 17604 12220 17632 12251
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 18371 12291 18429 12297
rect 18371 12257 18383 12291
rect 18417 12288 18429 12291
rect 19058 12288 19064 12300
rect 18417 12260 19064 12288
rect 18417 12257 18429 12260
rect 18371 12251 18429 12257
rect 18386 12220 18414 12251
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 21174 12288 21180 12300
rect 21135 12260 21180 12288
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 21453 12291 21511 12297
rect 21453 12257 21465 12291
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 24489 12291 24547 12297
rect 24489 12257 24501 12291
rect 24535 12288 24547 12291
rect 24762 12288 24768 12300
rect 24535 12260 24768 12288
rect 24535 12257 24547 12260
rect 24489 12251 24547 12257
rect 17604 12192 18414 12220
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 18598 12220 18604 12232
rect 18555 12192 18604 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 21468 12220 21496 12251
rect 24762 12248 24768 12260
rect 24820 12248 24826 12300
rect 25491 12297 25504 12300
rect 25476 12291 25504 12297
rect 25476 12288 25488 12291
rect 25411 12260 25488 12288
rect 25476 12257 25488 12260
rect 25476 12251 25504 12257
rect 25498 12248 25504 12251
rect 25556 12248 25562 12300
rect 20732 12192 21496 12220
rect 20732 12164 20760 12192
rect 16850 12112 16856 12164
rect 16908 12152 16914 12164
rect 20257 12155 20315 12161
rect 20257 12152 20269 12155
rect 16908 12124 20269 12152
rect 16908 12112 16914 12124
rect 20257 12121 20269 12124
rect 20303 12152 20315 12155
rect 20714 12152 20720 12164
rect 20303 12124 20720 12152
rect 20303 12121 20315 12124
rect 20257 12115 20315 12121
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 13173 12087 13231 12093
rect 13173 12084 13185 12087
rect 13044 12056 13185 12084
rect 13044 12044 13050 12056
rect 13173 12053 13185 12056
rect 13219 12053 13231 12087
rect 13173 12047 13231 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15427 12087 15485 12093
rect 15427 12084 15439 12087
rect 14792 12056 15439 12084
rect 14792 12044 14798 12056
rect 15427 12053 15439 12056
rect 15473 12053 15485 12087
rect 15427 12047 15485 12053
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 15654 12084 15660 12096
rect 15611 12056 15660 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 18046 12084 18052 12096
rect 17959 12056 18052 12084
rect 18046 12044 18052 12056
rect 18104 12084 18110 12096
rect 18279 12087 18337 12093
rect 18279 12084 18291 12087
rect 18104 12056 18291 12084
rect 18104 12044 18110 12056
rect 18279 12053 18291 12056
rect 18325 12053 18337 12087
rect 19150 12084 19156 12096
rect 19111 12056 19156 12084
rect 18279 12047 18337 12053
rect 19150 12044 19156 12056
rect 19208 12044 19214 12096
rect 20622 12084 20628 12096
rect 20583 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 24118 12084 24124 12096
rect 24079 12056 24124 12084
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 11790 11880 11796 11892
rect 11751 11852 11796 11880
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 14807 11840 14813 11892
rect 14865 11880 14871 11892
rect 16482 11880 16488 11892
rect 14865 11852 14910 11880
rect 16443 11852 16488 11880
rect 14865 11840 14871 11852
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 16850 11880 16856 11892
rect 16811 11852 16856 11880
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 18506 11880 18512 11892
rect 18467 11852 18512 11880
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 19058 11880 19064 11892
rect 19019 11852 19064 11880
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 21174 11840 21180 11892
rect 21232 11880 21238 11892
rect 21545 11883 21603 11889
rect 21545 11880 21557 11883
rect 21232 11852 21557 11880
rect 21232 11840 21238 11852
rect 21545 11849 21557 11852
rect 21591 11849 21603 11883
rect 24118 11880 24124 11892
rect 24079 11852 24124 11880
rect 21545 11843 21603 11849
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 25498 11880 25504 11892
rect 25459 11852 25504 11880
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 13446 11812 13452 11824
rect 10888 11784 13452 11812
rect 10888 11685 10916 11784
rect 13446 11772 13452 11784
rect 13504 11812 13510 11824
rect 13541 11815 13599 11821
rect 13541 11812 13553 11815
rect 13504 11784 13553 11812
rect 13504 11772 13510 11784
rect 13541 11781 13553 11784
rect 13587 11781 13599 11815
rect 13541 11775 13599 11781
rect 14553 11815 14611 11821
rect 14553 11781 14565 11815
rect 14599 11812 14611 11815
rect 14921 11815 14979 11821
rect 14921 11812 14933 11815
rect 14599 11784 14933 11812
rect 14599 11781 14611 11784
rect 14553 11775 14611 11781
rect 14921 11781 14933 11784
rect 14967 11812 14979 11815
rect 15378 11812 15384 11824
rect 14967 11784 15384 11812
rect 14967 11781 14979 11784
rect 14921 11775 14979 11781
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 18325 11815 18383 11821
rect 18325 11812 18337 11815
rect 17828 11784 18337 11812
rect 17828 11772 17834 11784
rect 18325 11781 18337 11784
rect 18371 11781 18383 11815
rect 18325 11775 18383 11781
rect 18598 11772 18604 11824
rect 18656 11812 18662 11824
rect 19429 11815 19487 11821
rect 19429 11812 19441 11815
rect 18656 11784 19441 11812
rect 18656 11772 18662 11784
rect 19429 11781 19441 11784
rect 19475 11781 19487 11815
rect 19429 11775 19487 11781
rect 11517 11747 11575 11753
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 13354 11744 13360 11756
rect 11563 11716 13360 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 14185 11747 14243 11753
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14231 11716 15025 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 15013 11713 15025 11716
rect 15059 11744 15071 11747
rect 16574 11744 16580 11756
rect 15059 11716 16580 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 18414 11744 18420 11756
rect 18327 11716 18420 11744
rect 18414 11704 18420 11716
rect 18472 11744 18478 11756
rect 19797 11747 19855 11753
rect 19797 11744 19809 11747
rect 18472 11716 19809 11744
rect 18472 11704 18478 11716
rect 19797 11713 19809 11716
rect 19843 11713 19855 11747
rect 19797 11707 19855 11713
rect 22186 11704 22192 11756
rect 22244 11744 22250 11756
rect 24581 11747 24639 11753
rect 24581 11744 24593 11747
rect 22244 11716 24593 11744
rect 22244 11704 22250 11716
rect 24581 11713 24593 11716
rect 24627 11744 24639 11747
rect 24946 11744 24952 11756
rect 24627 11716 24952 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 10689 11679 10747 11685
rect 10689 11645 10701 11679
rect 10735 11676 10747 11679
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10735 11648 10885 11676
rect 10735 11645 10747 11648
rect 10689 11639 10747 11645
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11676 12679 11679
rect 12802 11676 12808 11688
rect 12667 11648 12808 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 12802 11636 12808 11648
rect 12860 11676 12866 11688
rect 13630 11676 13636 11688
rect 12860 11648 13636 11676
rect 12860 11636 12866 11648
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 13786 11648 15393 11676
rect 12942 11611 13000 11617
rect 12942 11608 12954 11611
rect 12544 11580 12954 11608
rect 12544 11552 12572 11580
rect 12942 11577 12954 11580
rect 12988 11577 13000 11611
rect 12942 11571 13000 11577
rect 13078 11568 13084 11620
rect 13136 11608 13142 11620
rect 13786 11608 13814 11648
rect 15381 11645 15393 11648
rect 15427 11645 15439 11679
rect 15381 11639 15439 11645
rect 16356 11679 16414 11685
rect 16356 11645 16368 11679
rect 16402 11645 16414 11679
rect 16356 11639 16414 11645
rect 14642 11608 14648 11620
rect 13136 11580 13814 11608
rect 14603 11580 14648 11608
rect 13136 11568 13142 11580
rect 14642 11568 14648 11580
rect 14700 11568 14706 11620
rect 15562 11568 15568 11620
rect 15620 11608 15626 11620
rect 16209 11611 16267 11617
rect 16209 11608 16221 11611
rect 15620 11580 16221 11608
rect 15620 11568 15626 11580
rect 16209 11577 16221 11580
rect 16255 11577 16267 11611
rect 16209 11571 16267 11577
rect 12158 11500 12164 11552
rect 12216 11540 12222 11552
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 12216 11512 12265 11540
rect 12216 11500 12222 11512
rect 12253 11509 12265 11512
rect 12299 11540 12311 11543
rect 12526 11540 12532 11552
rect 12299 11512 12532 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15654 11540 15660 11552
rect 15436 11512 15660 11540
rect 15436 11500 15442 11512
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16114 11540 16120 11552
rect 16075 11512 16120 11540
rect 16114 11500 16120 11512
rect 16172 11540 16178 11552
rect 16371 11540 16399 11639
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18196 11679 18254 11685
rect 18196 11676 18208 11679
rect 17920 11648 18208 11676
rect 17920 11636 17926 11648
rect 18196 11645 18208 11648
rect 18242 11676 18254 11679
rect 19150 11676 19156 11688
rect 18242 11648 19156 11676
rect 18242 11645 18254 11648
rect 18196 11639 18254 11645
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 20346 11636 20352 11688
rect 20404 11676 20410 11688
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 20404 11648 20545 11676
rect 20404 11636 20410 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20772 11648 21005 11676
rect 20772 11636 20778 11648
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 17497 11611 17555 11617
rect 17497 11577 17509 11611
rect 17543 11608 17555 11611
rect 18049 11611 18107 11617
rect 18049 11608 18061 11611
rect 17543 11580 18061 11608
rect 17543 11577 17555 11580
rect 17497 11571 17555 11577
rect 18049 11577 18061 11580
rect 18095 11577 18107 11611
rect 21266 11608 21272 11620
rect 21227 11580 21272 11608
rect 18049 11571 18107 11577
rect 17770 11540 17776 11552
rect 16172 11512 16399 11540
rect 17731 11512 17776 11540
rect 16172 11500 16178 11512
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 18064 11540 18092 11571
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 22557 11611 22615 11617
rect 22557 11577 22569 11611
rect 22603 11608 22615 11611
rect 24302 11608 24308 11620
rect 22603 11580 24308 11608
rect 22603 11577 22615 11580
rect 22557 11571 22615 11577
rect 24302 11568 24308 11580
rect 24360 11568 24366 11620
rect 24397 11611 24455 11617
rect 24397 11577 24409 11611
rect 24443 11577 24455 11611
rect 24397 11571 24455 11577
rect 18138 11540 18144 11552
rect 18064 11512 18144 11540
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 23382 11540 23388 11552
rect 23343 11512 23388 11540
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 24118 11500 24124 11552
rect 24176 11540 24182 11552
rect 24412 11540 24440 11571
rect 24176 11512 24440 11540
rect 24176 11500 24182 11512
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 11885 11339 11943 11345
rect 11885 11305 11897 11339
rect 11931 11336 11943 11339
rect 13078 11336 13084 11348
rect 11931 11308 13084 11336
rect 11931 11305 11943 11308
rect 11885 11299 11943 11305
rect 13078 11296 13084 11308
rect 13136 11296 13142 11348
rect 13446 11336 13452 11348
rect 13407 11308 13452 11336
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14734 11336 14740 11348
rect 14695 11308 14740 11336
rect 14734 11296 14740 11308
rect 14792 11336 14798 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 14792 11308 15761 11336
rect 14792 11296 14798 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 15749 11299 15807 11305
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 21085 11339 21143 11345
rect 21085 11336 21097 11339
rect 20864 11308 21097 11336
rect 20864 11296 20870 11308
rect 21085 11305 21097 11308
rect 21131 11305 21143 11339
rect 21634 11336 21640 11348
rect 21595 11308 21640 11336
rect 21085 11299 21143 11305
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22189 11339 22247 11345
rect 22189 11305 22201 11339
rect 22235 11336 22247 11339
rect 23014 11336 23020 11348
rect 22235 11308 23020 11336
rect 22235 11305 22247 11308
rect 22189 11299 22247 11305
rect 23014 11296 23020 11308
rect 23072 11336 23078 11348
rect 24302 11336 24308 11348
rect 23072 11308 23244 11336
rect 24263 11308 24308 11336
rect 23072 11296 23078 11308
rect 12161 11271 12219 11277
rect 12161 11237 12173 11271
rect 12207 11268 12219 11271
rect 12250 11268 12256 11280
rect 12207 11240 12256 11268
rect 12207 11237 12219 11240
rect 12161 11231 12219 11237
rect 12250 11228 12256 11240
rect 12308 11228 12314 11280
rect 12342 11228 12348 11280
rect 12400 11268 12406 11280
rect 15105 11271 15163 11277
rect 12400 11240 13584 11268
rect 12400 11228 12406 11240
rect 1302 11160 1308 11212
rect 1360 11200 1366 11212
rect 13556 11209 13584 11240
rect 15105 11237 15117 11271
rect 15151 11268 15163 11271
rect 15562 11268 15568 11280
rect 15151 11240 15568 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15562 11228 15568 11240
rect 15620 11268 15626 11280
rect 16209 11271 16267 11277
rect 16209 11268 16221 11271
rect 15620 11240 16221 11268
rect 15620 11228 15626 11240
rect 16209 11237 16221 11240
rect 16255 11237 16267 11271
rect 16209 11231 16267 11237
rect 19061 11271 19119 11277
rect 19061 11237 19073 11271
rect 19107 11268 19119 11271
rect 20622 11268 20628 11280
rect 19107 11240 20628 11268
rect 19107 11237 19119 11240
rect 19061 11231 19119 11237
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 23106 11268 23112 11280
rect 23067 11240 23112 11268
rect 23106 11228 23112 11240
rect 23164 11228 23170 11280
rect 23216 11277 23244 11308
rect 24302 11296 24308 11308
rect 24360 11296 24366 11348
rect 23201 11271 23259 11277
rect 23201 11237 23213 11271
rect 23247 11237 23259 11271
rect 24762 11268 24768 11280
rect 24723 11240 24768 11268
rect 23201 11231 23259 11237
rect 24762 11228 24768 11240
rect 24820 11228 24826 11280
rect 1432 11203 1490 11209
rect 1432 11200 1444 11203
rect 1360 11172 1444 11200
rect 1360 11160 1366 11172
rect 1432 11169 1444 11172
rect 1478 11169 1490 11203
rect 1432 11163 1490 11169
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 13630 11200 13636 11212
rect 13587 11172 13636 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 14090 11200 14096 11212
rect 13786 11172 14096 11200
rect 13786 11144 13814 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 16022 11200 16028 11212
rect 15335 11172 16028 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 16022 11160 16028 11172
rect 16080 11200 16086 11212
rect 16853 11203 16911 11209
rect 16853 11200 16865 11203
rect 16080 11172 16865 11200
rect 16080 11160 16086 11172
rect 16853 11169 16865 11172
rect 16899 11169 16911 11203
rect 18322 11200 18328 11212
rect 18283 11172 18328 11200
rect 16853 11163 16911 11169
rect 18322 11160 18328 11172
rect 18380 11160 18386 11212
rect 12066 11132 12072 11144
rect 4126 11104 12072 11132
rect 1535 10999 1593 11005
rect 1535 10965 1547 10999
rect 1581 10996 1593 10999
rect 4126 10996 4154 11104
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11132 12771 11135
rect 12986 11132 12992 11144
rect 12759 11104 12992 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13722 11092 13728 11144
rect 13780 11104 13814 11144
rect 13780 11092 13786 11104
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16761 11135 16819 11141
rect 16761 11132 16773 11135
rect 16724 11104 16773 11132
rect 16724 11092 16730 11104
rect 16761 11101 16773 11104
rect 16807 11101 16819 11135
rect 16761 11095 16819 11101
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 18012 11104 18705 11132
rect 18012 11092 18018 11104
rect 18693 11101 18705 11104
rect 18739 11132 18751 11135
rect 19150 11132 19156 11144
rect 18739 11104 19156 11132
rect 18739 11101 18751 11104
rect 18693 11095 18751 11101
rect 19150 11092 19156 11104
rect 19208 11092 19214 11144
rect 21266 11132 21272 11144
rect 21227 11104 21272 11132
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11132 23811 11135
rect 24026 11132 24032 11144
rect 23799 11104 24032 11132
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 24026 11092 24032 11104
rect 24084 11132 24090 11144
rect 24673 11135 24731 11141
rect 24673 11132 24685 11135
rect 24084 11104 24685 11132
rect 24084 11092 24090 11104
rect 24673 11101 24685 11104
rect 24719 11101 24731 11135
rect 24946 11132 24952 11144
rect 24907 11104 24952 11132
rect 24673 11095 24731 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 18463 11067 18521 11073
rect 18463 11064 18475 11067
rect 17880 11036 18475 11064
rect 17880 11008 17908 11036
rect 18463 11033 18475 11036
rect 18509 11033 18521 11067
rect 18463 11027 18521 11033
rect 1581 10968 4154 10996
rect 1581 10965 1593 10968
rect 1535 10959 1593 10965
rect 15378 10956 15384 11008
rect 15436 10996 15442 11008
rect 15473 10999 15531 11005
rect 15473 10996 15485 10999
rect 15436 10968 15485 10996
rect 15436 10956 15442 10968
rect 15473 10965 15485 10968
rect 15519 10965 15531 10999
rect 15473 10959 15531 10965
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 16669 10999 16727 11005
rect 16669 10996 16681 10999
rect 16632 10968 16681 10996
rect 16632 10956 16638 10968
rect 16669 10965 16681 10968
rect 16715 10996 16727 10999
rect 17126 10996 17132 11008
rect 16715 10968 17132 10996
rect 16715 10965 16727 10968
rect 16669 10959 16727 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17862 10996 17868 11008
rect 17823 10968 17868 10996
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 18138 10996 18144 11008
rect 18099 10968 18144 10996
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 18601 10999 18659 11005
rect 18601 10965 18613 10999
rect 18647 10996 18659 10999
rect 18690 10996 18696 11008
rect 18647 10968 18696 10996
rect 18647 10965 18659 10968
rect 18601 10959 18659 10965
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 20625 10999 20683 11005
rect 20625 10965 20637 10999
rect 20671 10996 20683 10999
rect 20714 10996 20720 11008
rect 20671 10968 20720 10996
rect 20671 10965 20683 10968
rect 20625 10959 20683 10965
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1302 10752 1308 10804
rect 1360 10792 1366 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1360 10764 1593 10792
rect 1360 10752 1366 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 13630 10792 13636 10804
rect 13591 10764 13636 10792
rect 1581 10755 1639 10761
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 14148 10764 15485 10792
rect 14148 10752 14154 10764
rect 15473 10761 15485 10764
rect 15519 10761 15531 10795
rect 15473 10755 15531 10761
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 17770 10792 17776 10804
rect 17727 10764 17776 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 17770 10752 17776 10764
rect 17828 10792 17834 10804
rect 18325 10795 18383 10801
rect 18325 10792 18337 10795
rect 17828 10764 18337 10792
rect 17828 10752 17834 10764
rect 18325 10761 18337 10764
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 18693 10795 18751 10801
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 18782 10792 18788 10804
rect 18739 10764 18788 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 23014 10792 23020 10804
rect 22975 10764 23020 10792
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 24762 10792 24768 10804
rect 23446 10764 24768 10792
rect 23446 10736 23474 10764
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 10689 10727 10747 10733
rect 10689 10693 10701 10727
rect 10735 10724 10747 10727
rect 11790 10724 11796 10736
rect 10735 10696 11796 10724
rect 10735 10693 10747 10696
rect 10689 10687 10747 10693
rect 10796 10597 10824 10696
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 12253 10727 12311 10733
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12526 10724 12532 10736
rect 12299 10696 12532 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 15151 10727 15209 10733
rect 15151 10724 15163 10727
rect 14792 10696 15163 10724
rect 14792 10684 14798 10696
rect 15151 10693 15163 10696
rect 15197 10693 15209 10727
rect 15151 10687 15209 10693
rect 15289 10727 15347 10733
rect 15289 10693 15301 10727
rect 15335 10724 15347 10727
rect 16482 10724 16488 10736
rect 15335 10696 16488 10724
rect 15335 10693 15347 10696
rect 15289 10687 15347 10693
rect 15488 10668 15516 10696
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 17126 10724 17132 10736
rect 17039 10696 17132 10724
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 17862 10684 17868 10736
rect 17920 10724 17926 10736
rect 18187 10727 18245 10733
rect 18187 10724 18199 10727
rect 17920 10696 18199 10724
rect 17920 10684 17926 10696
rect 18187 10693 18199 10696
rect 18233 10693 18245 10727
rect 18187 10687 18245 10693
rect 22741 10727 22799 10733
rect 22741 10693 22753 10727
rect 22787 10724 22799 10727
rect 23382 10724 23388 10736
rect 22787 10696 23388 10724
rect 22787 10693 22799 10696
rect 22741 10687 22799 10693
rect 23382 10684 23388 10696
rect 23440 10696 23474 10736
rect 25774 10724 25780 10736
rect 25735 10696 25780 10724
rect 23440 10684 23446 10696
rect 25774 10684 25780 10696
rect 25832 10684 25838 10736
rect 13722 10656 13728 10668
rect 11348 10628 13728 10656
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 11348 10597 11376 10628
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14884 10628 15393 10656
rect 14884 10616 14890 10628
rect 15381 10625 15393 10628
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 15470 10616 15476 10668
rect 15528 10616 15534 10668
rect 17144 10656 17172 10684
rect 18414 10656 18420 10668
rect 17144 10628 18420 10656
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 21174 10656 21180 10668
rect 20548 10628 21180 10656
rect 11333 10591 11391 10597
rect 11333 10588 11345 10591
rect 10928 10560 11345 10588
rect 10928 10548 10934 10560
rect 11333 10557 11345 10560
rect 11379 10557 11391 10591
rect 11333 10551 11391 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10588 11575 10591
rect 12434 10588 12440 10600
rect 11563 10560 12440 10588
rect 11563 10557 11575 10560
rect 11517 10551 11575 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 14366 10548 14372 10600
rect 14424 10588 14430 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 14424 10560 14565 10588
rect 14424 10548 14430 10560
rect 14553 10557 14565 10560
rect 14599 10588 14611 10591
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14599 10560 15025 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 15013 10557 15025 10560
rect 15059 10588 15071 10591
rect 15562 10588 15568 10600
rect 15059 10560 15568 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16850 10588 16856 10600
rect 16531 10560 16856 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 16850 10548 16856 10560
rect 16908 10588 16914 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16908 10560 16957 10588
rect 16908 10548 16914 10560
rect 16945 10557 16957 10560
rect 16991 10588 17003 10591
rect 18598 10588 18604 10600
rect 16991 10560 18604 10588
rect 16991 10557 17003 10560
rect 16945 10551 17003 10557
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 20438 10548 20444 10600
rect 20496 10588 20502 10600
rect 20548 10597 20576 10628
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 24026 10616 24032 10628
rect 24084 10656 24090 10668
rect 25041 10659 25099 10665
rect 25041 10656 25053 10659
rect 24084 10628 25053 10656
rect 24084 10616 24090 10628
rect 25041 10625 25053 10628
rect 25087 10625 25099 10659
rect 25041 10619 25099 10625
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 20496 10560 20545 10588
rect 20496 10548 20502 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 20714 10588 20720 10600
rect 20675 10560 20720 10588
rect 20533 10551 20591 10557
rect 20714 10548 20720 10560
rect 20772 10548 20778 10600
rect 20993 10591 21051 10597
rect 20993 10557 21005 10591
rect 21039 10588 21051 10591
rect 21818 10588 21824 10600
rect 21039 10560 21824 10588
rect 21039 10557 21051 10560
rect 20993 10551 21051 10557
rect 21818 10548 21824 10560
rect 21876 10548 21882 10600
rect 25292 10591 25350 10597
rect 25292 10557 25304 10591
rect 25338 10588 25350 10591
rect 25792 10588 25820 10684
rect 25338 10560 25820 10588
rect 25338 10557 25350 10560
rect 25292 10551 25350 10557
rect 11885 10523 11943 10529
rect 11885 10489 11897 10523
rect 11931 10520 11943 10523
rect 12250 10520 12256 10532
rect 11931 10492 12256 10520
rect 11931 10489 11943 10492
rect 11885 10483 11943 10489
rect 12250 10480 12256 10492
rect 12308 10520 12314 10532
rect 12308 10492 12474 10520
rect 12308 10480 12314 10492
rect 12446 10452 12474 10492
rect 12526 10480 12532 10532
rect 12584 10520 12590 10532
rect 12758 10523 12816 10529
rect 12758 10520 12770 10523
rect 12584 10492 12770 10520
rect 12584 10480 12590 10492
rect 12758 10489 12770 10492
rect 12804 10489 12816 10523
rect 12758 10483 12816 10489
rect 14185 10523 14243 10529
rect 14185 10489 14197 10523
rect 14231 10520 14243 10523
rect 15470 10520 15476 10532
rect 14231 10492 15476 10520
rect 14231 10489 14243 10492
rect 14185 10483 14243 10489
rect 15470 10480 15476 10492
rect 15528 10480 15534 10532
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 17497 10523 17555 10529
rect 17497 10520 17509 10523
rect 16632 10492 17509 10520
rect 16632 10480 16638 10492
rect 17497 10489 17509 10492
rect 17543 10520 17555 10523
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 17543 10492 18061 10520
rect 17543 10489 17555 10492
rect 17497 10483 17555 10489
rect 18049 10489 18061 10492
rect 18095 10520 18107 10523
rect 18322 10520 18328 10532
rect 18095 10492 18328 10520
rect 18095 10489 18107 10492
rect 18049 10483 18107 10489
rect 18322 10480 18328 10492
rect 18380 10520 18386 10532
rect 22142 10523 22200 10529
rect 18380 10492 19564 10520
rect 18380 10480 18386 10492
rect 19536 10464 19564 10492
rect 22142 10489 22154 10523
rect 22188 10489 22200 10523
rect 23750 10520 23756 10532
rect 23711 10492 23756 10520
rect 22142 10483 22200 10489
rect 13078 10452 13084 10464
rect 12446 10424 13084 10452
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 13357 10455 13415 10461
rect 13357 10452 13369 10455
rect 13136 10424 13369 10452
rect 13136 10412 13142 10424
rect 13357 10421 13369 10424
rect 13403 10421 13415 10455
rect 14826 10452 14832 10464
rect 14787 10424 14832 10452
rect 13357 10415 13415 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 16022 10452 16028 10464
rect 15983 10424 16028 10452
rect 16022 10412 16028 10424
rect 16080 10452 16086 10464
rect 16761 10455 16819 10461
rect 16761 10452 16773 10455
rect 16080 10424 16773 10452
rect 16080 10412 16086 10424
rect 16761 10421 16773 10424
rect 16807 10452 16819 10455
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 16807 10424 17693 10452
rect 16807 10421 16819 10424
rect 16761 10415 16819 10421
rect 17681 10421 17693 10424
rect 17727 10452 17739 10455
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 17727 10424 17785 10452
rect 17727 10421 17739 10424
rect 17681 10415 17739 10421
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 19150 10452 19156 10464
rect 19111 10424 19156 10452
rect 17773 10415 17831 10421
rect 19150 10412 19156 10424
rect 19208 10412 19214 10464
rect 19518 10452 19524 10464
rect 19479 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19889 10455 19947 10461
rect 19889 10421 19901 10455
rect 19935 10452 19947 10455
rect 19978 10452 19984 10464
rect 19935 10424 19984 10452
rect 19935 10421 19947 10424
rect 19889 10415 19947 10421
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 21174 10412 21180 10464
rect 21232 10452 21238 10464
rect 21269 10455 21327 10461
rect 21269 10452 21281 10455
rect 21232 10424 21281 10452
rect 21232 10412 21238 10424
rect 21269 10421 21281 10424
rect 21315 10452 21327 10455
rect 21634 10452 21640 10464
rect 21315 10424 21640 10452
rect 21315 10421 21327 10424
rect 21269 10415 21327 10421
rect 21634 10412 21640 10424
rect 21692 10452 21698 10464
rect 22157 10452 22185 10483
rect 23750 10480 23756 10492
rect 23808 10480 23814 10532
rect 23845 10523 23903 10529
rect 23845 10489 23857 10523
rect 23891 10489 23903 10523
rect 23845 10483 23903 10489
rect 23382 10452 23388 10464
rect 21692 10424 22185 10452
rect 23343 10424 23388 10452
rect 21692 10412 21698 10424
rect 23382 10412 23388 10424
rect 23440 10452 23446 10464
rect 23860 10452 23888 10483
rect 23440 10424 23888 10452
rect 23440 10412 23446 10424
rect 24762 10412 24768 10464
rect 24820 10452 24826 10464
rect 25363 10455 25421 10461
rect 25363 10452 25375 10455
rect 24820 10424 25375 10452
rect 24820 10412 24826 10424
rect 25363 10421 25375 10424
rect 25409 10421 25421 10455
rect 25363 10415 25421 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 10870 10248 10876 10260
rect 10831 10220 10876 10248
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12066 10248 12072 10260
rect 12027 10220 12072 10248
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 12434 10248 12440 10260
rect 12395 10220 12440 10248
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 13722 10248 13728 10260
rect 13683 10220 13728 10248
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14792 10220 15025 10248
rect 14792 10208 14798 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 16850 10248 16856 10260
rect 16811 10220 16856 10248
rect 15013 10211 15071 10217
rect 12802 10180 12808 10192
rect 12763 10152 12808 10180
rect 12802 10140 12808 10152
rect 12860 10140 12866 10192
rect 14185 10115 14243 10121
rect 14185 10081 14197 10115
rect 14231 10081 14243 10115
rect 14660 10112 14688 10208
rect 15028 10180 15056 10211
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17865 10251 17923 10257
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 18414 10248 18420 10260
rect 17911 10220 18420 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 18414 10208 18420 10220
rect 18472 10208 18478 10260
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 20438 10248 20444 10260
rect 20395 10220 20444 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 21876 10220 22293 10248
rect 21876 10208 21882 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 23106 10208 23112 10260
rect 23164 10248 23170 10260
rect 23569 10251 23627 10257
rect 23569 10248 23581 10251
rect 23164 10220 23581 10248
rect 23164 10208 23170 10220
rect 23569 10217 23581 10220
rect 23615 10217 23627 10251
rect 23569 10211 23627 10217
rect 24535 10251 24593 10257
rect 24535 10217 24547 10251
rect 24581 10248 24593 10251
rect 24854 10248 24860 10260
rect 24581 10220 24860 10248
rect 24581 10217 24593 10220
rect 24535 10211 24593 10217
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 19061 10183 19119 10189
rect 15028 10152 15479 10180
rect 15286 10112 15292 10124
rect 14660 10084 15292 10112
rect 14185 10075 14243 10081
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 12986 10044 12992 10056
rect 12947 10016 12992 10044
rect 12986 10004 12992 10016
rect 13044 10004 13050 10056
rect 14200 10044 14228 10075
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15451 10121 15479 10152
rect 19061 10149 19073 10183
rect 19107 10180 19119 10183
rect 20625 10183 20683 10189
rect 20625 10180 20637 10183
rect 19107 10152 20637 10180
rect 19107 10149 19119 10152
rect 19061 10143 19119 10149
rect 20625 10149 20637 10152
rect 20671 10180 20683 10183
rect 20714 10180 20720 10192
rect 20671 10152 20720 10180
rect 20671 10149 20683 10152
rect 20625 10143 20683 10149
rect 20714 10140 20720 10152
rect 20772 10140 20778 10192
rect 21266 10140 21272 10192
rect 21324 10180 21330 10192
rect 21913 10183 21971 10189
rect 21913 10180 21925 10183
rect 21324 10152 21925 10180
rect 21324 10140 21330 10152
rect 21913 10149 21925 10152
rect 21959 10149 21971 10183
rect 21913 10143 21971 10149
rect 23293 10183 23351 10189
rect 23293 10149 23305 10183
rect 23339 10180 23351 10183
rect 23382 10180 23388 10192
rect 23339 10152 23388 10180
rect 23339 10149 23351 10152
rect 23293 10143 23351 10149
rect 23382 10140 23388 10152
rect 23440 10140 23446 10192
rect 23750 10140 23756 10192
rect 23808 10180 23814 10192
rect 24029 10183 24087 10189
rect 24029 10180 24041 10183
rect 23808 10152 24041 10180
rect 23808 10140 23814 10152
rect 24029 10149 24041 10152
rect 24075 10180 24087 10183
rect 24762 10180 24768 10192
rect 24075 10152 24768 10180
rect 24075 10149 24087 10152
rect 24029 10143 24087 10149
rect 24762 10140 24768 10152
rect 24820 10140 24826 10192
rect 15436 10115 15494 10121
rect 15436 10081 15448 10115
rect 15482 10081 15494 10115
rect 15436 10075 15494 10081
rect 17313 10115 17371 10121
rect 17313 10081 17325 10115
rect 17359 10112 17371 10115
rect 17494 10112 17500 10124
rect 17359 10084 17500 10112
rect 17359 10081 17371 10084
rect 17313 10075 17371 10081
rect 17494 10072 17500 10084
rect 17552 10112 17558 10124
rect 18046 10112 18052 10124
rect 17552 10084 18052 10112
rect 17552 10072 17558 10084
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 18138 10072 18144 10124
rect 18196 10112 18202 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 18196 10084 18337 10112
rect 18196 10072 18202 10084
rect 18325 10081 18337 10084
rect 18371 10081 18383 10115
rect 18325 10075 18383 10081
rect 20346 10072 20352 10124
rect 20404 10112 20410 10124
rect 20898 10112 20904 10124
rect 20404 10084 20904 10112
rect 20404 10072 20410 10084
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 21358 10112 21364 10124
rect 21319 10084 21364 10112
rect 21358 10072 21364 10084
rect 21416 10072 21422 10124
rect 23014 10112 23020 10124
rect 22975 10084 23020 10112
rect 23014 10072 23020 10084
rect 23072 10072 23078 10124
rect 24464 10115 24522 10121
rect 24464 10081 24476 10115
rect 24510 10112 24522 10115
rect 24670 10112 24676 10124
rect 24510 10084 24676 10112
rect 24510 10081 24522 10084
rect 24464 10075 24522 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 25476 10115 25534 10121
rect 25476 10081 25488 10115
rect 25522 10112 25534 10115
rect 26142 10112 26148 10124
rect 25522 10084 26148 10112
rect 25522 10081 25534 10084
rect 25476 10075 25534 10081
rect 26142 10072 26148 10084
rect 26200 10072 26206 10124
rect 15657 10047 15715 10053
rect 14200 10016 14688 10044
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 14200 9908 14228 10016
rect 14660 9976 14688 10016
rect 15657 10013 15669 10047
rect 15703 10044 15715 10047
rect 15930 10044 15936 10056
rect 15703 10016 15936 10044
rect 15703 10013 15715 10016
rect 15657 10007 15715 10013
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 19150 10044 19156 10056
rect 18739 10016 19156 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 19150 10004 19156 10016
rect 19208 10004 19214 10056
rect 21450 10044 21456 10056
rect 21411 10016 21456 10044
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 16574 9976 16580 9988
rect 14660 9948 16580 9976
rect 16574 9936 16580 9948
rect 16632 9936 16638 9988
rect 17497 9979 17555 9985
rect 17497 9945 17509 9979
rect 17543 9976 17555 9979
rect 17862 9976 17868 9988
rect 17543 9948 17868 9976
rect 17543 9945 17555 9948
rect 17497 9939 17555 9945
rect 17862 9936 17868 9948
rect 17920 9976 17926 9988
rect 18490 9979 18548 9985
rect 18490 9976 18502 9979
rect 17920 9948 18502 9976
rect 17920 9936 17926 9948
rect 18490 9945 18502 9948
rect 18536 9976 18548 9979
rect 18536 9948 19288 9976
rect 18536 9945 18548 9948
rect 18490 9939 18548 9945
rect 19260 9920 19288 9948
rect 13780 9880 14228 9908
rect 13780 9868 13786 9880
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15565 9911 15623 9917
rect 15565 9908 15577 9911
rect 15528 9880 15577 9908
rect 15528 9868 15534 9880
rect 15565 9877 15577 9880
rect 15611 9877 15623 9911
rect 15746 9908 15752 9920
rect 15707 9880 15752 9908
rect 15565 9871 15623 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16485 9911 16543 9917
rect 16485 9877 16497 9911
rect 16531 9908 16543 9911
rect 16666 9908 16672 9920
rect 16531 9880 16672 9908
rect 16531 9877 16543 9880
rect 16485 9871 16543 9877
rect 16666 9868 16672 9880
rect 16724 9868 16730 9920
rect 18230 9908 18236 9920
rect 18191 9880 18236 9908
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18598 9908 18604 9920
rect 18559 9880 18604 9908
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 19337 9911 19395 9917
rect 19337 9908 19349 9911
rect 19300 9880 19349 9908
rect 19300 9868 19306 9880
rect 19337 9877 19349 9880
rect 19383 9877 19395 9911
rect 19337 9871 19395 9877
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25547 9911 25605 9917
rect 25547 9908 25559 9911
rect 25004 9880 25559 9908
rect 25004 9868 25010 9880
rect 25547 9877 25559 9880
rect 25593 9877 25605 9911
rect 25547 9871 25605 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 14369 9707 14427 9713
rect 14369 9673 14381 9707
rect 14415 9704 14427 9707
rect 14734 9704 14740 9716
rect 14415 9676 14740 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 14734 9664 14740 9676
rect 14792 9704 14798 9716
rect 14967 9707 15025 9713
rect 14967 9704 14979 9707
rect 14792 9676 14979 9704
rect 14792 9664 14798 9676
rect 14967 9673 14979 9676
rect 15013 9704 15025 9707
rect 15654 9704 15660 9716
rect 15013 9676 15660 9704
rect 15013 9673 15025 9676
rect 14967 9667 15025 9673
rect 15654 9664 15660 9676
rect 15712 9704 15718 9716
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 15712 9676 16221 9704
rect 15712 9664 15718 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 16209 9667 16267 9673
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 16853 9707 16911 9713
rect 16853 9704 16865 9707
rect 16356 9676 16865 9704
rect 16356 9664 16362 9676
rect 16853 9673 16865 9676
rect 16899 9673 16911 9707
rect 16853 9667 16911 9673
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 19613 9707 19671 9713
rect 19613 9704 19625 9707
rect 18656 9676 19625 9704
rect 18656 9664 18662 9676
rect 19613 9673 19625 9676
rect 19659 9704 19671 9707
rect 19978 9704 19984 9716
rect 19659 9676 19984 9704
rect 19659 9673 19671 9676
rect 19613 9667 19671 9673
rect 19978 9664 19984 9676
rect 20036 9664 20042 9716
rect 20438 9704 20444 9716
rect 20399 9676 20444 9704
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21637 9707 21695 9713
rect 21637 9704 21649 9707
rect 20956 9676 21649 9704
rect 20956 9664 20962 9676
rect 21637 9673 21649 9676
rect 21683 9673 21695 9707
rect 21637 9667 21695 9673
rect 22649 9707 22707 9713
rect 22649 9673 22661 9707
rect 22695 9704 22707 9707
rect 23014 9704 23020 9716
rect 22695 9676 23020 9704
rect 22695 9673 22707 9676
rect 22649 9667 22707 9673
rect 23014 9664 23020 9676
rect 23072 9664 23078 9716
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 25130 9664 25136 9716
rect 25188 9704 25194 9716
rect 25363 9707 25421 9713
rect 25363 9704 25375 9707
rect 25188 9676 25375 9704
rect 25188 9664 25194 9676
rect 25363 9673 25375 9676
rect 25409 9673 25421 9707
rect 26142 9704 26148 9716
rect 26103 9676 26148 9704
rect 25363 9667 25421 9673
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 9030 9596 9036 9648
rect 9088 9636 9094 9648
rect 13722 9636 13728 9648
rect 9088 9608 13728 9636
rect 9088 9596 9094 9608
rect 13722 9596 13728 9608
rect 13780 9636 13786 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13780 9608 13921 9636
rect 13780 9596 13786 9608
rect 13909 9605 13921 9608
rect 13955 9605 13967 9639
rect 13909 9599 13967 9605
rect 14826 9596 14832 9648
rect 14884 9596 14890 9648
rect 15105 9639 15163 9645
rect 15105 9605 15117 9639
rect 15151 9636 15163 9639
rect 15378 9636 15384 9648
rect 15151 9608 15384 9636
rect 15151 9605 15163 9608
rect 15105 9599 15163 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 16666 9636 16672 9648
rect 16627 9608 16672 9636
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 18230 9596 18236 9648
rect 18288 9636 18294 9648
rect 18417 9639 18475 9645
rect 18417 9636 18429 9639
rect 18288 9608 18429 9636
rect 18288 9596 18294 9608
rect 18417 9605 18429 9608
rect 18463 9636 18475 9639
rect 19334 9636 19340 9648
rect 18463 9608 19340 9636
rect 18463 9605 18475 9608
rect 18417 9599 18475 9605
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12860 9540 13185 9568
rect 12860 9528 12866 9540
rect 13173 9537 13185 9540
rect 13219 9568 13231 9571
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13219 9540 13461 9568
rect 13219 9537 13231 9540
rect 13173 9531 13231 9537
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 14844 9568 14872 9596
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14783 9540 15209 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15197 9537 15209 9540
rect 15243 9568 15255 9571
rect 15930 9568 15936 9580
rect 15243 9540 15936 9568
rect 15243 9537 15255 9540
rect 15197 9531 15255 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 16761 9571 16819 9577
rect 16761 9537 16773 9571
rect 16807 9568 16819 9571
rect 16850 9568 16856 9580
rect 16807 9540 16856 9568
rect 16807 9537 16819 9540
rect 16761 9531 16819 9537
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 17865 9571 17923 9577
rect 17865 9537 17877 9571
rect 17911 9568 17923 9571
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 17911 9540 18521 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 18509 9537 18521 9540
rect 18555 9568 18567 9571
rect 18782 9568 18788 9580
rect 18555 9540 18788 9568
rect 18555 9537 18567 9540
rect 18509 9531 18567 9537
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 13078 9500 13084 9512
rect 12299 9472 13084 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14424 9472 14841 9500
rect 14424 9460 14430 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 16390 9500 16396 9512
rect 16351 9472 16396 9500
rect 14829 9463 14887 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16540 9503 16598 9509
rect 16540 9469 16552 9503
rect 16586 9500 16598 9503
rect 17494 9500 17500 9512
rect 16586 9472 17500 9500
rect 16586 9469 16598 9472
rect 16540 9463 16598 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 17880 9432 17908 9531
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 21266 9568 21272 9580
rect 21227 9540 21272 9568
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 25777 9571 25835 9577
rect 25777 9568 25789 9571
rect 25307 9540 25789 9568
rect 18288 9503 18346 9509
rect 18288 9469 18300 9503
rect 18334 9500 18346 9503
rect 19242 9500 19248 9512
rect 18334 9472 19248 9500
rect 18334 9469 18346 9472
rect 18288 9463 18346 9469
rect 19242 9460 19248 9472
rect 19300 9500 19306 9512
rect 19889 9503 19947 9509
rect 19889 9500 19901 9503
rect 19300 9472 19901 9500
rect 19300 9460 19306 9472
rect 19889 9469 19901 9472
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 20438 9460 20444 9512
rect 20496 9500 20502 9512
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 20496 9472 20637 9500
rect 20496 9460 20502 9472
rect 20625 9469 20637 9472
rect 20671 9500 20683 9503
rect 20806 9500 20812 9512
rect 20671 9472 20812 9500
rect 20671 9469 20683 9472
rect 20625 9463 20683 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 21177 9503 21235 9509
rect 21177 9469 21189 9503
rect 21223 9500 21235 9503
rect 21358 9500 21364 9512
rect 21223 9472 21364 9500
rect 21223 9469 21235 9472
rect 21177 9463 21235 9469
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 25307 9509 25335 9540
rect 25777 9537 25789 9540
rect 25823 9568 25835 9571
rect 27614 9568 27620 9580
rect 25823 9540 27620 9568
rect 25823 9537 25835 9540
rect 25777 9531 25835 9537
rect 27614 9528 27620 9540
rect 27672 9528 27678 9580
rect 23477 9503 23535 9509
rect 23477 9500 23489 9503
rect 22336 9472 23489 9500
rect 22336 9460 22342 9472
rect 23477 9469 23489 9472
rect 23523 9500 23535 9503
rect 23753 9503 23811 9509
rect 23753 9500 23765 9503
rect 23523 9472 23765 9500
rect 23523 9469 23535 9472
rect 23477 9463 23535 9469
rect 23753 9469 23765 9472
rect 23799 9469 23811 9503
rect 23753 9463 23811 9469
rect 25292 9503 25350 9509
rect 25292 9469 25304 9503
rect 25338 9469 25350 9503
rect 25292 9463 25350 9469
rect 18138 9432 18144 9444
rect 16494 9404 17908 9432
rect 18051 9404 18144 9432
rect 11885 9367 11943 9373
rect 11885 9333 11897 9367
rect 11931 9364 11943 9367
rect 12710 9364 12716 9376
rect 11931 9336 12716 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 15470 9364 15476 9376
rect 15431 9336 15476 9364
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 15930 9364 15936 9376
rect 15843 9336 15936 9364
rect 15930 9324 15936 9336
rect 15988 9364 15994 9376
rect 16494 9364 16522 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 18877 9435 18935 9441
rect 18877 9401 18889 9435
rect 18923 9432 18935 9435
rect 19426 9432 19432 9444
rect 18923 9404 19432 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 17402 9364 17408 9376
rect 15988 9336 16522 9364
rect 17363 9336 17408 9364
rect 15988 9324 15994 9336
rect 17402 9324 17408 9336
rect 17460 9364 17466 9376
rect 18156 9364 18184 9392
rect 19150 9364 19156 9376
rect 17460 9336 18184 9364
rect 19111 9336 19156 9364
rect 17460 9324 17466 9336
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 23934 9364 23940 9376
rect 23895 9336 23940 9364
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 14093 9163 14151 9169
rect 14093 9129 14105 9163
rect 14139 9160 14151 9163
rect 14274 9160 14280 9172
rect 14139 9132 14280 9160
rect 14139 9129 14151 9132
rect 14093 9123 14151 9129
rect 14274 9120 14280 9132
rect 14332 9120 14338 9172
rect 14369 9163 14427 9169
rect 14369 9129 14381 9163
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 16485 9163 16543 9169
rect 16485 9129 16497 9163
rect 16531 9160 16543 9163
rect 16574 9160 16580 9172
rect 16531 9132 16580 9160
rect 16531 9129 16543 9132
rect 16485 9123 16543 9129
rect 12342 9092 12348 9104
rect 12268 9064 12348 9092
rect 12268 9033 12296 9064
rect 12342 9052 12348 9064
rect 12400 9052 12406 9104
rect 14384 9092 14412 9123
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 17221 9163 17279 9169
rect 17221 9129 17233 9163
rect 17267 9160 17279 9163
rect 17494 9160 17500 9172
rect 17267 9132 17500 9160
rect 17267 9129 17279 9132
rect 17221 9123 17279 9129
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18785 9163 18843 9169
rect 18785 9160 18797 9163
rect 18196 9132 18797 9160
rect 18196 9120 18202 9132
rect 18785 9129 18797 9132
rect 18831 9129 18843 9163
rect 18785 9123 18843 9129
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 19981 9163 20039 9169
rect 19981 9160 19993 9163
rect 19576 9132 19993 9160
rect 19576 9120 19582 9132
rect 19981 9129 19993 9132
rect 20027 9129 20039 9163
rect 19981 9123 20039 9129
rect 20254 9120 20260 9172
rect 20312 9160 20318 9172
rect 20717 9163 20775 9169
rect 20717 9160 20729 9163
rect 20312 9132 20729 9160
rect 20312 9120 20318 9132
rect 20717 9129 20729 9132
rect 20763 9160 20775 9163
rect 21177 9163 21235 9169
rect 21177 9160 21189 9163
rect 20763 9132 21189 9160
rect 20763 9129 20775 9132
rect 20717 9123 20775 9129
rect 21177 9129 21189 9132
rect 21223 9160 21235 9163
rect 21358 9160 21364 9172
rect 21223 9132 21364 9160
rect 21223 9129 21235 9132
rect 21177 9123 21235 9129
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 24946 9160 24952 9172
rect 23768 9132 24952 9160
rect 14734 9092 14740 9104
rect 14384 9064 14740 9092
rect 14734 9052 14740 9064
rect 14792 9092 14798 9104
rect 15286 9092 15292 9104
rect 14792 9064 15292 9092
rect 14792 9052 14798 9064
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 22278 9092 22284 9104
rect 22239 9064 22284 9092
rect 22278 9052 22284 9064
rect 22336 9052 22342 9104
rect 23768 9101 23796 9132
rect 24946 9120 24952 9132
rect 25004 9120 25010 9172
rect 23753 9095 23811 9101
rect 23753 9061 23765 9095
rect 23799 9061 23811 9095
rect 23753 9055 23811 9061
rect 23845 9095 23903 9101
rect 23845 9061 23857 9095
rect 23891 9092 23903 9095
rect 23934 9092 23940 9104
rect 23891 9064 23940 9092
rect 23891 9061 23903 9064
rect 23845 9055 23903 9061
rect 23934 9052 23940 9064
rect 23992 9052 23998 9104
rect 24210 9052 24216 9104
rect 24268 9092 24274 9104
rect 25225 9095 25283 9101
rect 25225 9092 25237 9095
rect 24268 9064 25237 9092
rect 24268 9052 24274 9064
rect 25225 9061 25237 9064
rect 25271 9061 25283 9095
rect 25225 9055 25283 9061
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 12342 8956 12348 8968
rect 11296 8928 12348 8956
rect 11296 8916 11302 8928
rect 12342 8916 12348 8928
rect 12400 8956 12406 8968
rect 12544 8956 12572 8987
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13872 8996 14197 9024
rect 13872 8984 13878 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 15436 9027 15494 9033
rect 15436 8993 15448 9027
rect 15482 9024 15494 9027
rect 15562 9024 15568 9036
rect 15482 8996 15568 9024
rect 15482 8993 15494 8996
rect 15436 8987 15494 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 9024 18107 9027
rect 18230 9024 18236 9036
rect 18095 8996 18236 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 8993 18383 9027
rect 18325 8987 18383 8993
rect 15657 8959 15715 8965
rect 12400 8928 13814 8956
rect 12400 8916 12406 8928
rect 13786 8888 13814 8928
rect 15657 8925 15669 8959
rect 15703 8956 15715 8959
rect 15930 8956 15936 8968
rect 15703 8928 15936 8956
rect 15703 8925 15715 8928
rect 15657 8919 15715 8925
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 18340 8956 18368 8987
rect 22186 8956 22192 8968
rect 17828 8928 18368 8956
rect 22147 8928 22192 8956
rect 17828 8916 17834 8928
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 24026 8916 24032 8968
rect 24084 8956 24090 8968
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 24084 8928 24409 8956
rect 24084 8916 24090 8928
rect 24397 8925 24409 8928
rect 24443 8956 24455 8959
rect 24673 8959 24731 8965
rect 24673 8956 24685 8959
rect 24443 8928 24685 8956
rect 24443 8925 24455 8928
rect 24397 8919 24455 8925
rect 24673 8925 24685 8928
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 15749 8891 15807 8897
rect 15749 8888 15761 8891
rect 13786 8860 15761 8888
rect 15749 8857 15761 8860
rect 15795 8857 15807 8891
rect 15749 8851 15807 8857
rect 17494 8848 17500 8900
rect 17552 8888 17558 8900
rect 17865 8891 17923 8897
rect 17865 8888 17877 8891
rect 17552 8860 17877 8888
rect 17552 8848 17558 8860
rect 17865 8857 17877 8860
rect 17911 8857 17923 8891
rect 17865 8851 17923 8857
rect 22741 8891 22799 8897
rect 22741 8857 22753 8891
rect 22787 8888 22799 8891
rect 24044 8888 24072 8916
rect 22787 8860 24072 8888
rect 22787 8857 22799 8860
rect 22741 8851 22799 8857
rect 8662 8820 8668 8832
rect 8623 8792 8668 8820
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12584 8792 13001 8820
rect 12584 8780 12590 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 12989 8783 13047 8789
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15378 8820 15384 8832
rect 14967 8792 15384 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15378 8780 15384 8792
rect 15436 8820 15442 8832
rect 15565 8823 15623 8829
rect 15565 8820 15577 8823
rect 15436 8792 15577 8820
rect 15436 8780 15442 8792
rect 15565 8789 15577 8792
rect 15611 8820 15623 8823
rect 15838 8820 15844 8832
rect 15611 8792 15844 8820
rect 15611 8789 15623 8792
rect 15565 8783 15623 8789
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 16853 8823 16911 8829
rect 16853 8789 16865 8823
rect 16899 8820 16911 8823
rect 18598 8820 18604 8832
rect 16899 8792 18604 8820
rect 16899 8789 16911 8792
rect 16853 8783 16911 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 19242 8820 19248 8832
rect 19203 8792 19248 8820
rect 19242 8780 19248 8792
rect 19300 8780 19306 8832
rect 19334 8780 19340 8832
rect 19392 8820 19398 8832
rect 19702 8820 19708 8832
rect 19392 8792 19708 8820
rect 19392 8780 19398 8792
rect 19702 8780 19708 8792
rect 19760 8780 19766 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 11238 8616 11244 8628
rect 11199 8588 11244 8616
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12250 8616 12256 8628
rect 11931 8588 12256 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12250 8576 12256 8588
rect 12308 8616 12314 8628
rect 13078 8616 13084 8628
rect 12308 8588 13084 8616
rect 12308 8576 12314 8588
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 15654 8576 15660 8628
rect 15712 8616 15718 8628
rect 15749 8619 15807 8625
rect 15749 8616 15761 8619
rect 15712 8588 15761 8616
rect 15712 8576 15718 8588
rect 15749 8585 15761 8588
rect 15795 8585 15807 8619
rect 15749 8579 15807 8585
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 16117 8619 16175 8625
rect 16117 8616 16129 8619
rect 15896 8588 16129 8616
rect 15896 8576 15902 8588
rect 16117 8585 16129 8588
rect 16163 8616 16175 8619
rect 19702 8616 19708 8628
rect 16163 8588 19708 8616
rect 16163 8585 16175 8588
rect 16117 8579 16175 8585
rect 19702 8576 19708 8588
rect 19760 8616 19766 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19760 8588 19901 8616
rect 19760 8576 19766 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 20254 8616 20260 8628
rect 20215 8588 20260 8616
rect 19889 8579 19947 8585
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 22189 8619 22247 8625
rect 22189 8585 22201 8619
rect 22235 8616 22247 8619
rect 22278 8616 22284 8628
rect 22235 8588 22284 8616
rect 22235 8585 22247 8588
rect 22189 8579 22247 8585
rect 22278 8576 22284 8588
rect 22336 8616 22342 8628
rect 22465 8619 22523 8625
rect 22465 8616 22477 8619
rect 22336 8588 22477 8616
rect 22336 8576 22342 8588
rect 22465 8585 22477 8588
rect 22511 8585 22523 8619
rect 22465 8579 22523 8585
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23934 8616 23940 8628
rect 23523 8588 23940 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23934 8576 23940 8588
rect 23992 8576 23998 8628
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25547 8619 25605 8625
rect 25547 8616 25559 8619
rect 25464 8588 25559 8616
rect 25464 8576 25470 8588
rect 25547 8585 25559 8588
rect 25593 8585 25605 8619
rect 25547 8579 25605 8585
rect 14366 8508 14372 8560
rect 14424 8548 14430 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 14424 8520 15393 8548
rect 14424 8508 14430 8520
rect 15381 8517 15393 8520
rect 15427 8548 15439 8551
rect 15930 8548 15936 8560
rect 15427 8520 15936 8548
rect 15427 8517 15439 8520
rect 15381 8511 15439 8517
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 17402 8548 17408 8560
rect 16408 8520 17408 8548
rect 9030 8480 9036 8492
rect 8991 8452 9036 8480
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 12526 8480 12532 8492
rect 11379 8452 12532 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12894 8480 12900 8492
rect 12855 8452 12900 8480
rect 12894 8440 12900 8452
rect 12952 8440 12958 8492
rect 13814 8480 13820 8492
rect 13775 8452 13820 8480
rect 13814 8440 13820 8452
rect 13872 8480 13878 8492
rect 16408 8480 16436 8520
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 19337 8551 19395 8557
rect 19337 8517 19349 8551
rect 19383 8548 19395 8551
rect 22646 8548 22652 8560
rect 19383 8520 22652 8548
rect 19383 8517 19395 8520
rect 19337 8511 19395 8517
rect 22646 8508 22652 8520
rect 22704 8508 22710 8560
rect 13872 8452 16436 8480
rect 16485 8483 16543 8489
rect 13872 8440 13878 8452
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16531 8452 18736 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 14274 8412 14280 8424
rect 14235 8384 14280 8412
rect 9217 8375 9275 8381
rect 9232 8344 9260 8375
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 15470 8412 15476 8424
rect 14599 8384 15476 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 8588 8316 9260 8344
rect 12621 8347 12679 8353
rect 8588 8288 8616 8316
rect 12621 8313 12633 8347
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 13541 8347 13599 8353
rect 13541 8313 13553 8347
rect 13587 8344 13599 8347
rect 13998 8344 14004 8356
rect 13587 8316 14004 8344
rect 13587 8313 13599 8316
rect 13541 8307 13599 8313
rect 8570 8276 8576 8288
rect 8531 8248 8576 8276
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 12158 8276 12164 8288
rect 12119 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8276 12222 8288
rect 12636 8276 12664 8307
rect 13998 8304 14004 8316
rect 14056 8344 14062 8356
rect 14568 8344 14596 8375
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 16114 8412 16120 8424
rect 15611 8384 16120 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 16114 8372 16120 8384
rect 16172 8412 16178 8424
rect 16592 8421 16620 8452
rect 18708 8421 18736 8452
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 19521 8483 19579 8489
rect 19521 8480 19533 8483
rect 18840 8452 19533 8480
rect 18840 8440 18846 8452
rect 19521 8449 19533 8452
rect 19567 8480 19579 8483
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19567 8452 19993 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21450 8480 21456 8492
rect 21315 8452 21456 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22244 8452 22845 8480
rect 22244 8440 22250 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8480 23995 8483
rect 24026 8480 24032 8492
rect 23983 8452 24032 8480
rect 23983 8449 23995 8452
rect 23937 8443 23995 8449
rect 24026 8440 24032 8452
rect 24084 8440 24090 8492
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8480 24639 8483
rect 24670 8480 24676 8492
rect 24627 8452 24676 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 16577 8415 16635 8421
rect 16172 8384 16522 8412
rect 16172 8372 16178 8384
rect 14056 8316 14596 8344
rect 14056 8304 14062 8316
rect 14090 8276 14096 8288
rect 12216 8248 12664 8276
rect 14051 8248 14096 8276
rect 12216 8236 12222 8248
rect 14090 8236 14096 8248
rect 14148 8236 14154 8288
rect 16494 8276 16522 8384
rect 16577 8381 16589 8415
rect 16623 8381 16635 8415
rect 16577 8375 16635 8381
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8412 16819 8415
rect 18693 8415 18751 8421
rect 16807 8384 16988 8412
rect 16807 8381 16819 8384
rect 16761 8375 16819 8381
rect 16850 8276 16856 8288
rect 16494 8248 16856 8276
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 16960 8276 16988 8384
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 18708 8344 18736 8375
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 19760 8415 19818 8421
rect 19760 8412 19772 8415
rect 19300 8384 19772 8412
rect 19300 8372 19306 8384
rect 19760 8381 19772 8384
rect 19806 8412 19818 8415
rect 20625 8415 20683 8421
rect 20625 8412 20637 8415
rect 19806 8384 20637 8412
rect 19806 8381 19818 8384
rect 19760 8375 19818 8381
rect 20625 8381 20637 8384
rect 20671 8381 20683 8415
rect 21174 8412 21180 8424
rect 21087 8384 21180 8412
rect 20625 8375 20683 8381
rect 21174 8372 21180 8384
rect 21232 8412 21238 8424
rect 22002 8412 22008 8424
rect 21232 8384 22008 8412
rect 21232 8372 21238 8384
rect 19153 8347 19211 8353
rect 19153 8344 19165 8347
rect 18708 8316 19165 8344
rect 19153 8313 19165 8316
rect 19199 8344 19211 8347
rect 19337 8347 19395 8353
rect 19337 8344 19349 8347
rect 19199 8316 19349 8344
rect 19199 8313 19211 8316
rect 19153 8307 19211 8313
rect 19337 8313 19349 8316
rect 19383 8313 19395 8347
rect 19337 8307 19395 8313
rect 19518 8304 19524 8356
rect 19576 8344 19582 8356
rect 21646 8353 21674 8384
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 25476 8415 25534 8421
rect 25476 8381 25488 8415
rect 25522 8412 25534 8415
rect 25522 8384 26004 8412
rect 25522 8381 25534 8384
rect 25476 8375 25534 8381
rect 19612 8347 19670 8353
rect 19612 8344 19624 8347
rect 19576 8316 19624 8344
rect 19576 8304 19582 8316
rect 19612 8313 19624 8316
rect 19658 8313 19670 8347
rect 21631 8347 21689 8353
rect 21631 8344 21643 8347
rect 21609 8316 21643 8344
rect 19612 8307 19670 8313
rect 21631 8313 21643 8316
rect 21677 8313 21689 8347
rect 24026 8344 24032 8356
rect 23987 8316 24032 8344
rect 21631 8307 21689 8313
rect 24026 8304 24032 8316
rect 24084 8304 24090 8356
rect 17497 8279 17555 8285
rect 17497 8276 17509 8279
rect 16960 8248 17509 8276
rect 17497 8245 17509 8248
rect 17543 8276 17555 8279
rect 17770 8276 17776 8288
rect 17543 8248 17776 8276
rect 17543 8245 17555 8248
rect 17497 8239 17555 8245
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 18322 8276 18328 8288
rect 18283 8248 18328 8276
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 25976 8285 26004 8384
rect 25961 8279 26019 8285
rect 25961 8245 25973 8279
rect 26007 8276 26019 8279
rect 27614 8276 27620 8288
rect 26007 8248 27620 8276
rect 26007 8245 26019 8248
rect 25961 8239 26019 8245
rect 27614 8236 27620 8248
rect 27672 8236 27678 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 12434 8072 12440 8084
rect 12395 8044 12440 8072
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 14366 8072 14372 8084
rect 14327 8044 14372 8072
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 14734 8072 14740 8084
rect 14695 8044 14740 8072
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15105 8075 15163 8081
rect 15105 8041 15117 8075
rect 15151 8072 15163 8075
rect 15654 8072 15660 8084
rect 15151 8044 15660 8072
rect 15151 8041 15163 8044
rect 15105 8035 15163 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16850 8072 16856 8084
rect 16439 8044 16856 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 17092 8044 18245 8072
rect 17092 8032 17098 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 18233 8035 18291 8041
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 21450 8072 21456 8084
rect 21407 8044 21456 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 23937 8075 23995 8081
rect 23937 8041 23949 8075
rect 23983 8072 23995 8075
rect 24026 8072 24032 8084
rect 23983 8044 24032 8072
rect 23983 8041 23995 8044
rect 23937 8035 23995 8041
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 8754 8004 8760 8016
rect 8715 7976 8760 8004
rect 8754 7964 8760 7976
rect 8812 7964 8818 8016
rect 11241 8007 11299 8013
rect 11241 7973 11253 8007
rect 11287 8004 11299 8007
rect 12158 8004 12164 8016
rect 11287 7976 12164 8004
rect 11287 7973 11299 7976
rect 11241 7967 11299 7973
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 20346 8004 20352 8016
rect 19352 7976 20352 8004
rect 19352 7948 19380 7976
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 22002 7964 22008 8016
rect 22060 8004 22066 8016
rect 22234 8007 22292 8013
rect 22234 8004 22246 8007
rect 22060 7976 22246 8004
rect 22060 7964 22066 7976
rect 22234 7973 22246 7976
rect 22280 7973 22292 8007
rect 24210 8004 24216 8016
rect 24171 7976 24216 8004
rect 22234 7967 22292 7973
rect 24210 7964 24216 7976
rect 24268 7964 24274 8016
rect 24305 8007 24363 8013
rect 24305 7973 24317 8007
rect 24351 8004 24363 8007
rect 24670 8004 24676 8016
rect 24351 7976 24676 8004
rect 24351 7973 24363 7976
rect 24305 7967 24363 7973
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 8202 7936 8208 7948
rect 8163 7908 8208 7936
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8570 7936 8576 7948
rect 8435 7908 8576 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 10594 7936 10600 7948
rect 10555 7908 10600 7936
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 12066 7936 12072 7948
rect 12027 7908 12072 7936
rect 12066 7896 12072 7908
rect 12124 7896 12130 7948
rect 14182 7936 14188 7948
rect 14143 7908 14188 7936
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 15286 7936 15292 7948
rect 15247 7908 15292 7936
rect 15286 7896 15292 7908
rect 15344 7896 15350 7948
rect 15746 7936 15752 7948
rect 15707 7908 15752 7936
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 17000 7908 17601 7936
rect 17000 7896 17006 7908
rect 17589 7905 17601 7908
rect 17635 7936 17647 7939
rect 18322 7936 18328 7948
rect 17635 7908 18328 7936
rect 17635 7905 17647 7908
rect 17589 7899 17647 7905
rect 18322 7896 18328 7908
rect 18380 7936 18386 7948
rect 18601 7939 18659 7945
rect 18601 7936 18613 7939
rect 18380 7908 18613 7936
rect 18380 7896 18386 7908
rect 18601 7905 18613 7908
rect 18647 7905 18659 7939
rect 19334 7936 19340 7948
rect 19247 7908 19340 7936
rect 18601 7899 18659 7905
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 19426 7896 19432 7948
rect 19484 7936 19490 7948
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 19484 7908 19717 7936
rect 19484 7896 19490 7908
rect 19705 7905 19717 7908
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 21266 7896 21272 7948
rect 21324 7936 21330 7948
rect 21913 7939 21971 7945
rect 21913 7936 21925 7939
rect 21324 7908 21925 7936
rect 21324 7896 21330 7908
rect 21913 7905 21925 7908
rect 21959 7936 21971 7939
rect 22370 7936 22376 7948
rect 21959 7908 22376 7936
rect 21959 7905 21971 7908
rect 21913 7899 21971 7905
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14274 7868 14280 7880
rect 14139 7840 14280 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 14108 7800 14136 7831
rect 14274 7828 14280 7840
rect 14332 7868 14338 7880
rect 15304 7868 15332 7896
rect 16022 7868 16028 7880
rect 14332 7840 15332 7868
rect 15983 7840 16028 7868
rect 14332 7828 14338 7840
rect 16022 7828 16028 7840
rect 16080 7828 16086 7880
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17276 7840 17969 7868
rect 17276 7828 17282 7840
rect 17957 7837 17969 7840
rect 18003 7868 18015 7871
rect 19150 7868 19156 7880
rect 18003 7840 19156 7868
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 19150 7828 19156 7840
rect 19208 7828 19214 7880
rect 19978 7868 19984 7880
rect 19939 7840 19984 7868
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 24578 7868 24584 7880
rect 24539 7840 24584 7868
rect 24578 7828 24584 7840
rect 24636 7828 24642 7880
rect 11848 7772 14136 7800
rect 11848 7760 11854 7772
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 12802 7732 12808 7744
rect 10652 7704 12808 7732
rect 10652 7692 10658 7704
rect 12802 7692 12808 7704
rect 12860 7732 12866 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12860 7704 13001 7732
rect 12860 7692 12866 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 17494 7732 17500 7744
rect 17455 7704 17500 7732
rect 12989 7695 13047 7701
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 17770 7741 17776 7744
rect 17754 7735 17776 7741
rect 17754 7701 17766 7735
rect 17754 7695 17776 7701
rect 17770 7692 17776 7695
rect 17828 7692 17834 7744
rect 17862 7692 17868 7744
rect 17920 7732 17926 7744
rect 22833 7735 22891 7741
rect 17920 7704 17965 7732
rect 17920 7692 17926 7704
rect 22833 7701 22845 7735
rect 22879 7732 22891 7735
rect 24026 7732 24032 7744
rect 22879 7704 24032 7732
rect 22879 7701 22891 7704
rect 22833 7695 22891 7701
rect 24026 7692 24032 7704
rect 24084 7692 24090 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 10594 7528 10600 7540
rect 10555 7500 10600 7528
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 12066 7528 12072 7540
rect 11839 7500 12072 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 12161 7531 12219 7537
rect 12161 7497 12173 7531
rect 12207 7528 12219 7531
rect 12434 7528 12440 7540
rect 12207 7500 12440 7528
rect 12207 7497 12219 7500
rect 12161 7491 12219 7497
rect 12434 7488 12440 7500
rect 12492 7528 12498 7540
rect 13630 7528 13636 7540
rect 12492 7500 13636 7528
rect 12492 7488 12498 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 15013 7531 15071 7537
rect 15013 7497 15025 7531
rect 15059 7528 15071 7531
rect 15286 7528 15292 7540
rect 15059 7500 15292 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 19334 7528 19340 7540
rect 19295 7500 19340 7528
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 19613 7531 19671 7537
rect 19613 7528 19625 7531
rect 19484 7500 19625 7528
rect 19484 7488 19490 7500
rect 19613 7497 19625 7500
rect 19659 7528 19671 7531
rect 20441 7531 20499 7537
rect 20441 7528 20453 7531
rect 19659 7500 20453 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 20441 7497 20453 7500
rect 20487 7497 20499 7531
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20441 7491 20499 7497
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 15930 7460 15936 7472
rect 12584 7432 15936 7460
rect 12584 7420 12590 7432
rect 15930 7420 15936 7432
rect 15988 7460 15994 7472
rect 17589 7463 17647 7469
rect 17589 7460 17601 7463
rect 15988 7432 17601 7460
rect 15988 7420 15994 7432
rect 17589 7429 17601 7432
rect 17635 7460 17647 7463
rect 17862 7460 17868 7472
rect 17635 7432 17868 7460
rect 17635 7429 17647 7432
rect 17589 7423 17647 7429
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8202 7392 8208 7404
rect 7975 7364 8208 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8202 7352 8208 7364
rect 8260 7392 8266 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8260 7364 8493 7392
rect 8260 7352 8266 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12952 7364 13001 7392
rect 12952 7352 12958 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 20456 7392 20484 7491
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 22370 7528 22376 7540
rect 22331 7500 22376 7528
rect 22370 7488 22376 7500
rect 22428 7488 22434 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 24210 7528 24216 7540
rect 23523 7500 24216 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 25222 7488 25228 7540
rect 25280 7528 25286 7540
rect 25455 7531 25513 7537
rect 25455 7528 25467 7531
rect 25280 7500 25467 7528
rect 25280 7488 25286 7500
rect 25455 7497 25467 7500
rect 25501 7497 25513 7531
rect 25455 7491 25513 7497
rect 24489 7395 24547 7401
rect 20456 7364 21496 7392
rect 12989 7355 13047 7361
rect 1210 7284 1216 7336
rect 1268 7324 1274 7336
rect 1432 7327 1490 7333
rect 1432 7324 1444 7327
rect 1268 7296 1444 7324
rect 1268 7284 1274 7296
rect 1432 7293 1444 7296
rect 1478 7324 1490 7327
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1478 7296 1869 7324
rect 1478 7293 1490 7296
rect 1432 7287 1490 7293
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 8662 7324 8668 7336
rect 8623 7296 8668 7324
rect 1857 7287 1915 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 15473 7327 15531 7333
rect 15473 7293 15485 7327
rect 15519 7293 15531 7327
rect 15473 7287 15531 7293
rect 1535 7259 1593 7265
rect 1535 7225 1547 7259
rect 1581 7256 1593 7259
rect 7742 7256 7748 7268
rect 1581 7228 7748 7256
rect 1581 7225 1593 7228
rect 1535 7219 1593 7225
rect 7742 7216 7748 7228
rect 7800 7216 7806 7268
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7225 12771 7259
rect 12713 7219 12771 7225
rect 8297 7191 8355 7197
rect 8297 7157 8309 7191
rect 8343 7188 8355 7191
rect 8570 7188 8576 7200
rect 8343 7160 8576 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 12728 7188 12756 7219
rect 12802 7216 12808 7268
rect 12860 7256 12866 7268
rect 12860 7228 12905 7256
rect 12860 7216 12866 7228
rect 13078 7216 13084 7268
rect 13136 7256 13142 7268
rect 13722 7256 13728 7268
rect 13136 7228 13728 7256
rect 13136 7216 13142 7228
rect 13722 7216 13728 7228
rect 13780 7256 13786 7268
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 13780 7228 15301 7256
rect 13780 7216 13786 7228
rect 15289 7225 15301 7228
rect 15335 7256 15347 7259
rect 15488 7256 15516 7287
rect 15746 7284 15752 7336
rect 15804 7324 15810 7336
rect 15933 7327 15991 7333
rect 15933 7324 15945 7327
rect 15804 7296 15945 7324
rect 15804 7284 15810 7296
rect 15933 7293 15945 7296
rect 15979 7293 15991 7327
rect 15933 7287 15991 7293
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 17954 7324 17960 7336
rect 17552 7296 17960 7324
rect 17552 7284 17558 7296
rect 17954 7284 17960 7296
rect 18012 7324 18018 7336
rect 18141 7327 18199 7333
rect 18141 7324 18153 7327
rect 18012 7296 18153 7324
rect 18012 7284 18018 7296
rect 18141 7293 18153 7296
rect 18187 7324 18199 7327
rect 18782 7324 18788 7336
rect 18187 7296 18788 7324
rect 18187 7293 18199 7296
rect 18141 7287 18199 7293
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21468 7333 21496 7364
rect 24489 7361 24501 7395
rect 24535 7392 24547 7395
rect 24670 7392 24676 7404
rect 24535 7364 24676 7392
rect 24535 7361 24547 7364
rect 24489 7355 24547 7361
rect 24670 7352 24676 7364
rect 24728 7392 24734 7404
rect 24765 7395 24823 7401
rect 24765 7392 24777 7395
rect 24728 7364 24777 7392
rect 24728 7352 24734 7364
rect 24765 7361 24777 7364
rect 24811 7361 24823 7395
rect 24765 7355 24823 7361
rect 20993 7327 21051 7333
rect 20993 7324 21005 7327
rect 20864 7296 21005 7324
rect 20864 7284 20870 7296
rect 20993 7293 21005 7296
rect 21039 7293 21051 7327
rect 20993 7287 21051 7293
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7293 21511 7327
rect 24026 7324 24032 7336
rect 23987 7296 24032 7324
rect 21453 7287 21511 7293
rect 24026 7284 24032 7296
rect 24084 7284 24090 7336
rect 25384 7327 25442 7333
rect 25384 7293 25396 7327
rect 25430 7324 25442 7327
rect 25869 7327 25927 7333
rect 25869 7324 25881 7327
rect 25430 7296 25881 7324
rect 25430 7293 25442 7296
rect 25384 7287 25442 7293
rect 25869 7293 25881 7296
rect 25915 7324 25927 7327
rect 27614 7324 27620 7336
rect 25915 7296 27620 7324
rect 25915 7293 25927 7296
rect 25869 7287 25927 7293
rect 27614 7284 27620 7296
rect 27672 7284 27678 7336
rect 16206 7256 16212 7268
rect 15335 7228 15516 7256
rect 16167 7228 16212 7256
rect 15335 7225 15347 7228
rect 15289 7219 15347 7225
rect 16206 7216 16212 7228
rect 16264 7216 16270 7268
rect 21726 7256 21732 7268
rect 21687 7228 21732 7256
rect 21726 7216 21732 7228
rect 21784 7216 21790 7268
rect 13262 7188 13268 7200
rect 12728 7160 13268 7188
rect 13262 7148 13268 7160
rect 13320 7188 13326 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13320 7160 13645 7188
rect 13320 7148 13326 7160
rect 13633 7157 13645 7160
rect 13679 7157 13691 7191
rect 13633 7151 13691 7157
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 14240 7160 14289 7188
rect 14240 7148 14246 7160
rect 14277 7157 14289 7160
rect 14323 7188 14335 7191
rect 15470 7188 15476 7200
rect 14323 7160 15476 7188
rect 14323 7157 14335 7160
rect 14277 7151 14335 7157
rect 15470 7148 15476 7160
rect 15528 7188 15534 7200
rect 17218 7188 17224 7200
rect 15528 7160 17224 7188
rect 15528 7148 15534 7160
rect 17218 7148 17224 7160
rect 17276 7148 17282 7200
rect 18322 7188 18328 7200
rect 18283 7160 18328 7188
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 22002 7188 22008 7200
rect 21963 7160 22008 7188
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 12158 6984 12164 6996
rect 12119 6956 12164 6984
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12860 6956 12909 6984
rect 12860 6944 12866 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 15565 6987 15623 6993
rect 15565 6953 15577 6987
rect 15611 6984 15623 6987
rect 15746 6984 15752 6996
rect 15611 6956 15752 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 15746 6944 15752 6956
rect 15804 6984 15810 6996
rect 15841 6987 15899 6993
rect 15841 6984 15853 6987
rect 15804 6956 15853 6984
rect 15804 6944 15810 6956
rect 15841 6953 15853 6956
rect 15887 6953 15899 6987
rect 18782 6984 18788 6996
rect 18743 6956 18788 6984
rect 15841 6947 15899 6953
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 23845 6987 23903 6993
rect 23845 6953 23857 6987
rect 23891 6984 23903 6987
rect 24026 6984 24032 6996
rect 23891 6956 24032 6984
rect 23891 6953 23903 6956
rect 23845 6947 23903 6953
rect 24026 6944 24032 6956
rect 24084 6944 24090 6996
rect 15930 6876 15936 6928
rect 15988 6916 15994 6928
rect 16438 6919 16496 6925
rect 16438 6916 16450 6919
rect 15988 6888 16450 6916
rect 15988 6876 15994 6888
rect 16438 6885 16450 6888
rect 16484 6916 16496 6919
rect 18186 6919 18244 6925
rect 18186 6916 18198 6919
rect 16484 6888 18198 6916
rect 16484 6885 16496 6888
rect 16438 6879 16496 6885
rect 18186 6885 18198 6888
rect 18232 6916 18244 6919
rect 22002 6916 22008 6928
rect 18232 6888 22008 6916
rect 18232 6885 18244 6888
rect 18186 6879 18244 6885
rect 22002 6876 22008 6888
rect 22060 6916 22066 6928
rect 22694 6919 22752 6925
rect 22694 6916 22706 6919
rect 22060 6888 22706 6916
rect 22060 6876 22066 6888
rect 22694 6885 22706 6888
rect 22740 6885 22752 6919
rect 22694 6879 22752 6885
rect 11790 6808 11796 6860
rect 11848 6848 11854 6860
rect 11885 6851 11943 6857
rect 11885 6848 11897 6851
rect 11848 6820 11897 6848
rect 11848 6808 11854 6820
rect 11885 6817 11897 6820
rect 11931 6817 11943 6851
rect 12342 6848 12348 6860
rect 12303 6820 12348 6848
rect 11885 6811 11943 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 13722 6848 13728 6860
rect 13683 6820 13728 6848
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 14056 6820 14105 6848
rect 14056 6808 14062 6820
rect 14093 6817 14105 6820
rect 14139 6817 14151 6851
rect 14093 6811 14151 6817
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16117 6851 16175 6857
rect 16117 6848 16129 6851
rect 16080 6820 16129 6848
rect 16080 6808 16086 6820
rect 16117 6817 16129 6820
rect 16163 6817 16175 6851
rect 16117 6811 16175 6817
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 16264 6820 17877 6848
rect 16264 6808 16270 6820
rect 17865 6817 17877 6820
rect 17911 6848 17923 6851
rect 19426 6848 19432 6860
rect 17911 6820 19432 6848
rect 17911 6817 17923 6820
rect 17865 6811 17923 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 21726 6808 21732 6860
rect 21784 6848 21790 6860
rect 22373 6851 22431 6857
rect 22373 6848 22385 6851
rect 21784 6820 22385 6848
rect 21784 6808 21790 6820
rect 22373 6817 22385 6820
rect 22419 6848 22431 6851
rect 23014 6848 23020 6860
rect 22419 6820 23020 6848
rect 22419 6817 22431 6820
rect 22373 6811 22431 6817
rect 23014 6808 23020 6820
rect 23072 6808 23078 6860
rect 23293 6851 23351 6857
rect 23293 6817 23305 6851
rect 23339 6848 23351 6851
rect 24210 6848 24216 6860
rect 23339 6820 24216 6848
rect 23339 6817 23351 6820
rect 23293 6811 23351 6817
rect 24210 6808 24216 6820
rect 24268 6808 24274 6860
rect 14182 6780 14188 6792
rect 14143 6752 14188 6780
rect 14182 6740 14188 6752
rect 14240 6740 14246 6792
rect 24118 6780 24124 6792
rect 24079 6752 24124 6780
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 2188 6616 8493 6644
rect 2188 6604 2194 6616
rect 8481 6613 8493 6616
rect 8527 6644 8539 6647
rect 8662 6644 8668 6656
rect 8527 6616 8668 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16632 6616 17049 6644
rect 16632 6604 16638 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 17681 6647 17739 6653
rect 17681 6613 17693 6647
rect 17727 6644 17739 6647
rect 17770 6644 17776 6656
rect 17727 6616 17776 6644
rect 17727 6613 17739 6616
rect 17681 6607 17739 6613
rect 17770 6604 17776 6616
rect 17828 6644 17834 6656
rect 19058 6644 19064 6656
rect 17828 6616 19064 6644
rect 17828 6604 17834 6616
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12342 6440 12348 6452
rect 12023 6412 12348 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13998 6440 14004 6452
rect 13219 6412 14004 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 15841 6443 15899 6449
rect 15841 6409 15853 6443
rect 15887 6440 15899 6443
rect 16022 6440 16028 6452
rect 15887 6412 16028 6440
rect 15887 6409 15899 6412
rect 15841 6403 15899 6409
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 19426 6440 19432 6452
rect 19387 6412 19432 6440
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 22002 6400 22008 6452
rect 22060 6440 22066 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 22060 6412 22385 6440
rect 22060 6400 22066 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 22554 6400 22560 6452
rect 22612 6440 22618 6452
rect 22695 6443 22753 6449
rect 22695 6440 22707 6443
rect 22612 6412 22707 6440
rect 22612 6400 22618 6412
rect 22695 6409 22707 6412
rect 22741 6409 22753 6443
rect 23014 6440 23020 6452
rect 22975 6412 23020 6440
rect 22695 6403 22753 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 24029 6443 24087 6449
rect 24029 6409 24041 6443
rect 24075 6440 24087 6443
rect 24118 6440 24124 6452
rect 24075 6412 24124 6440
rect 24075 6409 24087 6412
rect 24029 6403 24087 6409
rect 24118 6400 24124 6412
rect 24176 6400 24182 6452
rect 11790 6332 11796 6384
rect 11848 6372 11854 6384
rect 12621 6375 12679 6381
rect 12621 6372 12633 6375
rect 11848 6344 12633 6372
rect 11848 6332 11854 6344
rect 12621 6341 12633 6344
rect 12667 6341 12679 6375
rect 12621 6335 12679 6341
rect 13541 6375 13599 6381
rect 13541 6341 13553 6375
rect 13587 6372 13599 6375
rect 13722 6372 13728 6384
rect 13587 6344 13728 6372
rect 13587 6341 13599 6344
rect 13541 6335 13599 6341
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 16298 6332 16304 6384
rect 16356 6372 16362 6384
rect 18506 6372 18512 6384
rect 16356 6344 18512 6372
rect 16356 6332 16362 6344
rect 18506 6332 18512 6344
rect 18564 6372 18570 6384
rect 18693 6375 18751 6381
rect 18693 6372 18705 6375
rect 18564 6344 18705 6372
rect 18564 6332 18570 6344
rect 18693 6341 18705 6344
rect 18739 6341 18751 6375
rect 18693 6335 18751 6341
rect 24210 6332 24216 6384
rect 24268 6372 24274 6384
rect 25133 6375 25191 6381
rect 25133 6372 25145 6375
rect 24268 6344 25145 6372
rect 24268 6332 24274 6344
rect 25133 6341 25145 6344
rect 25179 6341 25191 6375
rect 25133 6335 25191 6341
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6304 14059 6307
rect 14182 6304 14188 6316
rect 14047 6276 14188 6304
rect 14047 6273 14059 6276
rect 14001 6267 14059 6273
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 16482 6304 16488 6316
rect 16443 6276 16488 6304
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6304 18199 6307
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 18187 6276 19073 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 19061 6273 19073 6276
rect 19107 6304 19119 6307
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19107 6276 19625 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 24489 6307 24547 6313
rect 24489 6304 24501 6307
rect 19613 6267 19671 6273
rect 23446 6276 24501 6304
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 22592 6239 22650 6245
rect 22592 6236 22604 6239
rect 22143 6208 22604 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 22592 6205 22604 6208
rect 22638 6236 22650 6239
rect 23446 6236 23474 6276
rect 24489 6273 24501 6276
rect 24535 6304 24547 6307
rect 24578 6304 24584 6316
rect 24535 6276 24584 6304
rect 24535 6273 24547 6276
rect 24489 6267 24547 6273
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 22638 6208 23474 6236
rect 22638 6205 22650 6208
rect 22592 6199 22650 6205
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 13817 6171 13875 6177
rect 13817 6168 13829 6171
rect 13688 6140 13829 6168
rect 13688 6128 13694 6140
rect 13817 6137 13829 6140
rect 13863 6168 13875 6171
rect 14322 6171 14380 6177
rect 14322 6168 14334 6171
rect 13863 6140 14334 6168
rect 13863 6137 13875 6140
rect 13817 6131 13875 6137
rect 14322 6137 14334 6140
rect 14368 6168 14380 6171
rect 15930 6168 15936 6180
rect 14368 6140 15936 6168
rect 14368 6137 14380 6140
rect 14322 6131 14380 6137
rect 15930 6128 15936 6140
rect 15988 6168 15994 6180
rect 16117 6171 16175 6177
rect 16117 6168 16129 6171
rect 15988 6140 16129 6168
rect 15988 6128 15994 6140
rect 16117 6137 16129 6140
rect 16163 6137 16175 6171
rect 16117 6131 16175 6137
rect 14921 6103 14979 6109
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15378 6100 15384 6112
rect 14967 6072 15384 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 16132 6100 16160 6131
rect 16574 6128 16580 6180
rect 16632 6168 16638 6180
rect 17126 6168 17132 6180
rect 16632 6140 16677 6168
rect 17087 6140 17132 6168
rect 16632 6128 16638 6140
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 17497 6171 17555 6177
rect 17497 6137 17509 6171
rect 17543 6168 17555 6171
rect 18233 6171 18291 6177
rect 18233 6168 18245 6171
rect 17543 6140 18245 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 18233 6137 18245 6140
rect 18279 6168 18291 6171
rect 18322 6168 18328 6180
rect 18279 6140 18328 6168
rect 18279 6137 18291 6140
rect 18233 6131 18291 6137
rect 18322 6128 18328 6140
rect 18380 6128 18386 6180
rect 21545 6171 21603 6177
rect 21545 6137 21557 6171
rect 21591 6168 21603 6171
rect 23385 6171 23443 6177
rect 23385 6168 23397 6171
rect 21591 6140 23397 6168
rect 21591 6137 21603 6140
rect 21545 6131 21603 6137
rect 23385 6137 23397 6140
rect 23431 6168 23443 6171
rect 24213 6171 24271 6177
rect 24213 6168 24225 6171
rect 23431 6140 24225 6168
rect 23431 6137 23443 6140
rect 23385 6131 23443 6137
rect 24213 6137 24225 6140
rect 24259 6137 24271 6171
rect 24213 6131 24271 6137
rect 24305 6171 24363 6177
rect 24305 6137 24317 6171
rect 24351 6137 24363 6171
rect 24305 6131 24363 6137
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 16132 6072 17785 6100
rect 17773 6069 17785 6072
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 24118 6060 24124 6112
rect 24176 6100 24182 6112
rect 24320 6100 24348 6131
rect 24176 6072 24348 6100
rect 24176 6060 24182 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 14182 5856 14188 5908
rect 14240 5896 14246 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 14240 5868 14657 5896
rect 14240 5856 14246 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16761 5899 16819 5905
rect 16761 5896 16773 5899
rect 16540 5868 16773 5896
rect 16540 5856 16546 5868
rect 16761 5865 16773 5868
rect 16807 5865 16819 5899
rect 16761 5859 16819 5865
rect 24210 5856 24216 5908
rect 24268 5896 24274 5908
rect 24268 5868 24440 5896
rect 24268 5856 24274 5868
rect 13817 5831 13875 5837
rect 13817 5797 13829 5831
rect 13863 5828 13875 5831
rect 13863 5800 15332 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5760 14427 5763
rect 14458 5760 14464 5772
rect 14415 5732 14464 5760
rect 14415 5729 14427 5732
rect 14369 5723 14427 5729
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 15304 5704 15332 5800
rect 17126 5788 17132 5840
rect 17184 5828 17190 5840
rect 17862 5828 17868 5840
rect 17184 5800 17868 5828
rect 17184 5788 17190 5800
rect 17862 5788 17868 5800
rect 17920 5788 17926 5840
rect 17954 5788 17960 5840
rect 18012 5828 18018 5840
rect 18506 5828 18512 5840
rect 18012 5800 18057 5828
rect 18467 5800 18512 5828
rect 18012 5788 18018 5800
rect 18506 5788 18512 5800
rect 18564 5788 18570 5840
rect 22002 5788 22008 5840
rect 22060 5828 22066 5840
rect 24412 5837 24440 5868
rect 22694 5831 22752 5837
rect 22694 5828 22706 5831
rect 22060 5800 22706 5828
rect 22060 5788 22066 5800
rect 22694 5797 22706 5800
rect 22740 5797 22752 5831
rect 22694 5791 22752 5797
rect 24397 5831 24455 5837
rect 24397 5797 24409 5831
rect 24443 5797 24455 5831
rect 24397 5791 24455 5797
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 15436 5732 15481 5760
rect 15436 5720 15442 5732
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 22373 5763 22431 5769
rect 22373 5760 22385 5763
rect 20036 5732 22385 5760
rect 20036 5720 20042 5732
rect 22373 5729 22385 5732
rect 22419 5760 22431 5763
rect 22554 5760 22560 5772
rect 22419 5732 22560 5760
rect 22419 5729 22431 5732
rect 22373 5723 22431 5729
rect 22554 5720 22560 5732
rect 22612 5720 22618 5772
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 13722 5692 13728 5704
rect 12667 5664 13728 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 23474 5652 23480 5704
rect 23532 5692 23538 5704
rect 24305 5695 24363 5701
rect 24305 5692 24317 5695
rect 23532 5664 24317 5692
rect 23532 5652 23538 5664
rect 24305 5661 24317 5664
rect 24351 5661 24363 5695
rect 24578 5692 24584 5704
rect 24539 5664 24584 5692
rect 24305 5655 24363 5661
rect 16485 5627 16543 5633
rect 16485 5593 16497 5627
rect 16531 5624 16543 5627
rect 16574 5624 16580 5636
rect 16531 5596 16580 5624
rect 16531 5593 16543 5596
rect 16485 5587 16543 5593
rect 16574 5584 16580 5596
rect 16632 5624 16638 5636
rect 17402 5624 17408 5636
rect 16632 5596 17408 5624
rect 16632 5584 16638 5596
rect 17402 5584 17408 5596
rect 17460 5584 17466 5636
rect 24320 5624 24348 5655
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 24670 5624 24676 5636
rect 24320 5596 24676 5624
rect 24670 5584 24676 5596
rect 24728 5584 24734 5636
rect 23293 5559 23351 5565
rect 23293 5525 23305 5559
rect 23339 5556 23351 5559
rect 24026 5556 24032 5568
rect 23339 5528 24032 5556
rect 23339 5525 23351 5528
rect 23293 5519 23351 5525
rect 24026 5516 24032 5528
rect 24084 5516 24090 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12943 5355 13001 5361
rect 12943 5352 12955 5355
rect 12768 5324 12955 5352
rect 12768 5312 12774 5324
rect 12943 5321 12955 5324
rect 12989 5321 13001 5355
rect 12943 5315 13001 5321
rect 15105 5355 15163 5361
rect 15105 5321 15117 5355
rect 15151 5352 15163 5355
rect 15286 5352 15292 5364
rect 15151 5324 15292 5352
rect 15151 5321 15163 5324
rect 15105 5315 15163 5321
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17954 5352 17960 5364
rect 17543 5324 17960 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 22002 5312 22008 5364
rect 22060 5352 22066 5364
rect 22373 5355 22431 5361
rect 22373 5352 22385 5355
rect 22060 5324 22385 5352
rect 22060 5312 22066 5324
rect 22373 5321 22385 5324
rect 22419 5321 22431 5355
rect 22373 5315 22431 5321
rect 13722 5244 13728 5296
rect 13780 5284 13786 5296
rect 15381 5287 15439 5293
rect 15381 5284 15393 5287
rect 13780 5256 15393 5284
rect 13780 5244 13786 5256
rect 15381 5253 15393 5256
rect 15427 5253 15439 5287
rect 15381 5247 15439 5253
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5216 13875 5219
rect 14090 5216 14096 5228
rect 13863 5188 14096 5216
rect 13863 5185 13875 5188
rect 13817 5179 13875 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 14516 5188 15945 5216
rect 14516 5176 14522 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 17920 5188 18429 5216
rect 17920 5176 17926 5188
rect 18417 5185 18429 5188
rect 18463 5216 18475 5219
rect 19061 5219 19119 5225
rect 19061 5216 19073 5219
rect 18463 5188 19073 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 19061 5185 19073 5188
rect 19107 5185 19119 5219
rect 19061 5179 19119 5185
rect 12872 5151 12930 5157
rect 12872 5117 12884 5151
rect 12918 5148 12930 5151
rect 13354 5148 13360 5160
rect 12918 5120 13360 5148
rect 12918 5117 12930 5120
rect 12872 5111 12930 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 13964 5120 14749 5148
rect 13964 5108 13970 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 13630 5080 13636 5092
rect 13543 5052 13636 5080
rect 13630 5040 13636 5052
rect 13688 5080 13694 5092
rect 13688 5052 13814 5080
rect 13688 5040 13694 5052
rect 13786 5012 13814 5052
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 15654 5080 15660 5092
rect 14424 5052 15660 5080
rect 14424 5040 14430 5052
rect 15654 5040 15660 5052
rect 15712 5040 15718 5092
rect 15749 5083 15807 5089
rect 15749 5049 15761 5083
rect 15795 5049 15807 5083
rect 18138 5080 18144 5092
rect 18099 5052 18144 5080
rect 15749 5043 15807 5049
rect 14185 5015 14243 5021
rect 14185 5012 14197 5015
rect 13786 4984 14197 5012
rect 14185 4981 14197 4984
rect 14231 4981 14243 5015
rect 14185 4975 14243 4981
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15764 5012 15792 5043
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 18233 5083 18291 5089
rect 18233 5049 18245 5083
rect 18279 5049 18291 5083
rect 22388 5080 22416 5315
rect 22554 5312 22560 5364
rect 22612 5352 22618 5364
rect 22741 5355 22799 5361
rect 22741 5352 22753 5355
rect 22612 5324 22753 5352
rect 22612 5312 22618 5324
rect 22741 5321 22753 5324
rect 22787 5321 22799 5355
rect 22741 5315 22799 5321
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 23532 5324 23577 5352
rect 23532 5312 23538 5324
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 24949 5355 25007 5361
rect 24949 5352 24961 5355
rect 24268 5324 24961 5352
rect 24268 5312 24274 5324
rect 24949 5321 24961 5324
rect 24995 5321 25007 5355
rect 26050 5352 26056 5364
rect 26011 5324 26056 5352
rect 24949 5315 25007 5321
rect 26050 5312 26056 5324
rect 26108 5312 26114 5364
rect 24026 5148 24032 5160
rect 23987 5120 24032 5148
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 25568 5151 25626 5157
rect 25568 5117 25580 5151
rect 25614 5148 25626 5151
rect 26050 5148 26056 5160
rect 25614 5120 26056 5148
rect 25614 5117 25626 5120
rect 25568 5111 25626 5117
rect 26050 5108 26056 5120
rect 26108 5108 26114 5160
rect 25958 5080 25964 5092
rect 22388 5052 25964 5080
rect 18233 5043 18291 5049
rect 16577 5015 16635 5021
rect 16577 5012 16589 5015
rect 15436 4984 16589 5012
rect 15436 4972 15442 4984
rect 16577 4981 16589 4984
rect 16623 5012 16635 5015
rect 16945 5015 17003 5021
rect 16945 5012 16957 5015
rect 16623 4984 16957 5012
rect 16623 4981 16635 4984
rect 16577 4975 16635 4981
rect 16945 4981 16957 4984
rect 16991 4981 17003 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 16945 4975 17003 4981
rect 17770 4972 17776 4984
rect 17828 5012 17834 5024
rect 18248 5012 18276 5043
rect 25958 5040 25964 5052
rect 26016 5040 26022 5092
rect 24394 5012 24400 5024
rect 17828 4984 18276 5012
rect 24355 4984 24400 5012
rect 17828 4972 17834 4984
rect 24394 4972 24400 4984
rect 24452 4972 24458 5024
rect 25038 4972 25044 5024
rect 25096 5012 25102 5024
rect 25639 5015 25697 5021
rect 25639 5012 25651 5015
rect 25096 4984 25651 5012
rect 25096 4972 25102 4984
rect 25639 4981 25651 4984
rect 25685 4981 25697 5015
rect 25639 4975 25697 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14645 4811 14703 4817
rect 14645 4808 14657 4811
rect 14148 4780 14657 4808
rect 14148 4768 14154 4780
rect 14645 4777 14657 4780
rect 14691 4777 14703 4811
rect 14645 4771 14703 4777
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 16301 4811 16359 4817
rect 16301 4808 16313 4811
rect 15712 4780 16313 4808
rect 15712 4768 15718 4780
rect 16301 4777 16313 4780
rect 16347 4777 16359 4811
rect 17770 4808 17776 4820
rect 17731 4780 17776 4808
rect 16301 4771 16359 4777
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 18138 4768 18144 4820
rect 18196 4808 18202 4820
rect 18325 4811 18383 4817
rect 18325 4808 18337 4811
rect 18196 4780 18337 4808
rect 18196 4768 18202 4780
rect 18325 4777 18337 4780
rect 18371 4808 18383 4811
rect 19015 4811 19073 4817
rect 19015 4808 19027 4811
rect 18371 4780 19027 4808
rect 18371 4777 18383 4780
rect 18325 4771 18383 4777
rect 19015 4777 19027 4780
rect 19061 4777 19073 4811
rect 24026 4808 24032 4820
rect 23987 4780 24032 4808
rect 19015 4771 19073 4777
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 13814 4700 13820 4752
rect 13872 4740 13878 4752
rect 13872 4712 15424 4740
rect 13872 4700 13878 4712
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1578 4672 1584 4684
rect 1510 4644 1584 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 15396 4681 15424 4712
rect 24118 4700 24124 4752
rect 24176 4740 24182 4752
rect 24394 4740 24400 4752
rect 24176 4712 24400 4740
rect 24176 4700 24182 4712
rect 24394 4700 24400 4712
rect 24452 4740 24458 4752
rect 24489 4743 24547 4749
rect 24489 4740 24501 4743
rect 24452 4712 24501 4740
rect 24452 4700 24458 4712
rect 24489 4709 24501 4712
rect 24535 4709 24547 4743
rect 24489 4703 24547 4709
rect 24670 4700 24676 4752
rect 24728 4740 24734 4752
rect 25041 4743 25099 4749
rect 25041 4740 25053 4743
rect 24728 4712 25053 4740
rect 24728 4700 24734 4712
rect 25041 4709 25053 4712
rect 25087 4709 25099 4743
rect 25041 4703 25099 4709
rect 15381 4675 15439 4681
rect 15381 4641 15393 4675
rect 15427 4672 15439 4675
rect 15838 4672 15844 4684
rect 15427 4644 15844 4672
rect 15427 4641 15439 4644
rect 15381 4635 15439 4641
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 17402 4672 17408 4684
rect 17363 4644 17408 4672
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 18966 4672 18972 4684
rect 18923 4644 18972 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 15286 4604 15292 4616
rect 15247 4576 15292 4604
rect 15286 4564 15292 4576
rect 15344 4564 15350 4616
rect 24397 4607 24455 4613
rect 24397 4573 24409 4607
rect 24443 4604 24455 4607
rect 25222 4604 25228 4616
rect 24443 4576 25228 4604
rect 24443 4573 24455 4576
rect 24397 4567 24455 4573
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 1535 4539 1593 4545
rect 1535 4505 1547 4539
rect 1581 4536 1593 4539
rect 10502 4536 10508 4548
rect 1581 4508 10508 4536
rect 1581 4505 1593 4508
rect 1535 4499 1593 4505
rect 10502 4496 10508 4508
rect 10560 4496 10566 4548
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 13722 4264 13728 4276
rect 10560 4236 13728 4264
rect 10560 4224 10566 4236
rect 13722 4224 13728 4236
rect 13780 4264 13786 4276
rect 14001 4267 14059 4273
rect 14001 4264 14013 4267
rect 13780 4236 14013 4264
rect 13780 4224 13786 4236
rect 14001 4233 14013 4236
rect 14047 4233 14059 4267
rect 15838 4264 15844 4276
rect 15799 4236 15844 4264
rect 14001 4227 14059 4233
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 18966 4264 18972 4276
rect 18927 4236 18972 4264
rect 18966 4224 18972 4236
rect 19024 4224 19030 4276
rect 24118 4264 24124 4276
rect 24079 4236 24124 4264
rect 24118 4224 24124 4236
rect 24176 4224 24182 4276
rect 25222 4264 25228 4276
rect 25183 4236 25228 4264
rect 25222 4224 25228 4236
rect 25280 4224 25286 4276
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 13814 4128 13820 4140
rect 13771 4100 13820 4128
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15197 4131 15255 4137
rect 15197 4128 15209 4131
rect 14424 4100 15209 4128
rect 14424 4088 14430 4100
rect 15197 4097 15209 4100
rect 15243 4097 15255 4131
rect 24670 4128 24676 4140
rect 24631 4100 24676 4128
rect 15197 4091 15255 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4060 12311 4063
rect 12529 4063 12587 4069
rect 12529 4060 12541 4063
rect 12299 4032 12541 4060
rect 12299 4029 12311 4032
rect 12253 4023 12311 4029
rect 12529 4029 12541 4032
rect 12575 4060 12587 4063
rect 12986 4060 12992 4072
rect 12575 4032 12992 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 14918 3992 14924 4004
rect 14879 3964 14924 3992
rect 14918 3952 14924 3964
rect 14976 3952 14982 4004
rect 15013 3995 15071 4001
rect 15013 3961 15025 3995
rect 15059 3992 15071 3995
rect 15286 3992 15292 4004
rect 15059 3964 15292 3992
rect 15059 3961 15071 3964
rect 15013 3955 15071 3961
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 14737 3927 14795 3933
rect 14737 3893 14749 3927
rect 14783 3924 14795 3927
rect 15028 3924 15056 3955
rect 15286 3952 15292 3964
rect 15344 3952 15350 4004
rect 23477 3995 23535 4001
rect 23477 3961 23489 3995
rect 23523 3992 23535 3995
rect 24302 3992 24308 4004
rect 23523 3964 24308 3992
rect 23523 3961 23535 3964
rect 23477 3955 23535 3961
rect 24302 3952 24308 3964
rect 24360 3952 24366 4004
rect 24397 3995 24455 4001
rect 24397 3961 24409 3995
rect 24443 3961 24455 3995
rect 24397 3955 24455 3961
rect 14783 3896 15056 3924
rect 14783 3893 14795 3896
rect 14737 3887 14795 3893
rect 24026 3884 24032 3936
rect 24084 3924 24090 3936
rect 24412 3924 24440 3955
rect 24084 3896 24440 3924
rect 24084 3884 24090 3896
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 12986 3720 12992 3732
rect 12947 3692 12992 3720
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 14918 3720 14924 3732
rect 14879 3692 14924 3720
rect 14918 3680 14924 3692
rect 14976 3720 14982 3732
rect 15427 3723 15485 3729
rect 15427 3720 15439 3723
rect 14976 3692 15439 3720
rect 14976 3680 14982 3692
rect 15427 3689 15439 3692
rect 15473 3689 15485 3723
rect 15427 3683 15485 3689
rect 24026 3680 24032 3732
rect 24084 3720 24090 3732
rect 24213 3723 24271 3729
rect 24213 3720 24225 3723
rect 24084 3692 24225 3720
rect 24084 3680 24090 3692
rect 24213 3689 24225 3692
rect 24259 3689 24271 3723
rect 24213 3683 24271 3689
rect 24302 3680 24308 3732
rect 24360 3720 24366 3732
rect 24719 3723 24777 3729
rect 24719 3720 24731 3723
rect 24360 3692 24731 3720
rect 24360 3680 24366 3692
rect 24719 3689 24731 3692
rect 24765 3689 24777 3723
rect 24719 3683 24777 3689
rect 12250 3612 12256 3664
rect 12308 3652 12314 3664
rect 12431 3655 12489 3661
rect 12431 3652 12443 3655
rect 12308 3624 12443 3652
rect 12308 3612 12314 3624
rect 12431 3621 12443 3624
rect 12477 3652 12489 3655
rect 13630 3652 13636 3664
rect 12477 3624 13636 3652
rect 12477 3621 12489 3624
rect 12431 3615 12489 3621
rect 13630 3612 13636 3624
rect 13688 3612 13694 3664
rect 12069 3587 12127 3593
rect 12069 3553 12081 3587
rect 12115 3584 12127 3587
rect 12158 3584 12164 3596
rect 12115 3556 12164 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 15197 3587 15255 3593
rect 15197 3553 15209 3587
rect 15243 3584 15255 3587
rect 15378 3584 15384 3596
rect 15243 3556 15384 3584
rect 15243 3553 15255 3556
rect 15197 3547 15255 3553
rect 15378 3544 15384 3556
rect 15436 3544 15442 3596
rect 13354 3380 13360 3392
rect 13315 3352 13360 3380
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 24489 3383 24547 3389
rect 24489 3349 24501 3383
rect 24535 3380 24547 3383
rect 24670 3380 24676 3392
rect 24535 3352 24676 3380
rect 24535 3349 24547 3352
rect 24489 3343 24547 3349
rect 24670 3340 24676 3352
rect 24728 3340 24734 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 11793 3179 11851 3185
rect 11793 3145 11805 3179
rect 11839 3176 11851 3179
rect 12158 3176 12164 3188
rect 11839 3148 12164 3176
rect 11839 3145 11851 3148
rect 11793 3139 11851 3145
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 13354 3108 13360 3120
rect 12820 3080 13360 3108
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12250 3040 12256 3052
rect 12207 3012 12256 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12820 3049 12848 3080
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 12805 3043 12863 3049
rect 12805 3009 12817 3043
rect 12851 3009 12863 3043
rect 13262 3040 13268 3052
rect 13223 3012 13268 3040
rect 12805 3003 12863 3009
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 12894 2904 12900 2916
rect 12855 2876 12900 2904
rect 12894 2864 12900 2876
rect 12952 2904 12958 2916
rect 13725 2907 13783 2913
rect 13725 2904 13737 2907
rect 12952 2876 13737 2904
rect 12952 2864 12958 2876
rect 13725 2873 13737 2876
rect 13771 2873 13783 2907
rect 13725 2867 13783 2873
rect 24670 2836 24676 2848
rect 24631 2808 24676 2836
rect 24670 2796 24676 2808
rect 24728 2796 24734 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12986 2632 12992 2644
rect 12483 2604 12992 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12820 2573 12848 2604
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 13354 2592 13360 2644
rect 13412 2632 13418 2644
rect 14323 2635 14381 2641
rect 14323 2632 14335 2635
rect 13412 2604 14335 2632
rect 13412 2592 13418 2604
rect 14323 2601 14335 2604
rect 14369 2601 14381 2635
rect 14323 2595 14381 2601
rect 24719 2635 24777 2641
rect 24719 2601 24731 2635
rect 24765 2632 24777 2635
rect 25222 2632 25228 2644
rect 24765 2604 25228 2632
rect 24765 2601 24777 2604
rect 24719 2595 24777 2601
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12783 2536 12817 2564
rect 12805 2533 12817 2536
rect 12851 2533 12863 2567
rect 12805 2527 12863 2533
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1854 2496 1860 2508
rect 1510 2468 1860 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 14252 2499 14310 2505
rect 14252 2465 14264 2499
rect 14298 2465 14310 2499
rect 14252 2459 14310 2465
rect 24648 2499 24706 2505
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 25130 2496 25136 2508
rect 24694 2468 25136 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 11992 2400 12725 2428
rect 11992 2369 12020 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 14267 2428 14295 2459
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 14734 2428 14740 2440
rect 14267 2400 14740 2428
rect 12713 2391 12771 2397
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 1535 2363 1593 2369
rect 1535 2329 1547 2363
rect 1581 2360 1593 2363
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 1581 2332 11989 2360
rect 1581 2329 1593 2332
rect 1535 2323 1593 2329
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 13262 2360 13268 2372
rect 13223 2332 13268 2360
rect 11977 2323 12035 2329
rect 13262 2320 13268 2332
rect 13320 2320 13326 2372
rect 25130 2292 25136 2304
rect 25091 2264 25136 2292
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 5258 76 5264 128
rect 5316 116 5322 128
rect 11974 116 11980 128
rect 5316 88 11980 116
rect 5316 76 5322 88
rect 11974 76 11980 88
rect 12032 76 12038 128
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 27160 25440 27212 25492
rect 24676 25304 24728 25356
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 25596 24896 25648 24948
rect 18880 24828 18932 24880
rect 25228 24828 25280 24880
rect 19432 24735 19484 24744
rect 19432 24701 19476 24735
rect 19476 24701 19484 24735
rect 19432 24692 19484 24701
rect 18788 24667 18840 24676
rect 18788 24633 18797 24667
rect 18797 24633 18831 24667
rect 18831 24633 18840 24667
rect 18788 24624 18840 24633
rect 20352 24624 20404 24676
rect 16948 24599 17000 24608
rect 16948 24565 16957 24599
rect 16957 24565 16991 24599
rect 16991 24565 17000 24599
rect 16948 24556 17000 24565
rect 20996 24556 21048 24608
rect 24216 24692 24268 24744
rect 23204 24556 23256 24608
rect 23756 24556 23808 24608
rect 24676 24556 24728 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 22468 24352 22520 24404
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 20628 24284 20680 24336
rect 21088 24327 21140 24336
rect 21088 24293 21097 24327
rect 21097 24293 21131 24327
rect 21131 24293 21140 24327
rect 21088 24284 21140 24293
rect 756 24216 808 24268
rect 1860 24216 1912 24268
rect 13176 24216 13228 24268
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 17408 24216 17460 24268
rect 18604 24216 18656 24268
rect 19156 24216 19208 24268
rect 22468 24259 22520 24268
rect 22468 24225 22477 24259
rect 22477 24225 22511 24259
rect 22511 24225 22520 24259
rect 22468 24216 22520 24225
rect 23848 24216 23900 24268
rect 25136 24216 25188 24268
rect 20996 24191 21048 24200
rect 20996 24157 21005 24191
rect 21005 24157 21039 24191
rect 21039 24157 21048 24191
rect 20996 24148 21048 24157
rect 21272 24191 21324 24200
rect 21272 24157 21281 24191
rect 21281 24157 21315 24191
rect 21315 24157 21324 24191
rect 21272 24148 21324 24157
rect 24124 24080 24176 24132
rect 2688 24012 2740 24064
rect 13268 24012 13320 24064
rect 19248 24012 19300 24064
rect 20444 24055 20496 24064
rect 20444 24021 20453 24055
rect 20453 24021 20487 24055
rect 20487 24021 20496 24055
rect 20444 24012 20496 24021
rect 20536 24012 20588 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1860 23851 1912 23860
rect 1860 23817 1869 23851
rect 1869 23817 1903 23851
rect 1903 23817 1912 23851
rect 1860 23808 1912 23817
rect 11704 23851 11756 23860
rect 11704 23817 11713 23851
rect 11713 23817 11747 23851
rect 11747 23817 11756 23851
rect 11704 23808 11756 23817
rect 13176 23808 13228 23860
rect 14740 23808 14792 23860
rect 15292 23808 15344 23860
rect 15568 23851 15620 23860
rect 15568 23817 15577 23851
rect 15577 23817 15611 23851
rect 15611 23817 15620 23851
rect 15568 23808 15620 23817
rect 17408 23851 17460 23860
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 17408 23808 17460 23817
rect 19156 23808 19208 23860
rect 21088 23808 21140 23860
rect 21364 23851 21416 23860
rect 21364 23817 21373 23851
rect 21373 23817 21407 23851
rect 21407 23817 21416 23851
rect 21364 23808 21416 23817
rect 23664 23808 23716 23860
rect 23848 23851 23900 23860
rect 23848 23817 23857 23851
rect 23857 23817 23891 23851
rect 23891 23817 23900 23851
rect 23848 23808 23900 23817
rect 24952 23808 25004 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 15936 23740 15988 23792
rect 17500 23740 17552 23792
rect 19340 23740 19392 23792
rect 20996 23740 21048 23792
rect 1308 23672 1360 23724
rect 16948 23672 17000 23724
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 21272 23672 21324 23724
rect 22468 23672 22520 23724
rect 11704 23604 11756 23656
rect 13544 23604 13596 23656
rect 15292 23604 15344 23656
rect 15752 23647 15804 23656
rect 15752 23613 15761 23647
rect 15761 23613 15795 23647
rect 15795 23613 15804 23647
rect 15752 23604 15804 23613
rect 16672 23604 16724 23656
rect 22008 23647 22060 23656
rect 22008 23613 22017 23647
rect 22017 23613 22051 23647
rect 22051 23613 22060 23647
rect 22008 23604 22060 23613
rect 24400 23604 24452 23656
rect 18788 23579 18840 23588
rect 1768 23468 1820 23520
rect 14740 23468 14792 23520
rect 17776 23468 17828 23520
rect 18788 23545 18797 23579
rect 18797 23545 18831 23579
rect 18831 23545 18840 23579
rect 18788 23536 18840 23545
rect 20444 23579 20496 23588
rect 20444 23545 20453 23579
rect 20453 23545 20487 23579
rect 20487 23545 20496 23579
rect 20444 23536 20496 23545
rect 20996 23468 21048 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 15568 23264 15620 23316
rect 16672 23264 16724 23316
rect 18144 23307 18196 23316
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 15752 23196 15804 23248
rect 17776 23239 17828 23248
rect 17776 23205 17785 23239
rect 17785 23205 17819 23239
rect 17819 23205 17828 23239
rect 17776 23196 17828 23205
rect 19432 23196 19484 23248
rect 19892 23196 19944 23248
rect 20536 23264 20588 23316
rect 21364 23307 21416 23316
rect 21364 23273 21373 23307
rect 21373 23273 21407 23307
rect 21407 23273 21416 23307
rect 21364 23264 21416 23273
rect 22008 23307 22060 23316
rect 22008 23273 22017 23307
rect 22017 23273 22051 23307
rect 22051 23273 22060 23307
rect 22008 23264 22060 23273
rect 24216 23264 24268 23316
rect 25504 23264 25556 23316
rect 13636 23128 13688 23180
rect 16120 23128 16172 23180
rect 17132 23171 17184 23180
rect 17132 23137 17141 23171
rect 17141 23137 17175 23171
rect 17175 23137 17184 23171
rect 17132 23128 17184 23137
rect 20996 23171 21048 23180
rect 20996 23137 21005 23171
rect 21005 23137 21039 23171
rect 21039 23137 21048 23171
rect 20996 23128 21048 23137
rect 22468 23171 22520 23180
rect 22468 23137 22477 23171
rect 22477 23137 22511 23171
rect 22511 23137 22520 23171
rect 22468 23128 22520 23137
rect 23112 23128 23164 23180
rect 24124 23128 24176 23180
rect 24676 23128 24728 23180
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 20444 22992 20496 23044
rect 12808 22924 12860 22976
rect 14556 22967 14608 22976
rect 14556 22933 14565 22967
rect 14565 22933 14599 22967
rect 14599 22933 14608 22967
rect 14556 22924 14608 22933
rect 18144 22924 18196 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 13544 22720 13596 22772
rect 19432 22720 19484 22772
rect 24676 22763 24728 22772
rect 16120 22652 16172 22704
rect 20444 22695 20496 22704
rect 20444 22661 20453 22695
rect 20453 22661 20487 22695
rect 20487 22661 20496 22695
rect 20444 22652 20496 22661
rect 14556 22627 14608 22636
rect 14556 22593 14565 22627
rect 14565 22593 14599 22627
rect 14599 22593 14608 22627
rect 14556 22584 14608 22593
rect 14740 22584 14792 22636
rect 16212 22627 16264 22636
rect 16212 22593 16221 22627
rect 16221 22593 16255 22627
rect 16255 22593 16264 22627
rect 16212 22584 16264 22593
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 19984 22584 20036 22636
rect 13084 22516 13136 22568
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 23204 22584 23256 22636
rect 25228 22559 25280 22568
rect 25228 22525 25237 22559
rect 25237 22525 25271 22559
rect 25271 22525 25280 22559
rect 25228 22516 25280 22525
rect 12808 22423 12860 22432
rect 12808 22389 12817 22423
rect 12817 22389 12851 22423
rect 12851 22389 12860 22423
rect 12808 22380 12860 22389
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 15384 22448 15436 22500
rect 14280 22380 14332 22389
rect 16396 22448 16448 22500
rect 18144 22491 18196 22500
rect 18144 22457 18153 22491
rect 18153 22457 18187 22491
rect 18187 22457 18196 22491
rect 18144 22448 18196 22457
rect 19892 22491 19944 22500
rect 17132 22423 17184 22432
rect 17132 22389 17141 22423
rect 17141 22389 17175 22423
rect 17175 22389 17184 22423
rect 17132 22380 17184 22389
rect 19892 22457 19901 22491
rect 19901 22457 19935 22491
rect 19935 22457 19944 22491
rect 19892 22448 19944 22457
rect 19984 22491 20036 22500
rect 19984 22457 19993 22491
rect 19993 22457 20027 22491
rect 20027 22457 20036 22491
rect 19984 22448 20036 22457
rect 20536 22448 20588 22500
rect 22468 22491 22520 22500
rect 22468 22457 22477 22491
rect 22477 22457 22511 22491
rect 22511 22457 22520 22491
rect 22468 22448 22520 22457
rect 23756 22491 23808 22500
rect 23756 22457 23765 22491
rect 23765 22457 23799 22491
rect 23799 22457 23808 22491
rect 23756 22448 23808 22457
rect 23848 22491 23900 22500
rect 23848 22457 23857 22491
rect 23857 22457 23891 22491
rect 23891 22457 23900 22491
rect 23848 22448 23900 22457
rect 19432 22380 19484 22432
rect 20076 22380 20128 22432
rect 20996 22380 21048 22432
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 13636 22176 13688 22228
rect 14556 22176 14608 22228
rect 15292 22176 15344 22228
rect 16212 22219 16264 22228
rect 16212 22185 16221 22219
rect 16221 22185 16255 22219
rect 16255 22185 16264 22219
rect 16212 22176 16264 22185
rect 19524 22219 19576 22228
rect 19524 22185 19533 22219
rect 19533 22185 19567 22219
rect 19567 22185 19576 22219
rect 19524 22176 19576 22185
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 18236 22108 18288 22160
rect 21088 22151 21140 22160
rect 21088 22117 21097 22151
rect 21097 22117 21131 22151
rect 21131 22117 21140 22151
rect 21088 22108 21140 22117
rect 22652 22151 22704 22160
rect 22652 22117 22661 22151
rect 22661 22117 22695 22151
rect 22695 22117 22704 22151
rect 22652 22108 22704 22117
rect 23204 22151 23256 22160
rect 23204 22117 23213 22151
rect 23213 22117 23247 22151
rect 23247 22117 23256 22151
rect 23204 22108 23256 22117
rect 23848 22108 23900 22160
rect 15476 22040 15528 22092
rect 16396 22083 16448 22092
rect 16396 22049 16405 22083
rect 16405 22049 16439 22083
rect 16439 22049 16448 22083
rect 16396 22040 16448 22049
rect 20812 22040 20864 22092
rect 24124 22083 24176 22092
rect 24124 22049 24133 22083
rect 24133 22049 24167 22083
rect 24167 22049 24176 22083
rect 24124 22040 24176 22049
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 18144 21972 18196 22024
rect 20352 21972 20404 22024
rect 22560 22015 22612 22024
rect 22560 21981 22569 22015
rect 22569 21981 22603 22015
rect 22603 21981 22612 22015
rect 22560 21972 22612 21981
rect 19156 21879 19208 21888
rect 19156 21845 19165 21879
rect 19165 21845 19199 21879
rect 19199 21845 19208 21879
rect 19156 21836 19208 21845
rect 22008 21836 22060 21888
rect 22744 21836 22796 21888
rect 23756 21836 23808 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 20076 21675 20128 21684
rect 20076 21641 20085 21675
rect 20085 21641 20119 21675
rect 20119 21641 20128 21675
rect 20076 21632 20128 21641
rect 21088 21632 21140 21684
rect 22652 21632 22704 21684
rect 24124 21675 24176 21684
rect 24124 21641 24133 21675
rect 24133 21641 24167 21675
rect 24167 21641 24176 21675
rect 24124 21632 24176 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 19708 21564 19760 21616
rect 22560 21607 22612 21616
rect 22560 21573 22569 21607
rect 22569 21573 22603 21607
rect 22603 21573 22612 21607
rect 22560 21564 22612 21573
rect 14280 21539 14332 21548
rect 14280 21505 14289 21539
rect 14289 21505 14323 21539
rect 14323 21505 14332 21539
rect 14280 21496 14332 21505
rect 17960 21496 18012 21548
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 15292 21428 15344 21480
rect 14372 21360 14424 21412
rect 15384 21360 15436 21412
rect 18052 21428 18104 21480
rect 19156 21471 19208 21480
rect 19156 21437 19165 21471
rect 19165 21437 19199 21471
rect 19199 21437 19208 21471
rect 19156 21428 19208 21437
rect 24216 21428 24268 21480
rect 14464 21292 14516 21344
rect 15476 21292 15528 21344
rect 16396 21335 16448 21344
rect 16396 21301 16405 21335
rect 16405 21301 16439 21335
rect 16439 21301 16448 21335
rect 16396 21292 16448 21301
rect 19340 21292 19392 21344
rect 20812 21292 20864 21344
rect 21456 21335 21508 21344
rect 21456 21301 21465 21335
rect 21465 21301 21499 21335
rect 21499 21301 21508 21335
rect 21456 21292 21508 21301
rect 21732 21335 21784 21344
rect 21732 21301 21741 21335
rect 21741 21301 21775 21335
rect 21775 21301 21784 21335
rect 21732 21292 21784 21301
rect 22468 21292 22520 21344
rect 22652 21292 22704 21344
rect 23020 21292 23072 21344
rect 23664 21292 23716 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 16120 21088 16172 21140
rect 16396 21088 16448 21140
rect 19432 21131 19484 21140
rect 19432 21097 19441 21131
rect 19441 21097 19475 21131
rect 19475 21097 19484 21131
rect 19432 21088 19484 21097
rect 20352 21088 20404 21140
rect 21732 21088 21784 21140
rect 22744 21131 22796 21140
rect 22744 21097 22753 21131
rect 22753 21097 22787 21131
rect 22787 21097 22796 21131
rect 22744 21088 22796 21097
rect 25504 21131 25556 21140
rect 25504 21097 25513 21131
rect 25513 21097 25547 21131
rect 25547 21097 25556 21131
rect 25504 21088 25556 21097
rect 13820 21063 13872 21072
rect 13820 21029 13829 21063
rect 13829 21029 13863 21063
rect 13863 21029 13872 21063
rect 14372 21063 14424 21072
rect 13820 21020 13872 21029
rect 14372 21029 14381 21063
rect 14381 21029 14415 21063
rect 14415 21029 14424 21063
rect 14372 21020 14424 21029
rect 19340 21020 19392 21072
rect 1124 20952 1176 21004
rect 10048 20952 10100 21004
rect 11796 20995 11848 21004
rect 11796 20961 11840 20995
rect 11840 20961 11848 20995
rect 11796 20952 11848 20961
rect 21088 20952 21140 21004
rect 23940 20995 23992 21004
rect 23940 20961 23949 20995
rect 23949 20961 23983 20995
rect 23983 20961 23992 20995
rect 23940 20952 23992 20961
rect 25136 20952 25188 21004
rect 16580 20884 16632 20936
rect 18604 20884 18656 20936
rect 24032 20884 24084 20936
rect 27620 20884 27672 20936
rect 3240 20748 3292 20800
rect 12900 20748 12952 20800
rect 13728 20748 13780 20800
rect 17408 20748 17460 20800
rect 18696 20748 18748 20800
rect 19800 20791 19852 20800
rect 19800 20757 19809 20791
rect 19809 20757 19843 20791
rect 19843 20757 19852 20791
rect 19800 20748 19852 20757
rect 24032 20791 24084 20800
rect 24032 20757 24041 20791
rect 24041 20757 24075 20791
rect 24075 20757 24084 20791
rect 24032 20748 24084 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1124 20544 1176 20596
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 11796 20587 11848 20596
rect 11796 20553 11805 20587
rect 11805 20553 11839 20587
rect 11839 20553 11848 20587
rect 11796 20544 11848 20553
rect 13820 20544 13872 20596
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 21088 20587 21140 20596
rect 21088 20553 21097 20587
rect 21097 20553 21131 20587
rect 21131 20553 21140 20587
rect 21088 20544 21140 20553
rect 22468 20587 22520 20596
rect 22468 20553 22477 20587
rect 22477 20553 22511 20587
rect 22511 20553 22520 20587
rect 22468 20544 22520 20553
rect 24032 20587 24084 20596
rect 24032 20553 24041 20587
rect 24041 20553 24075 20587
rect 24075 20553 24084 20587
rect 24032 20544 24084 20553
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 5540 20340 5592 20392
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 12992 20315 13044 20324
rect 12992 20281 13001 20315
rect 13001 20281 13035 20315
rect 13035 20281 13044 20315
rect 12992 20272 13044 20281
rect 13728 20272 13780 20324
rect 16120 20519 16172 20528
rect 16120 20485 16129 20519
rect 16129 20485 16163 20519
rect 16163 20485 16172 20519
rect 16120 20476 16172 20485
rect 16488 20476 16540 20528
rect 19340 20476 19392 20528
rect 19800 20451 19852 20460
rect 19800 20417 19809 20451
rect 19809 20417 19843 20451
rect 19843 20417 19852 20451
rect 19800 20408 19852 20417
rect 25320 20408 25372 20460
rect 16120 20340 16172 20392
rect 9680 20204 9732 20256
rect 12900 20204 12952 20256
rect 18696 20383 18748 20392
rect 18696 20349 18705 20383
rect 18705 20349 18739 20383
rect 18739 20349 18748 20383
rect 18696 20340 18748 20349
rect 21548 20383 21600 20392
rect 21548 20349 21557 20383
rect 21557 20349 21591 20383
rect 21591 20349 21600 20383
rect 21548 20340 21600 20349
rect 16488 20204 16540 20256
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 19340 20247 19392 20256
rect 19340 20213 19349 20247
rect 19349 20213 19383 20247
rect 19383 20213 19392 20247
rect 19340 20204 19392 20213
rect 23296 20204 23348 20256
rect 23940 20272 23992 20324
rect 24032 20204 24084 20256
rect 24492 20272 24544 20324
rect 25136 20204 25188 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 14372 20000 14424 20052
rect 25136 20000 25188 20052
rect 25320 20043 25372 20052
rect 25320 20009 25329 20043
rect 25329 20009 25363 20043
rect 25363 20009 25372 20043
rect 25320 20000 25372 20009
rect 18052 19975 18104 19984
rect 18052 19941 18061 19975
rect 18061 19941 18095 19975
rect 18095 19941 18104 19975
rect 18052 19932 18104 19941
rect 18696 19932 18748 19984
rect 12992 19864 13044 19916
rect 13176 19864 13228 19916
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 15844 19864 15896 19916
rect 17776 19907 17828 19916
rect 15936 19796 15988 19848
rect 17776 19873 17785 19907
rect 17785 19873 17819 19907
rect 17819 19873 17828 19907
rect 17776 19864 17828 19873
rect 21548 19932 21600 19984
rect 22376 19975 22428 19984
rect 22376 19941 22385 19975
rect 22385 19941 22419 19975
rect 22419 19941 22428 19975
rect 22376 19932 22428 19941
rect 23940 19975 23992 19984
rect 23940 19941 23949 19975
rect 23949 19941 23983 19975
rect 23983 19941 23992 19975
rect 23940 19932 23992 19941
rect 24492 19975 24544 19984
rect 24492 19941 24501 19975
rect 24501 19941 24535 19975
rect 24535 19941 24544 19975
rect 24492 19932 24544 19941
rect 20076 19864 20128 19916
rect 21916 19864 21968 19916
rect 22284 19839 22336 19848
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 24032 19796 24084 19848
rect 23112 19728 23164 19780
rect 23664 19728 23716 19780
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 13636 19703 13688 19712
rect 13636 19669 13645 19703
rect 13645 19669 13679 19703
rect 13679 19669 13688 19703
rect 13636 19660 13688 19669
rect 16580 19660 16632 19712
rect 18604 19660 18656 19712
rect 19156 19660 19208 19712
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 24492 19728 24544 19780
rect 23204 19660 23256 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 16580 19499 16632 19508
rect 16580 19465 16589 19499
rect 16589 19465 16623 19499
rect 16623 19465 16632 19499
rect 20076 19499 20128 19508
rect 16580 19456 16632 19465
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 25412 19499 25464 19508
rect 25412 19465 25421 19499
rect 25421 19465 25455 19499
rect 25455 19465 25464 19499
rect 25412 19456 25464 19465
rect 24216 19388 24268 19440
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 22284 19320 22336 19372
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 17776 19295 17828 19304
rect 12624 19184 12676 19236
rect 12900 19227 12952 19236
rect 12900 19193 12909 19227
rect 12909 19193 12943 19227
rect 12943 19193 12952 19227
rect 12900 19184 12952 19193
rect 14832 19184 14884 19236
rect 15292 19227 15344 19236
rect 15292 19193 15301 19227
rect 15301 19193 15335 19227
rect 15335 19193 15344 19227
rect 15292 19184 15344 19193
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 17776 19252 17828 19261
rect 18512 19252 18564 19304
rect 19156 19295 19208 19304
rect 17868 19184 17920 19236
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 20628 19252 20680 19304
rect 23204 19252 23256 19304
rect 25228 19295 25280 19304
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 13176 19116 13228 19168
rect 15844 19116 15896 19168
rect 18052 19116 18104 19168
rect 19340 19184 19392 19236
rect 22100 19184 22152 19236
rect 23756 19227 23808 19236
rect 23756 19193 23765 19227
rect 23765 19193 23799 19227
rect 23799 19193 23808 19227
rect 23756 19184 23808 19193
rect 18696 19116 18748 19168
rect 20996 19116 21048 19168
rect 22376 19116 22428 19168
rect 23388 19159 23440 19168
rect 23388 19125 23397 19159
rect 23397 19125 23431 19159
rect 23431 19125 23440 19159
rect 23388 19116 23440 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 13176 18955 13228 18964
rect 13176 18921 13185 18955
rect 13185 18921 13219 18955
rect 13219 18921 13228 18955
rect 13176 18912 13228 18921
rect 15936 18912 15988 18964
rect 16120 18955 16172 18964
rect 16120 18921 16129 18955
rect 16129 18921 16163 18955
rect 16163 18921 16172 18955
rect 16120 18912 16172 18921
rect 20628 18955 20680 18964
rect 20628 18921 20637 18955
rect 20637 18921 20671 18955
rect 20671 18921 20680 18955
rect 20628 18912 20680 18921
rect 21916 18955 21968 18964
rect 21916 18921 21925 18955
rect 21925 18921 21959 18955
rect 21959 18921 21968 18955
rect 21916 18912 21968 18921
rect 23296 18912 23348 18964
rect 24860 18912 24912 18964
rect 13636 18844 13688 18896
rect 15568 18776 15620 18828
rect 22284 18844 22336 18896
rect 18696 18819 18748 18828
rect 13728 18708 13780 18760
rect 18696 18785 18705 18819
rect 18705 18785 18739 18819
rect 18739 18785 18748 18819
rect 18696 18776 18748 18785
rect 19156 18819 19208 18828
rect 19156 18785 19165 18819
rect 19165 18785 19199 18819
rect 19199 18785 19208 18819
rect 19156 18776 19208 18785
rect 20996 18819 21048 18828
rect 20996 18785 21005 18819
rect 21005 18785 21039 18819
rect 21039 18785 21048 18819
rect 20996 18776 21048 18785
rect 23388 18776 23440 18828
rect 24216 18776 24268 18828
rect 15844 18640 15896 18692
rect 22836 18708 22888 18760
rect 14004 18572 14056 18624
rect 15568 18615 15620 18624
rect 15568 18581 15577 18615
rect 15577 18581 15611 18615
rect 15611 18581 15620 18615
rect 15568 18572 15620 18581
rect 23756 18572 23808 18624
rect 25044 18572 25096 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3792 18368 3844 18420
rect 13636 18411 13688 18420
rect 13636 18377 13645 18411
rect 13645 18377 13679 18411
rect 13679 18377 13688 18411
rect 13636 18368 13688 18377
rect 18696 18368 18748 18420
rect 20996 18368 21048 18420
rect 22836 18411 22888 18420
rect 22836 18377 22845 18411
rect 22845 18377 22879 18411
rect 22879 18377 22888 18411
rect 22836 18368 22888 18377
rect 24768 18411 24820 18420
rect 24768 18377 24777 18411
rect 24777 18377 24811 18411
rect 24811 18377 24820 18411
rect 24768 18368 24820 18377
rect 15936 18275 15988 18284
rect 15936 18241 15945 18275
rect 15945 18241 15979 18275
rect 15979 18241 15988 18275
rect 15936 18232 15988 18241
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 21916 18275 21968 18284
rect 21916 18241 21925 18275
rect 21925 18241 21959 18275
rect 21959 18241 21968 18275
rect 21916 18232 21968 18241
rect 3792 18164 3844 18216
rect 14832 18164 14884 18216
rect 12992 18096 13044 18148
rect 3884 18028 3936 18080
rect 14004 18071 14056 18080
rect 14004 18037 14013 18071
rect 14013 18037 14047 18071
rect 14047 18037 14056 18071
rect 14004 18028 14056 18037
rect 14832 18071 14884 18080
rect 14832 18037 14841 18071
rect 14841 18037 14875 18071
rect 14875 18037 14884 18071
rect 14832 18028 14884 18037
rect 15200 18096 15252 18148
rect 17040 18164 17092 18216
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 18788 18096 18840 18148
rect 19156 18096 19208 18148
rect 15568 18028 15620 18080
rect 17776 18071 17828 18080
rect 17776 18037 17785 18071
rect 17785 18037 17819 18071
rect 17819 18037 17828 18071
rect 17776 18028 17828 18037
rect 22008 18096 22060 18148
rect 22284 18028 22336 18080
rect 24216 18028 24268 18080
rect 24860 18028 24912 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 14004 17824 14056 17876
rect 15200 17756 15252 17808
rect 20720 17756 20772 17808
rect 21916 17756 21968 17808
rect 22008 17756 22060 17808
rect 1124 17688 1176 17740
rect 16120 17731 16172 17740
rect 16120 17697 16129 17731
rect 16129 17697 16163 17731
rect 16163 17697 16172 17731
rect 16120 17688 16172 17697
rect 18880 17688 18932 17740
rect 19984 17688 20036 17740
rect 22560 17731 22612 17740
rect 22560 17697 22569 17731
rect 22569 17697 22603 17731
rect 22603 17697 22612 17731
rect 22560 17688 22612 17697
rect 24952 17688 25004 17740
rect 17592 17663 17644 17672
rect 17592 17629 17601 17663
rect 17601 17629 17635 17663
rect 17635 17629 17644 17663
rect 17592 17620 17644 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 24032 17663 24084 17672
rect 24032 17629 24041 17663
rect 24041 17629 24075 17663
rect 24075 17629 24084 17663
rect 24032 17620 24084 17629
rect 8944 17484 8996 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 16304 17527 16356 17536
rect 16304 17493 16313 17527
rect 16313 17493 16347 17527
rect 16347 17493 16356 17527
rect 16304 17484 16356 17493
rect 16488 17484 16540 17536
rect 18512 17484 18564 17536
rect 19432 17527 19484 17536
rect 19432 17493 19441 17527
rect 19441 17493 19475 17527
rect 19475 17493 19484 17527
rect 19432 17484 19484 17493
rect 25228 17552 25280 17604
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1124 17280 1176 17332
rect 2412 17323 2464 17332
rect 2412 17289 2421 17323
rect 2421 17289 2455 17323
rect 2455 17289 2464 17323
rect 2412 17280 2464 17289
rect 16120 17280 16172 17332
rect 16304 17280 16356 17332
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 22284 17280 22336 17332
rect 22560 17323 22612 17332
rect 22560 17289 22569 17323
rect 22569 17289 22603 17323
rect 22603 17289 22612 17323
rect 22560 17280 22612 17289
rect 24032 17280 24084 17332
rect 17500 17212 17552 17264
rect 19984 17212 20036 17264
rect 24768 17212 24820 17264
rect 16396 17187 16448 17196
rect 16396 17153 16405 17187
rect 16405 17153 16439 17187
rect 16439 17153 16448 17187
rect 16396 17144 16448 17153
rect 17592 17144 17644 17196
rect 20996 17144 21048 17196
rect 21640 17144 21692 17196
rect 24124 17187 24176 17196
rect 24124 17153 24133 17187
rect 24133 17153 24167 17187
rect 24167 17153 24176 17187
rect 24124 17144 24176 17153
rect 2412 17076 2464 17128
rect 12900 17076 12952 17128
rect 15384 17119 15436 17128
rect 15384 17085 15393 17119
rect 15393 17085 15427 17119
rect 15427 17085 15436 17119
rect 15384 17076 15436 17085
rect 19064 17076 19116 17128
rect 19432 17119 19484 17128
rect 19432 17085 19441 17119
rect 19441 17085 19475 17119
rect 19475 17085 19484 17119
rect 19432 17076 19484 17085
rect 22560 17076 22612 17128
rect 23020 17076 23072 17128
rect 15476 17051 15528 17060
rect 15476 17017 15485 17051
rect 15485 17017 15519 17051
rect 15519 17017 15528 17051
rect 15476 17008 15528 17017
rect 19340 17051 19392 17060
rect 1952 16940 2004 16992
rect 12992 16983 13044 16992
rect 12992 16949 13001 16983
rect 13001 16949 13035 16983
rect 13035 16949 13044 16983
rect 12992 16940 13044 16949
rect 16304 16940 16356 16992
rect 19340 17017 19349 17051
rect 19349 17017 19383 17051
rect 19383 17017 19392 17051
rect 19340 17008 19392 17017
rect 21272 17051 21324 17060
rect 21272 17017 21281 17051
rect 21281 17017 21315 17051
rect 21315 17017 21324 17051
rect 21272 17008 21324 17017
rect 18880 16983 18932 16992
rect 18880 16949 18889 16983
rect 18889 16949 18923 16983
rect 18923 16949 18932 16983
rect 18880 16940 18932 16949
rect 20536 16940 20588 16992
rect 23388 16983 23440 16992
rect 23388 16949 23397 16983
rect 23397 16949 23431 16983
rect 23431 16949 23440 16983
rect 23388 16940 23440 16949
rect 24032 16940 24084 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 16396 16779 16448 16788
rect 16396 16745 16405 16779
rect 16405 16745 16439 16779
rect 16439 16745 16448 16779
rect 16396 16736 16448 16745
rect 19984 16736 20036 16788
rect 20996 16736 21048 16788
rect 21272 16736 21324 16788
rect 24124 16779 24176 16788
rect 24124 16745 24133 16779
rect 24133 16745 24167 16779
rect 24167 16745 24176 16779
rect 24124 16736 24176 16745
rect 12992 16711 13044 16720
rect 12992 16677 13001 16711
rect 13001 16677 13035 16711
rect 13035 16677 13044 16711
rect 12992 16668 13044 16677
rect 13544 16711 13596 16720
rect 13544 16677 13553 16711
rect 13553 16677 13587 16711
rect 13587 16677 13596 16711
rect 13544 16668 13596 16677
rect 15384 16668 15436 16720
rect 16120 16668 16172 16720
rect 16948 16668 17000 16720
rect 19340 16668 19392 16720
rect 21088 16711 21140 16720
rect 21088 16677 21097 16711
rect 21097 16677 21131 16711
rect 21131 16677 21140 16711
rect 21088 16668 21140 16677
rect 21640 16711 21692 16720
rect 21640 16677 21649 16711
rect 21649 16677 21683 16711
rect 21683 16677 21692 16711
rect 21640 16668 21692 16677
rect 22468 16668 22520 16720
rect 23388 16668 23440 16720
rect 24952 16668 25004 16720
rect 12256 16532 12308 16584
rect 14740 16532 14792 16584
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 21364 16532 21416 16584
rect 22928 16575 22980 16584
rect 22928 16541 22937 16575
rect 22937 16541 22971 16575
rect 22971 16541 22980 16575
rect 22928 16532 22980 16541
rect 24768 16575 24820 16584
rect 17500 16507 17552 16516
rect 17500 16473 17509 16507
rect 17509 16473 17543 16507
rect 17543 16473 17552 16507
rect 17500 16464 17552 16473
rect 20536 16464 20588 16516
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 24676 16464 24728 16516
rect 15844 16396 15896 16448
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 12256 16235 12308 16244
rect 12256 16201 12265 16235
rect 12265 16201 12299 16235
rect 12299 16201 12308 16235
rect 12256 16192 12308 16201
rect 12992 16192 13044 16244
rect 14740 16235 14792 16244
rect 14740 16201 14749 16235
rect 14749 16201 14783 16235
rect 14783 16201 14792 16235
rect 14740 16192 14792 16201
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 16948 16235 17000 16244
rect 16948 16201 16957 16235
rect 16957 16201 16991 16235
rect 16991 16201 17000 16235
rect 16948 16192 17000 16201
rect 19340 16235 19392 16244
rect 19340 16201 19349 16235
rect 19349 16201 19383 16235
rect 19383 16201 19392 16235
rect 19340 16192 19392 16201
rect 24216 16192 24268 16244
rect 24952 16192 25004 16244
rect 25044 16192 25096 16244
rect 22468 16167 22520 16176
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 16028 16099 16080 16108
rect 16028 16065 16037 16099
rect 16037 16065 16071 16099
rect 16071 16065 16080 16099
rect 16028 16056 16080 16065
rect 12900 15963 12952 15972
rect 12900 15929 12909 15963
rect 12909 15929 12943 15963
rect 12943 15929 12952 15963
rect 12900 15920 12952 15929
rect 12992 15963 13044 15972
rect 12992 15929 13001 15963
rect 13001 15929 13035 15963
rect 13035 15929 13044 15963
rect 12992 15920 13044 15929
rect 15384 15852 15436 15904
rect 15476 15852 15528 15904
rect 22468 16133 22477 16167
rect 22477 16133 22511 16167
rect 22511 16133 22520 16167
rect 22468 16124 22520 16133
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 21088 16056 21140 16108
rect 21364 16099 21416 16108
rect 21364 16065 21373 16099
rect 21373 16065 21407 16099
rect 21407 16065 21416 16099
rect 21364 16056 21416 16065
rect 25228 16056 25280 16108
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 20536 16031 20588 16040
rect 20536 15997 20545 16031
rect 20545 15997 20579 16031
rect 20579 15997 20588 16031
rect 20536 15988 20588 15997
rect 17684 15852 17736 15904
rect 18512 15852 18564 15904
rect 23940 15963 23992 15972
rect 23940 15929 23949 15963
rect 23949 15929 23983 15963
rect 23983 15929 23992 15963
rect 24492 15963 24544 15972
rect 23940 15920 23992 15929
rect 24492 15929 24501 15963
rect 24501 15929 24535 15963
rect 24535 15929 24544 15963
rect 24492 15920 24544 15929
rect 22192 15852 22244 15904
rect 23112 15895 23164 15904
rect 23112 15861 23121 15895
rect 23121 15861 23155 15895
rect 23155 15861 23164 15895
rect 23112 15852 23164 15861
rect 25228 15895 25280 15904
rect 25228 15861 25237 15895
rect 25237 15861 25271 15895
rect 25271 15861 25280 15895
rect 25228 15852 25280 15861
rect 25872 15895 25924 15904
rect 25872 15861 25881 15895
rect 25881 15861 25915 15895
rect 25915 15861 25924 15895
rect 25872 15852 25924 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 12624 15691 12676 15700
rect 12624 15657 12633 15691
rect 12633 15657 12667 15691
rect 12667 15657 12676 15691
rect 12624 15648 12676 15657
rect 12900 15648 12952 15700
rect 15844 15648 15896 15700
rect 16028 15648 16080 15700
rect 17868 15691 17920 15700
rect 17868 15657 17877 15691
rect 17877 15657 17911 15691
rect 17911 15657 17920 15691
rect 17868 15648 17920 15657
rect 23388 15648 23440 15700
rect 24492 15648 24544 15700
rect 15936 15580 15988 15632
rect 22284 15580 22336 15632
rect 22928 15580 22980 15632
rect 23940 15580 23992 15632
rect 12992 15512 13044 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 16120 15512 16172 15564
rect 16948 15512 17000 15564
rect 18328 15555 18380 15564
rect 18328 15521 18337 15555
rect 18337 15521 18371 15555
rect 18371 15521 18380 15555
rect 18328 15512 18380 15521
rect 18512 15555 18564 15564
rect 18512 15521 18521 15555
rect 18521 15521 18555 15555
rect 18555 15521 18564 15555
rect 18512 15512 18564 15521
rect 24768 15555 24820 15564
rect 24768 15521 24777 15555
rect 24777 15521 24811 15555
rect 24811 15521 24820 15555
rect 24768 15512 24820 15521
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 18604 15487 18656 15496
rect 18604 15453 18613 15487
rect 18613 15453 18647 15487
rect 18647 15453 18656 15487
rect 18604 15444 18656 15453
rect 22376 15487 22428 15496
rect 22376 15453 22385 15487
rect 22385 15453 22419 15487
rect 22419 15453 22428 15487
rect 22376 15444 22428 15453
rect 17776 15376 17828 15428
rect 18328 15376 18380 15428
rect 16580 15351 16632 15360
rect 16580 15317 16589 15351
rect 16589 15317 16623 15351
rect 16623 15317 16632 15351
rect 16580 15308 16632 15317
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 21640 15308 21692 15360
rect 24216 15308 24268 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 12164 15104 12216 15156
rect 12624 15104 12676 15156
rect 15384 15104 15436 15156
rect 15936 15147 15988 15156
rect 15936 15113 15945 15147
rect 15945 15113 15979 15147
rect 15979 15113 15988 15147
rect 15936 15104 15988 15113
rect 18144 15104 18196 15156
rect 18328 15104 18380 15156
rect 22468 15104 22520 15156
rect 24768 15104 24820 15156
rect 11520 14968 11572 15020
rect 12624 14968 12676 15020
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 18880 14968 18932 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20444 15011 20496 15020
rect 20444 14977 20453 15011
rect 20453 14977 20487 15011
rect 20487 14977 20496 15011
rect 20444 14968 20496 14977
rect 5448 14943 5500 14952
rect 5448 14909 5466 14943
rect 5466 14909 5500 14943
rect 5448 14900 5500 14909
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 12624 14875 12676 14884
rect 12624 14841 12633 14875
rect 12633 14841 12667 14875
rect 12667 14841 12676 14875
rect 15936 14900 15988 14952
rect 16580 14943 16632 14952
rect 16580 14909 16589 14943
rect 16589 14909 16623 14943
rect 16623 14909 16632 14943
rect 16580 14900 16632 14909
rect 17868 14900 17920 14952
rect 12624 14832 12676 14841
rect 15292 14832 15344 14884
rect 21640 14900 21692 14952
rect 24216 14943 24268 14952
rect 24216 14909 24225 14943
rect 24225 14909 24259 14943
rect 24259 14909 24268 14943
rect 24216 14900 24268 14909
rect 18328 14875 18380 14884
rect 18328 14841 18337 14875
rect 18337 14841 18371 14875
rect 18371 14841 18380 14875
rect 18328 14832 18380 14841
rect 19064 14832 19116 14884
rect 20076 14875 20128 14884
rect 20076 14841 20085 14875
rect 20085 14841 20119 14875
rect 20119 14841 20128 14875
rect 20076 14832 20128 14841
rect 22284 14832 22336 14884
rect 24676 14875 24728 14884
rect 24676 14841 24685 14875
rect 24685 14841 24719 14875
rect 24719 14841 24728 14875
rect 24676 14832 24728 14841
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 15660 14764 15712 14816
rect 16948 14764 17000 14816
rect 18512 14764 18564 14816
rect 24492 14764 24544 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 16580 14560 16632 14612
rect 18236 14560 18288 14612
rect 19984 14560 20036 14612
rect 22376 14603 22428 14612
rect 22376 14569 22385 14603
rect 22385 14569 22419 14603
rect 22419 14569 22428 14603
rect 22376 14560 22428 14569
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 14188 14467 14240 14476
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 18144 14492 18196 14544
rect 19340 14492 19392 14544
rect 20076 14492 20128 14544
rect 22928 14492 22980 14544
rect 24032 14492 24084 14544
rect 24492 14535 24544 14544
rect 24492 14501 24501 14535
rect 24501 14501 24535 14535
rect 24535 14501 24544 14535
rect 24492 14492 24544 14501
rect 24676 14492 24728 14544
rect 17408 14424 17460 14476
rect 21548 14467 21600 14476
rect 21548 14433 21557 14467
rect 21557 14433 21591 14467
rect 21591 14433 21600 14467
rect 21548 14424 21600 14433
rect 11796 14356 11848 14408
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 17132 14356 17184 14408
rect 22744 14356 22796 14408
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 23572 14356 23624 14365
rect 23664 14356 23716 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 13544 14288 13596 14340
rect 16396 14288 16448 14340
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 19524 14220 19576 14272
rect 24216 14263 24268 14272
rect 24216 14229 24225 14263
rect 24225 14229 24259 14263
rect 24259 14229 24268 14263
rect 24216 14220 24268 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 11520 14016 11572 14068
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 12624 14016 12676 14068
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 18144 14016 18196 14068
rect 18236 14016 18288 14068
rect 21548 14016 21600 14068
rect 22744 14016 22796 14068
rect 24032 14059 24084 14068
rect 24032 14025 24041 14059
rect 24041 14025 24075 14059
rect 24075 14025 24084 14059
rect 24032 14016 24084 14025
rect 24676 14016 24728 14068
rect 20444 13991 20496 14000
rect 20444 13957 20453 13991
rect 20453 13957 20487 13991
rect 20487 13957 20496 13991
rect 20444 13948 20496 13957
rect 12256 13880 12308 13932
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 22376 13948 22428 14000
rect 24768 13991 24820 14000
rect 24768 13957 24777 13991
rect 24777 13957 24811 13991
rect 24811 13957 24820 13991
rect 24768 13948 24820 13957
rect 17132 13880 17184 13889
rect 23572 13880 23624 13932
rect 24584 13880 24636 13932
rect 12532 13812 12584 13864
rect 14372 13812 14424 13864
rect 14832 13812 14884 13864
rect 16396 13855 16448 13864
rect 16396 13821 16405 13855
rect 16405 13821 16439 13855
rect 16439 13821 16448 13855
rect 16396 13812 16448 13821
rect 16488 13812 16540 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 21824 13855 21876 13864
rect 18144 13744 18196 13796
rect 19064 13744 19116 13796
rect 19340 13744 19392 13796
rect 12164 13719 12216 13728
rect 12164 13685 12173 13719
rect 12173 13685 12207 13719
rect 12207 13685 12216 13719
rect 12164 13676 12216 13685
rect 13544 13676 13596 13728
rect 15660 13676 15712 13728
rect 19524 13676 19576 13728
rect 21548 13744 21600 13796
rect 20628 13676 20680 13728
rect 21180 13719 21232 13728
rect 21180 13685 21189 13719
rect 21189 13685 21223 13719
rect 21223 13685 21232 13719
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 24308 13787 24360 13796
rect 24308 13753 24317 13787
rect 24317 13753 24351 13787
rect 24351 13753 24360 13787
rect 24308 13744 24360 13753
rect 22836 13719 22888 13728
rect 21180 13676 21232 13685
rect 22836 13685 22845 13719
rect 22845 13685 22879 13719
rect 22879 13685 22888 13719
rect 22836 13676 22888 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 12348 13515 12400 13524
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 18144 13515 18196 13524
rect 14648 13404 14700 13456
rect 18144 13481 18153 13515
rect 18153 13481 18187 13515
rect 18187 13481 18196 13515
rect 18144 13472 18196 13481
rect 22744 13472 22796 13524
rect 24308 13472 24360 13524
rect 18052 13404 18104 13456
rect 18880 13404 18932 13456
rect 21640 13447 21692 13456
rect 21640 13413 21649 13447
rect 21649 13413 21683 13447
rect 21683 13413 21692 13447
rect 21640 13404 21692 13413
rect 24676 13404 24728 13456
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 12624 13379 12676 13388
rect 12624 13345 12633 13379
rect 12633 13345 12667 13379
rect 12667 13345 12676 13379
rect 12624 13336 12676 13345
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 14832 13336 14884 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 16672 13379 16724 13388
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 16856 13336 16908 13388
rect 20352 13336 20404 13388
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19340 13311 19392 13320
rect 19340 13277 19349 13311
rect 19349 13277 19383 13311
rect 19383 13277 19392 13311
rect 19340 13268 19392 13277
rect 20628 13268 20680 13320
rect 21824 13336 21876 13388
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 24584 13311 24636 13320
rect 16396 13200 16448 13252
rect 21180 13200 21232 13252
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 25136 13200 25188 13252
rect 12532 13132 12584 13184
rect 13452 13175 13504 13184
rect 13452 13141 13461 13175
rect 13461 13141 13495 13175
rect 13495 13141 13504 13175
rect 13452 13132 13504 13141
rect 14832 13175 14884 13184
rect 14832 13141 14841 13175
rect 14841 13141 14875 13175
rect 14875 13141 14884 13175
rect 14832 13132 14884 13141
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 21916 13175 21968 13184
rect 21916 13141 21925 13175
rect 21925 13141 21959 13175
rect 21959 13141 21968 13175
rect 21916 13132 21968 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 11796 12928 11848 12980
rect 13912 12928 13964 12980
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 16856 12928 16908 12980
rect 18880 12928 18932 12980
rect 22836 12928 22888 12980
rect 12256 12860 12308 12912
rect 12808 12860 12860 12912
rect 16120 12860 16172 12912
rect 16488 12860 16540 12912
rect 19064 12860 19116 12912
rect 25412 12860 25464 12912
rect 13452 12792 13504 12844
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 16580 12792 16632 12844
rect 21916 12792 21968 12844
rect 24676 12835 24728 12844
rect 24676 12801 24685 12835
rect 24685 12801 24719 12835
rect 24719 12801 24728 12835
rect 24676 12792 24728 12801
rect 11980 12724 12032 12776
rect 13360 12724 13412 12776
rect 14740 12724 14792 12776
rect 17960 12724 18012 12776
rect 11888 12588 11940 12640
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 16672 12656 16724 12708
rect 20352 12724 20404 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 22836 12724 22888 12776
rect 15016 12631 15068 12640
rect 13360 12588 13412 12597
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 16580 12588 16632 12640
rect 17960 12588 18012 12640
rect 18604 12588 18656 12640
rect 21640 12631 21692 12640
rect 21640 12597 21649 12631
rect 21649 12597 21683 12631
rect 21683 12597 21692 12631
rect 21640 12588 21692 12597
rect 22744 12588 22796 12640
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 14740 12427 14792 12436
rect 14740 12393 14749 12427
rect 14749 12393 14783 12427
rect 14783 12393 14792 12427
rect 14740 12384 14792 12393
rect 15016 12384 15068 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 12532 12359 12584 12368
rect 12532 12325 12541 12359
rect 12541 12325 12575 12359
rect 12575 12325 12584 12359
rect 12532 12316 12584 12325
rect 13452 12316 13504 12368
rect 15568 12316 15620 12368
rect 16488 12316 16540 12368
rect 17500 12384 17552 12436
rect 25228 12384 25280 12436
rect 18696 12316 18748 12368
rect 22468 12359 22520 12368
rect 22468 12325 22477 12359
rect 22477 12325 22511 12359
rect 22511 12325 22520 12359
rect 22468 12316 22520 12325
rect 27620 12316 27672 12368
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 11888 12248 11940 12300
rect 12624 12248 12676 12300
rect 13084 12248 13136 12300
rect 16672 12248 16724 12300
rect 18144 12291 18196 12300
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 12992 12044 13044 12096
rect 13912 12223 13964 12232
rect 13912 12189 13921 12223
rect 13921 12189 13955 12223
rect 13955 12189 13964 12223
rect 13912 12180 13964 12189
rect 16580 12180 16632 12232
rect 18144 12257 18153 12291
rect 18153 12257 18187 12291
rect 18187 12257 18196 12291
rect 18144 12248 18196 12257
rect 19064 12248 19116 12300
rect 21180 12291 21232 12300
rect 21180 12257 21189 12291
rect 21189 12257 21223 12291
rect 21223 12257 21232 12291
rect 21180 12248 21232 12257
rect 18604 12180 18656 12232
rect 24768 12248 24820 12300
rect 25504 12291 25556 12300
rect 25504 12257 25522 12291
rect 25522 12257 25556 12291
rect 25504 12248 25556 12257
rect 16856 12112 16908 12164
rect 20720 12112 20772 12164
rect 14740 12044 14792 12096
rect 15660 12044 15712 12096
rect 18052 12087 18104 12096
rect 18052 12053 18061 12087
rect 18061 12053 18095 12087
rect 18095 12053 18104 12087
rect 18052 12044 18104 12053
rect 19156 12087 19208 12096
rect 19156 12053 19165 12087
rect 19165 12053 19199 12087
rect 19199 12053 19208 12087
rect 19156 12044 19208 12053
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 24124 12087 24176 12096
rect 24124 12053 24133 12087
rect 24133 12053 24167 12087
rect 24167 12053 24176 12087
rect 24124 12044 24176 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 11796 11883 11848 11892
rect 11796 11849 11805 11883
rect 11805 11849 11839 11883
rect 11839 11849 11848 11883
rect 11796 11840 11848 11849
rect 14813 11883 14865 11892
rect 14813 11849 14822 11883
rect 14822 11849 14856 11883
rect 14856 11849 14865 11883
rect 16488 11883 16540 11892
rect 14813 11840 14865 11849
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 16856 11883 16908 11892
rect 16856 11849 16865 11883
rect 16865 11849 16899 11883
rect 16899 11849 16908 11883
rect 16856 11840 16908 11849
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 21180 11840 21232 11892
rect 24124 11883 24176 11892
rect 24124 11849 24133 11883
rect 24133 11849 24167 11883
rect 24167 11849 24176 11883
rect 24124 11840 24176 11849
rect 25504 11883 25556 11892
rect 25504 11849 25513 11883
rect 25513 11849 25547 11883
rect 25547 11849 25556 11883
rect 25504 11840 25556 11849
rect 13452 11772 13504 11824
rect 15384 11772 15436 11824
rect 17776 11772 17828 11824
rect 18604 11772 18656 11824
rect 13360 11704 13412 11756
rect 16580 11747 16632 11756
rect 16580 11713 16589 11747
rect 16589 11713 16623 11747
rect 16623 11713 16632 11747
rect 16580 11704 16632 11713
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 22192 11704 22244 11756
rect 24952 11704 25004 11756
rect 12808 11636 12860 11688
rect 13636 11636 13688 11688
rect 13084 11568 13136 11620
rect 14648 11611 14700 11620
rect 14648 11577 14657 11611
rect 14657 11577 14691 11611
rect 14691 11577 14700 11611
rect 14648 11568 14700 11577
rect 15568 11568 15620 11620
rect 12164 11500 12216 11552
rect 12532 11500 12584 11552
rect 15384 11500 15436 11552
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 17868 11636 17920 11688
rect 19156 11636 19208 11688
rect 20352 11636 20404 11688
rect 20720 11636 20772 11688
rect 21272 11611 21324 11620
rect 17776 11543 17828 11552
rect 16120 11500 16172 11509
rect 17776 11509 17785 11543
rect 17785 11509 17819 11543
rect 17819 11509 17828 11543
rect 17776 11500 17828 11509
rect 21272 11577 21281 11611
rect 21281 11577 21315 11611
rect 21315 11577 21324 11611
rect 21272 11568 21324 11577
rect 24308 11611 24360 11620
rect 24308 11577 24317 11611
rect 24317 11577 24351 11611
rect 24351 11577 24360 11611
rect 24308 11568 24360 11577
rect 18144 11500 18196 11552
rect 23388 11543 23440 11552
rect 23388 11509 23397 11543
rect 23397 11509 23431 11543
rect 23431 11509 23440 11543
rect 23388 11500 23440 11509
rect 24124 11500 24176 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 13084 11296 13136 11348
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 20812 11296 20864 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 23020 11296 23072 11348
rect 24308 11339 24360 11348
rect 12256 11228 12308 11280
rect 12348 11228 12400 11280
rect 1308 11160 1360 11212
rect 15568 11228 15620 11280
rect 20628 11228 20680 11280
rect 23112 11271 23164 11280
rect 23112 11237 23121 11271
rect 23121 11237 23155 11271
rect 23155 11237 23164 11271
rect 23112 11228 23164 11237
rect 24308 11305 24317 11339
rect 24317 11305 24351 11339
rect 24351 11305 24360 11339
rect 24308 11296 24360 11305
rect 24768 11271 24820 11280
rect 24768 11237 24777 11271
rect 24777 11237 24811 11271
rect 24811 11237 24820 11271
rect 24768 11228 24820 11237
rect 13636 11160 13688 11212
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 16028 11160 16080 11212
rect 18328 11203 18380 11212
rect 18328 11169 18337 11203
rect 18337 11169 18371 11203
rect 18371 11169 18380 11203
rect 18328 11160 18380 11169
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12992 11092 13044 11144
rect 13728 11092 13780 11144
rect 16672 11092 16724 11144
rect 17960 11092 18012 11144
rect 19156 11092 19208 11144
rect 21272 11135 21324 11144
rect 21272 11101 21281 11135
rect 21281 11101 21315 11135
rect 21315 11101 21324 11135
rect 21272 11092 21324 11101
rect 24032 11092 24084 11144
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 15384 10956 15436 11008
rect 16580 10956 16632 11008
rect 17132 10956 17184 11008
rect 17868 10999 17920 11008
rect 17868 10965 17877 10999
rect 17877 10965 17911 10999
rect 17911 10965 17920 10999
rect 17868 10956 17920 10965
rect 18144 10999 18196 11008
rect 18144 10965 18153 10999
rect 18153 10965 18187 10999
rect 18187 10965 18196 10999
rect 18144 10956 18196 10965
rect 18696 10956 18748 11008
rect 20720 10956 20772 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1308 10752 1360 10804
rect 13636 10795 13688 10804
rect 13636 10761 13645 10795
rect 13645 10761 13679 10795
rect 13679 10761 13688 10795
rect 13636 10752 13688 10761
rect 14096 10752 14148 10804
rect 17776 10752 17828 10804
rect 18788 10752 18840 10804
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 24768 10795 24820 10804
rect 24768 10761 24777 10795
rect 24777 10761 24811 10795
rect 24811 10761 24820 10795
rect 24768 10752 24820 10761
rect 11796 10684 11848 10736
rect 12532 10684 12584 10736
rect 14740 10684 14792 10736
rect 16488 10684 16540 10736
rect 17132 10727 17184 10736
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 17868 10684 17920 10736
rect 23388 10684 23440 10736
rect 25780 10727 25832 10736
rect 25780 10693 25789 10727
rect 25789 10693 25823 10727
rect 25823 10693 25832 10727
rect 25780 10684 25832 10693
rect 10876 10548 10928 10600
rect 13728 10616 13780 10668
rect 14832 10616 14884 10668
rect 15476 10616 15528 10668
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 14372 10548 14424 10600
rect 15568 10548 15620 10600
rect 16856 10548 16908 10600
rect 18604 10548 18656 10600
rect 20444 10548 20496 10600
rect 21180 10616 21232 10668
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 20720 10591 20772 10600
rect 20720 10557 20729 10591
rect 20729 10557 20763 10591
rect 20763 10557 20772 10591
rect 20720 10548 20772 10557
rect 21824 10591 21876 10600
rect 21824 10557 21833 10591
rect 21833 10557 21867 10591
rect 21867 10557 21876 10591
rect 21824 10548 21876 10557
rect 12256 10480 12308 10532
rect 12532 10480 12584 10532
rect 15476 10480 15528 10532
rect 16580 10480 16632 10532
rect 18328 10480 18380 10532
rect 23756 10523 23808 10532
rect 13084 10412 13136 10464
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 19156 10455 19208 10464
rect 19156 10421 19165 10455
rect 19165 10421 19199 10455
rect 19199 10421 19208 10455
rect 19156 10412 19208 10421
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 19984 10412 20036 10464
rect 21180 10412 21232 10464
rect 21640 10455 21692 10464
rect 21640 10421 21649 10455
rect 21649 10421 21683 10455
rect 21683 10421 21692 10455
rect 23756 10489 23765 10523
rect 23765 10489 23799 10523
rect 23799 10489 23808 10523
rect 23756 10480 23808 10489
rect 23388 10455 23440 10464
rect 21640 10412 21692 10421
rect 23388 10421 23397 10455
rect 23397 10421 23431 10455
rect 23431 10421 23440 10455
rect 23388 10412 23440 10421
rect 24768 10412 24820 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 12072 10251 12124 10260
rect 12072 10217 12081 10251
rect 12081 10217 12115 10251
rect 12115 10217 12124 10251
rect 12072 10208 12124 10217
rect 12440 10251 12492 10260
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 14372 10251 14424 10260
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 14740 10208 14792 10260
rect 16856 10251 16908 10260
rect 12808 10183 12860 10192
rect 12808 10149 12817 10183
rect 12817 10149 12851 10183
rect 12851 10149 12860 10183
rect 12808 10140 12860 10149
rect 16856 10217 16865 10251
rect 16865 10217 16899 10251
rect 16899 10217 16908 10251
rect 16856 10208 16908 10217
rect 18420 10208 18472 10260
rect 20444 10208 20496 10260
rect 21824 10208 21876 10260
rect 23112 10208 23164 10260
rect 24860 10208 24912 10260
rect 15292 10115 15344 10124
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 20720 10140 20772 10192
rect 21272 10140 21324 10192
rect 23388 10140 23440 10192
rect 23756 10140 23808 10192
rect 24768 10140 24820 10192
rect 17500 10072 17552 10124
rect 18052 10072 18104 10124
rect 18144 10072 18196 10124
rect 20352 10072 20404 10124
rect 20904 10115 20956 10124
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 23020 10115 23072 10124
rect 23020 10081 23029 10115
rect 23029 10081 23063 10115
rect 23063 10081 23072 10115
rect 23020 10072 23072 10081
rect 24676 10072 24728 10124
rect 26148 10072 26200 10124
rect 13728 9868 13780 9920
rect 15936 10004 15988 10056
rect 19156 10004 19208 10056
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 16580 9936 16632 9988
rect 17868 9936 17920 9988
rect 15476 9868 15528 9920
rect 15752 9911 15804 9920
rect 15752 9877 15761 9911
rect 15761 9877 15795 9911
rect 15795 9877 15804 9911
rect 15752 9868 15804 9877
rect 16672 9868 16724 9920
rect 18236 9911 18288 9920
rect 18236 9877 18245 9911
rect 18245 9877 18279 9911
rect 18279 9877 18288 9911
rect 18236 9868 18288 9877
rect 18604 9911 18656 9920
rect 18604 9877 18613 9911
rect 18613 9877 18647 9911
rect 18647 9877 18656 9911
rect 18604 9868 18656 9877
rect 19248 9868 19300 9920
rect 24952 9868 25004 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 14740 9664 14792 9716
rect 15660 9664 15712 9716
rect 16304 9664 16356 9716
rect 18604 9664 18656 9716
rect 19984 9664 20036 9716
rect 20444 9707 20496 9716
rect 20444 9673 20453 9707
rect 20453 9673 20487 9707
rect 20487 9673 20496 9707
rect 20444 9664 20496 9673
rect 20904 9664 20956 9716
rect 23020 9664 23072 9716
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 25136 9664 25188 9716
rect 26148 9707 26200 9716
rect 26148 9673 26157 9707
rect 26157 9673 26191 9707
rect 26191 9673 26200 9707
rect 26148 9664 26200 9673
rect 9036 9596 9088 9648
rect 13728 9596 13780 9648
rect 14832 9596 14884 9648
rect 15384 9596 15436 9648
rect 16672 9639 16724 9648
rect 16672 9605 16681 9639
rect 16681 9605 16715 9639
rect 16715 9605 16724 9639
rect 16672 9596 16724 9605
rect 18236 9596 18288 9648
rect 19340 9596 19392 9648
rect 12808 9528 12860 9580
rect 15936 9528 15988 9580
rect 16856 9528 16908 9580
rect 13084 9503 13136 9512
rect 13084 9469 13093 9503
rect 13093 9469 13127 9503
rect 13127 9469 13136 9503
rect 13084 9460 13136 9469
rect 14372 9460 14424 9512
rect 16396 9503 16448 9512
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 17500 9460 17552 9512
rect 18788 9528 18840 9580
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 19248 9460 19300 9512
rect 20444 9460 20496 9512
rect 20812 9460 20864 9512
rect 21364 9460 21416 9512
rect 22284 9460 22336 9512
rect 27620 9528 27672 9580
rect 18144 9435 18196 9444
rect 12716 9324 12768 9376
rect 15476 9367 15528 9376
rect 15476 9333 15485 9367
rect 15485 9333 15519 9367
rect 15519 9333 15528 9367
rect 15476 9324 15528 9333
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 18144 9401 18153 9435
rect 18153 9401 18187 9435
rect 18187 9401 18196 9435
rect 18144 9392 18196 9401
rect 19432 9392 19484 9444
rect 17408 9367 17460 9376
rect 15936 9324 15988 9333
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 19156 9367 19208 9376
rect 17408 9324 17460 9333
rect 19156 9333 19165 9367
rect 19165 9333 19199 9367
rect 19199 9333 19208 9367
rect 19156 9324 19208 9333
rect 23940 9367 23992 9376
rect 23940 9333 23949 9367
rect 23949 9333 23983 9367
rect 23983 9333 23992 9367
rect 23940 9324 23992 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 14280 9120 14332 9172
rect 12348 9052 12400 9104
rect 16580 9120 16632 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 18144 9120 18196 9172
rect 19524 9120 19576 9172
rect 20260 9120 20312 9172
rect 21364 9120 21416 9172
rect 14740 9052 14792 9104
rect 15292 9095 15344 9104
rect 15292 9061 15301 9095
rect 15301 9061 15335 9095
rect 15335 9061 15344 9095
rect 15292 9052 15344 9061
rect 22284 9095 22336 9104
rect 22284 9061 22293 9095
rect 22293 9061 22327 9095
rect 22327 9061 22336 9095
rect 22284 9052 22336 9061
rect 24952 9120 25004 9172
rect 23940 9052 23992 9104
rect 24216 9052 24268 9104
rect 11244 8916 11296 8968
rect 12348 8916 12400 8968
rect 13820 8984 13872 9036
rect 15568 8984 15620 9036
rect 18236 8984 18288 9036
rect 15936 8916 15988 8968
rect 17776 8916 17828 8968
rect 22192 8959 22244 8968
rect 22192 8925 22201 8959
rect 22201 8925 22235 8959
rect 22235 8925 22244 8959
rect 22192 8916 22244 8925
rect 24032 8916 24084 8968
rect 17500 8848 17552 8900
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 12532 8780 12584 8832
rect 15384 8780 15436 8832
rect 15844 8780 15896 8832
rect 18604 8780 18656 8832
rect 19248 8823 19300 8832
rect 19248 8789 19257 8823
rect 19257 8789 19291 8823
rect 19291 8789 19300 8823
rect 19248 8780 19300 8789
rect 19340 8780 19392 8832
rect 19708 8823 19760 8832
rect 19708 8789 19717 8823
rect 19717 8789 19751 8823
rect 19751 8789 19760 8823
rect 19708 8780 19760 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 12256 8576 12308 8628
rect 13084 8576 13136 8628
rect 15660 8576 15712 8628
rect 15844 8576 15896 8628
rect 19708 8576 19760 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 22284 8576 22336 8628
rect 23940 8576 23992 8628
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 25412 8576 25464 8628
rect 14372 8508 14424 8560
rect 15936 8508 15988 8560
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12900 8483 12952 8492
rect 12900 8449 12909 8483
rect 12909 8449 12943 8483
rect 12943 8449 12952 8483
rect 12900 8440 12952 8449
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 17408 8508 17460 8560
rect 22652 8508 22704 8560
rect 13820 8440 13872 8449
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 14280 8415 14332 8424
rect 14280 8381 14289 8415
rect 14289 8381 14323 8415
rect 14323 8381 14332 8415
rect 14280 8372 14332 8381
rect 8576 8279 8628 8288
rect 8576 8245 8585 8279
rect 8585 8245 8619 8279
rect 8619 8245 8628 8279
rect 8576 8236 8628 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 14004 8304 14056 8356
rect 15476 8372 15528 8424
rect 16120 8372 16172 8424
rect 18788 8440 18840 8492
rect 21456 8440 21508 8492
rect 22192 8440 22244 8492
rect 24032 8440 24084 8492
rect 24676 8440 24728 8492
rect 14096 8279 14148 8288
rect 12164 8236 12216 8245
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 16856 8279 16908 8288
rect 16856 8245 16865 8279
rect 16865 8245 16899 8279
rect 16899 8245 16908 8279
rect 16856 8236 16908 8245
rect 19248 8372 19300 8424
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 19524 8304 19576 8356
rect 22008 8372 22060 8424
rect 24032 8347 24084 8356
rect 24032 8313 24041 8347
rect 24041 8313 24075 8347
rect 24075 8313 24084 8347
rect 24032 8304 24084 8313
rect 17776 8279 17828 8288
rect 17776 8245 17785 8279
rect 17785 8245 17819 8279
rect 17819 8245 17828 8279
rect 17776 8236 17828 8245
rect 18328 8279 18380 8288
rect 18328 8245 18337 8279
rect 18337 8245 18371 8279
rect 18371 8245 18380 8279
rect 18328 8236 18380 8245
rect 27620 8236 27672 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 14372 8075 14424 8084
rect 14372 8041 14381 8075
rect 14381 8041 14415 8075
rect 14415 8041 14424 8075
rect 14372 8032 14424 8041
rect 14740 8075 14792 8084
rect 14740 8041 14749 8075
rect 14749 8041 14783 8075
rect 14783 8041 14792 8075
rect 14740 8032 14792 8041
rect 15660 8032 15712 8084
rect 16856 8032 16908 8084
rect 17040 8032 17092 8084
rect 21456 8032 21508 8084
rect 24032 8032 24084 8084
rect 8760 8007 8812 8016
rect 8760 7973 8769 8007
rect 8769 7973 8803 8007
rect 8803 7973 8812 8007
rect 8760 7964 8812 7973
rect 12164 7964 12216 8016
rect 20352 7964 20404 8016
rect 22008 7964 22060 8016
rect 24216 8007 24268 8016
rect 24216 7973 24225 8007
rect 24225 7973 24259 8007
rect 24259 7973 24268 8007
rect 24216 7964 24268 7973
rect 24676 7964 24728 8016
rect 8208 7939 8260 7948
rect 8208 7905 8217 7939
rect 8217 7905 8251 7939
rect 8251 7905 8260 7939
rect 8208 7896 8260 7905
rect 8576 7896 8628 7948
rect 10600 7939 10652 7948
rect 10600 7905 10609 7939
rect 10609 7905 10643 7939
rect 10643 7905 10652 7939
rect 10600 7896 10652 7905
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 15292 7896 15344 7905
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 16948 7896 17000 7948
rect 18328 7896 18380 7948
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 19432 7896 19484 7948
rect 21272 7896 21324 7948
rect 22376 7896 22428 7948
rect 11796 7760 11848 7812
rect 14280 7828 14332 7880
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 17224 7828 17276 7880
rect 19156 7828 19208 7880
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 24584 7871 24636 7880
rect 24584 7837 24593 7871
rect 24593 7837 24627 7871
rect 24627 7837 24636 7871
rect 24584 7828 24636 7837
rect 10600 7692 10652 7744
rect 12808 7692 12860 7744
rect 17500 7735 17552 7744
rect 17500 7701 17509 7735
rect 17509 7701 17543 7735
rect 17543 7701 17552 7735
rect 17500 7692 17552 7701
rect 17776 7735 17828 7744
rect 17776 7701 17800 7735
rect 17800 7701 17828 7735
rect 17776 7692 17828 7701
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 24032 7692 24084 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 10600 7531 10652 7540
rect 10600 7497 10609 7531
rect 10609 7497 10643 7531
rect 10643 7497 10652 7531
rect 10600 7488 10652 7497
rect 12072 7488 12124 7540
rect 12440 7488 12492 7540
rect 13636 7488 13688 7540
rect 15292 7488 15344 7540
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 19340 7488 19392 7497
rect 19432 7488 19484 7540
rect 20812 7531 20864 7540
rect 12532 7420 12584 7472
rect 15936 7420 15988 7472
rect 17868 7420 17920 7472
rect 8208 7352 8260 7404
rect 12900 7352 12952 7404
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 24216 7488 24268 7540
rect 25228 7488 25280 7540
rect 1216 7284 1268 7336
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 7748 7216 7800 7268
rect 8576 7148 8628 7200
rect 12808 7259 12860 7268
rect 12808 7225 12817 7259
rect 12817 7225 12851 7259
rect 12851 7225 12860 7259
rect 12808 7216 12860 7225
rect 13084 7216 13136 7268
rect 13728 7216 13780 7268
rect 15752 7284 15804 7336
rect 17500 7284 17552 7336
rect 17960 7284 18012 7336
rect 18788 7284 18840 7336
rect 20812 7284 20864 7336
rect 24676 7352 24728 7404
rect 24032 7327 24084 7336
rect 24032 7293 24041 7327
rect 24041 7293 24075 7327
rect 24075 7293 24084 7327
rect 24032 7284 24084 7293
rect 27620 7284 27672 7336
rect 16212 7259 16264 7268
rect 16212 7225 16221 7259
rect 16221 7225 16255 7259
rect 16255 7225 16264 7259
rect 16212 7216 16264 7225
rect 21732 7259 21784 7268
rect 21732 7225 21741 7259
rect 21741 7225 21775 7259
rect 21775 7225 21784 7259
rect 21732 7216 21784 7225
rect 13268 7148 13320 7200
rect 14188 7148 14240 7200
rect 15476 7148 15528 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 18328 7191 18380 7200
rect 18328 7157 18337 7191
rect 18337 7157 18371 7191
rect 18371 7157 18380 7191
rect 18328 7148 18380 7157
rect 22008 7191 22060 7200
rect 22008 7157 22017 7191
rect 22017 7157 22051 7191
rect 22051 7157 22060 7191
rect 22008 7148 22060 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 12164 6987 12216 6996
rect 12164 6953 12173 6987
rect 12173 6953 12207 6987
rect 12207 6953 12216 6987
rect 12164 6944 12216 6953
rect 12808 6944 12860 6996
rect 15752 6944 15804 6996
rect 18788 6987 18840 6996
rect 18788 6953 18797 6987
rect 18797 6953 18831 6987
rect 18831 6953 18840 6987
rect 18788 6944 18840 6953
rect 24032 6944 24084 6996
rect 15936 6876 15988 6928
rect 22008 6876 22060 6928
rect 11796 6808 11848 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14004 6808 14056 6860
rect 16028 6808 16080 6860
rect 16212 6808 16264 6860
rect 19432 6808 19484 6860
rect 21732 6808 21784 6860
rect 23020 6808 23072 6860
rect 24216 6851 24268 6860
rect 24216 6817 24225 6851
rect 24225 6817 24259 6851
rect 24259 6817 24268 6851
rect 24216 6808 24268 6817
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 24124 6783 24176 6792
rect 24124 6749 24133 6783
rect 24133 6749 24167 6783
rect 24167 6749 24176 6783
rect 24124 6740 24176 6749
rect 2136 6604 2188 6656
rect 8668 6604 8720 6656
rect 16580 6604 16632 6656
rect 17776 6604 17828 6656
rect 19064 6604 19116 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 12348 6400 12400 6452
rect 14004 6400 14056 6452
rect 16028 6400 16080 6452
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 22008 6400 22060 6452
rect 22560 6400 22612 6452
rect 23020 6443 23072 6452
rect 23020 6409 23029 6443
rect 23029 6409 23063 6443
rect 23063 6409 23072 6443
rect 23020 6400 23072 6409
rect 24124 6400 24176 6452
rect 11796 6332 11848 6384
rect 13728 6332 13780 6384
rect 16304 6332 16356 6384
rect 18512 6332 18564 6384
rect 24216 6332 24268 6384
rect 14188 6264 14240 6316
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 24584 6264 24636 6316
rect 13636 6128 13688 6180
rect 15936 6128 15988 6180
rect 15384 6060 15436 6112
rect 16580 6171 16632 6180
rect 16580 6137 16589 6171
rect 16589 6137 16623 6171
rect 16623 6137 16632 6171
rect 17132 6171 17184 6180
rect 16580 6128 16632 6137
rect 17132 6137 17141 6171
rect 17141 6137 17175 6171
rect 17175 6137 17184 6171
rect 17132 6128 17184 6137
rect 18328 6128 18380 6180
rect 24124 6060 24176 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 14188 5856 14240 5908
rect 16488 5856 16540 5908
rect 24216 5856 24268 5908
rect 14464 5720 14516 5772
rect 17132 5788 17184 5840
rect 17868 5831 17920 5840
rect 17868 5797 17877 5831
rect 17877 5797 17911 5831
rect 17911 5797 17920 5831
rect 17868 5788 17920 5797
rect 17960 5831 18012 5840
rect 17960 5797 17969 5831
rect 17969 5797 18003 5831
rect 18003 5797 18012 5831
rect 18512 5831 18564 5840
rect 17960 5788 18012 5797
rect 18512 5797 18521 5831
rect 18521 5797 18555 5831
rect 18555 5797 18564 5831
rect 18512 5788 18564 5797
rect 22008 5788 22060 5840
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 19984 5720 20036 5772
rect 22560 5720 22612 5772
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 23480 5652 23532 5704
rect 24584 5695 24636 5704
rect 16580 5584 16632 5636
rect 17408 5584 17460 5636
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24676 5584 24728 5636
rect 24032 5516 24084 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 12716 5312 12768 5364
rect 15292 5312 15344 5364
rect 17960 5312 18012 5364
rect 22008 5312 22060 5364
rect 13728 5244 13780 5296
rect 14096 5176 14148 5228
rect 14464 5176 14516 5228
rect 17868 5176 17920 5228
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 13912 5108 13964 5160
rect 13636 5083 13688 5092
rect 13636 5049 13645 5083
rect 13645 5049 13679 5083
rect 13679 5049 13688 5083
rect 13636 5040 13688 5049
rect 14372 5040 14424 5092
rect 15660 5083 15712 5092
rect 15660 5049 15669 5083
rect 15669 5049 15703 5083
rect 15703 5049 15712 5083
rect 15660 5040 15712 5049
rect 18144 5083 18196 5092
rect 15384 4972 15436 5024
rect 18144 5049 18153 5083
rect 18153 5049 18187 5083
rect 18187 5049 18196 5083
rect 18144 5040 18196 5049
rect 22560 5312 22612 5364
rect 23480 5355 23532 5364
rect 23480 5321 23489 5355
rect 23489 5321 23523 5355
rect 23523 5321 23532 5355
rect 23480 5312 23532 5321
rect 24216 5312 24268 5364
rect 26056 5355 26108 5364
rect 26056 5321 26065 5355
rect 26065 5321 26099 5355
rect 26099 5321 26108 5355
rect 26056 5312 26108 5321
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 26056 5108 26108 5160
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 25964 5040 26016 5092
rect 24400 5015 24452 5024
rect 17776 4972 17828 4981
rect 24400 4981 24409 5015
rect 24409 4981 24443 5015
rect 24443 4981 24452 5015
rect 24400 4972 24452 4981
rect 25044 4972 25096 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 14096 4768 14148 4820
rect 15660 4768 15712 4820
rect 17776 4811 17828 4820
rect 17776 4777 17785 4811
rect 17785 4777 17819 4811
rect 17819 4777 17828 4811
rect 17776 4768 17828 4777
rect 18144 4768 18196 4820
rect 24032 4811 24084 4820
rect 24032 4777 24041 4811
rect 24041 4777 24075 4811
rect 24075 4777 24084 4811
rect 24032 4768 24084 4777
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 13820 4700 13872 4709
rect 1584 4632 1636 4684
rect 24124 4700 24176 4752
rect 24400 4700 24452 4752
rect 24676 4700 24728 4752
rect 15844 4632 15896 4684
rect 17408 4675 17460 4684
rect 17408 4641 17417 4675
rect 17417 4641 17451 4675
rect 17451 4641 17460 4675
rect 17408 4632 17460 4641
rect 18972 4632 19024 4684
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 15292 4607 15344 4616
rect 15292 4573 15301 4607
rect 15301 4573 15335 4607
rect 15335 4573 15344 4607
rect 15292 4564 15344 4573
rect 25228 4564 25280 4616
rect 10508 4496 10560 4548
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 10508 4224 10560 4276
rect 13728 4224 13780 4276
rect 15844 4267 15896 4276
rect 15844 4233 15853 4267
rect 15853 4233 15887 4267
rect 15887 4233 15896 4267
rect 15844 4224 15896 4233
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 18972 4267 19024 4276
rect 18972 4233 18981 4267
rect 18981 4233 19015 4267
rect 19015 4233 19024 4267
rect 18972 4224 19024 4233
rect 24124 4267 24176 4276
rect 24124 4233 24133 4267
rect 24133 4233 24167 4267
rect 24167 4233 24176 4267
rect 24124 4224 24176 4233
rect 25228 4267 25280 4276
rect 25228 4233 25237 4267
rect 25237 4233 25271 4267
rect 25271 4233 25280 4267
rect 25228 4224 25280 4233
rect 13820 4088 13872 4140
rect 14372 4088 14424 4140
rect 24676 4131 24728 4140
rect 24676 4097 24685 4131
rect 24685 4097 24719 4131
rect 24719 4097 24728 4131
rect 24676 4088 24728 4097
rect 12992 4020 13044 4072
rect 14924 3995 14976 4004
rect 14924 3961 14933 3995
rect 14933 3961 14967 3995
rect 14967 3961 14976 3995
rect 14924 3952 14976 3961
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 15292 3952 15344 4004
rect 24308 3995 24360 4004
rect 24308 3961 24317 3995
rect 24317 3961 24351 3995
rect 24351 3961 24360 3995
rect 24308 3952 24360 3961
rect 24032 3884 24084 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 12992 3723 13044 3732
rect 12992 3689 13001 3723
rect 13001 3689 13035 3723
rect 13035 3689 13044 3723
rect 12992 3680 13044 3689
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 24032 3680 24084 3732
rect 24308 3680 24360 3732
rect 12256 3612 12308 3664
rect 13636 3612 13688 3664
rect 12164 3544 12216 3596
rect 15384 3544 15436 3596
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 24676 3340 24728 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 12164 3136 12216 3188
rect 15384 3179 15436 3188
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 12256 3000 12308 3052
rect 13360 3068 13412 3120
rect 13268 3043 13320 3052
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 12900 2907 12952 2916
rect 12900 2873 12909 2907
rect 12909 2873 12943 2907
rect 12943 2873 12952 2907
rect 12900 2864 12952 2873
rect 24676 2839 24728 2848
rect 24676 2805 24685 2839
rect 24685 2805 24719 2839
rect 24719 2805 24728 2839
rect 24676 2796 24728 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 12992 2592 13044 2644
rect 13360 2592 13412 2644
rect 25228 2592 25280 2644
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 25136 2456 25188 2508
rect 14740 2431 14792 2440
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 25136 2295 25188 2304
rect 25136 2261 25145 2295
rect 25145 2261 25179 2295
rect 25179 2261 25188 2295
rect 25136 2252 25188 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 5264 76 5316 128
rect 11980 76 12032 128
<< metal2 >>
rect 754 27520 810 28000
rect 2226 27554 2282 28000
rect 2226 27526 2452 27554
rect 2226 27520 2282 27526
rect 768 24274 796 27520
rect 1306 25664 1362 25673
rect 1306 25599 1362 25608
rect 756 24268 808 24274
rect 756 24210 808 24216
rect 1320 23730 1348 25599
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 1872 23866 1900 24210
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1308 23724 1360 23730
rect 1308 23666 1360 23672
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1122 22128 1178 22137
rect 1122 22063 1178 22072
rect 1136 21010 1164 22063
rect 1124 21004 1176 21010
rect 1124 20946 1176 20952
rect 1136 20602 1164 20946
rect 1124 20596 1176 20602
rect 1124 20538 1176 20544
rect 1122 18592 1178 18601
rect 1122 18527 1178 18536
rect 1136 17746 1164 18527
rect 1124 17740 1176 17746
rect 1124 17682 1176 17688
rect 1136 17338 1164 17682
rect 1124 17332 1176 17338
rect 1124 17274 1176 17280
rect 1780 15065 1808 23462
rect 2424 17338 2452 27526
rect 3790 27520 3846 28000
rect 5354 27554 5410 28000
rect 5354 27526 5580 27554
rect 5354 27520 5410 27526
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2424 17134 2452 17274
rect 2412 17128 2464 17134
rect 1950 17096 2006 17105
rect 2412 17070 2464 17076
rect 1950 17031 2006 17040
rect 1964 16998 1992 17031
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1766 15056 1822 15065
rect 1766 14991 1822 15000
rect 2700 11665 2728 24006
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3252 16017 3280 20742
rect 3804 18426 3832 27520
rect 5552 20602 5580 27526
rect 6918 27520 6974 28000
rect 8482 27520 8538 28000
rect 10046 27520 10102 28000
rect 11610 27554 11666 28000
rect 11610 27526 11744 27554
rect 11610 27520 11666 27526
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6932 24313 6960 27520
rect 8496 24721 8524 27520
rect 8482 24712 8538 24721
rect 8482 24647 8538 24656
rect 6918 24304 6974 24313
rect 6918 24239 6974 24248
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 10060 21010 10088 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 11716 23866 11744 27526
rect 13174 27520 13230 28000
rect 14738 27520 14794 28000
rect 16210 27554 16266 28000
rect 17774 27554 17830 28000
rect 15948 27526 16266 27554
rect 13188 24274 13216 27520
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13188 23866 13216 24210
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 11716 23662 11744 23802
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12820 22438 12848 22918
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 11796 21004 11848 21010
rect 11796 20946 11848 20952
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 11808 20602 11836 20946
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 5552 20398 5580 20538
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 9692 19281 9720 20198
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 9678 19272 9734 19281
rect 9678 19207 9734 19216
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3804 18222 3832 18362
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17241 3924 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 3882 17232 3938 17241
rect 3882 17167 3938 17176
rect 8956 16561 8984 17478
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 12256 16584 12308 16590
rect 8942 16552 8998 16561
rect 12256 16526 12308 16532
rect 8942 16487 8998 16496
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 12268 16250 12296 16526
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 12636 15706 12664 19178
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5446 15192 5502 15201
rect 5622 15184 5918 15204
rect 5446 15127 5502 15136
rect 12164 15156 12216 15162
rect 5460 14958 5488 15127
rect 12164 15098 12216 15104
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 11532 14482 11560 14962
rect 11520 14476 11572 14482
rect 11520 14418 11572 14424
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 11532 14074 11560 14418
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 14074 11836 14350
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 12176 13734 12204 15098
rect 12268 14618 12296 15438
rect 12636 15162 12664 15642
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12636 14890 12664 14962
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12268 14260 12296 14554
rect 12268 14232 12388 14260
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 11808 12306 11836 12922
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 12306 11928 12582
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 11808 11898 11836 12242
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 1306 11656 1362 11665
rect 1306 11591 1362 11600
rect 2686 11656 2742 11665
rect 2686 11591 2742 11600
rect 1320 11218 1348 11591
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 1308 11212 1360 11218
rect 1308 11154 1360 11160
rect 1320 10810 1348 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 1308 10804 1360 10810
rect 1308 10746 1360 10752
rect 11808 10742 11836 11834
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10888 10266 10916 10542
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 8680 8430 8708 8774
rect 9048 8498 9076 9590
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11256 8634 11284 8910
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8758 8392 8814 8401
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 1214 8120 1270 8129
rect 1214 8055 1270 8064
rect 1228 7342 1256 8055
rect 8588 7954 8616 8230
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 8220 7410 8248 7890
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 1216 7336 1268 7342
rect 1216 7278 1268 7284
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7760 6905 7788 7210
rect 8588 7206 8616 7890
rect 8680 7342 8708 8366
rect 8758 8327 8814 8336
rect 8772 8022 8800 8327
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10612 7750 10640 7890
rect 11808 7818 11836 10678
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10612 7546 10640 7686
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 7746 6896 7802 6905
rect 7746 6831 7802 6840
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1596 4593 1624 4626
rect 1582 4584 1638 4593
rect 1582 4519 1638 4528
rect 1596 4282 1624 4519
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1872 2281 1900 2450
rect 1858 2272 1914 2281
rect 1858 2207 1914 2216
rect 1766 82 1822 480
rect 2148 82 2176 6598
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 1766 54 2176 82
rect 5262 128 5318 480
rect 5262 76 5264 128
rect 5316 76 5318 128
rect 1766 0 1822 54
rect 5262 0 5318 76
rect 8588 82 8616 7142
rect 8680 6662 8708 7278
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 11808 6866 11836 7754
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 11808 6390 11836 6802
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10520 4282 10548 4490
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 8758 82 8814 480
rect 11992 134 12020 12718
rect 12176 11558 12204 13670
rect 12268 13394 12296 13874
rect 12360 13530 12388 14232
rect 12636 14074 12664 14826
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 12918 12296 13330
rect 12544 13190 12572 13806
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12256 12912 12308 12918
rect 12308 12872 12388 12900
rect 12256 12854 12308 12860
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12360 11286 12388 12872
rect 12544 12374 12572 13126
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12636 12306 12664 13330
rect 12820 12918 12848 22374
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20466 12940 20742
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 19242 12940 20198
rect 13004 19922 13032 20266
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13004 19310 13032 19654
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 13004 18154 13032 19246
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12912 16130 12940 17070
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13004 16726 13032 16934
rect 12992 16720 13044 16726
rect 12992 16662 13044 16668
rect 13004 16250 13032 16662
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12912 16102 13032 16130
rect 13004 15978 13032 16102
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 12912 15706 12940 15914
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12912 15026 12940 15642
rect 13004 15570 13032 15914
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 14414 12940 14962
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 13096 13814 13124 22510
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13188 19174 13216 19858
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13188 18970 13216 19110
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 12912 13786 13124 13814
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11694 12848 12038
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 12084 10266 12112 11086
rect 12268 10538 12296 11222
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12084 7954 12112 9114
rect 12360 9110 12388 11222
rect 12544 10742 12572 11494
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10266 12480 10542
rect 12544 10538 12572 10678
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 10146 12572 10474
rect 12452 10118 12572 10146
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12348 9104 12400 9110
rect 12268 9052 12348 9058
rect 12268 9046 12400 9052
rect 12268 9030 12388 9046
rect 12268 8634 12296 9030
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 8022 12204 8230
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7546 12112 7890
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12176 3602 12204 6938
rect 12360 6866 12388 8910
rect 12452 8090 12480 10118
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9382 12756 9998
rect 12820 9586 12848 10134
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8498 12572 8774
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12452 7546 12480 8026
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12360 6458 12388 6802
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12176 3194 12204 3538
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12268 3058 12296 3606
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 8588 54 8814 82
rect 11980 128 12032 134
rect 11980 70 12032 76
rect 12254 82 12310 480
rect 12544 82 12572 7414
rect 12728 5370 12756 9318
rect 12912 8498 12940 13786
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11150 13032 12038
rect 13096 11626 13124 12242
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11354 13124 11562
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 10062 13032 11086
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13096 9518 13124 10406
rect 13280 9625 13308 24006
rect 14752 23866 14780 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23866 15332 24210
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 13556 22778 13584 23598
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 13636 23180 13688 23186
rect 13636 23122 13688 23128
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13648 22234 13676 23122
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22642 14596 22918
rect 14752 22642 14780 23462
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13648 19802 13676 22170
rect 14292 21554 14320 22374
rect 14568 22234 14596 22578
rect 15304 22234 15332 23598
rect 15580 23322 15608 23802
rect 15948 23798 15976 27526
rect 16210 27520 16266 27526
rect 17512 27526 17830 27554
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 16960 23730 16988 24550
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17420 23866 17448 24210
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15764 23254 15792 23598
rect 16684 23322 16712 23598
rect 17420 23474 17448 23802
rect 17512 23798 17540 27526
rect 17774 27520 17830 27526
rect 19338 27520 19394 28000
rect 20902 27554 20958 28000
rect 20640 27526 20958 27554
rect 18880 24880 18932 24886
rect 18880 24822 18932 24828
rect 18602 24712 18658 24721
rect 18602 24647 18658 24656
rect 18788 24676 18840 24682
rect 18616 24274 18644 24647
rect 18788 24618 18840 24624
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 17776 23520 17828 23526
rect 17420 23446 17540 23474
rect 17776 23462 17828 23468
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 15752 23248 15804 23254
rect 15752 23190 15804 23196
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 16132 22710 16160 23122
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 14556 22228 14608 22234
rect 14556 22170 14608 22176
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14384 21078 14412 21354
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13740 20330 13768 20742
rect 13832 20602 13860 21014
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13556 19774 13676 19802
rect 13556 16726 13584 19774
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 18902 13676 19654
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13648 18426 13676 18838
rect 13740 18766 13768 20266
rect 14384 20058 14412 20334
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 14016 18086 14044 18566
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14016 17882 14044 18022
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13556 16114 13584 16662
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14200 14822 14228 15506
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 14482 14228 14758
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 13544 14340 13596 14346
rect 13544 14282 13596 14288
rect 13556 13734 13584 14282
rect 14200 14074 14228 14418
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14384 13870 14412 14214
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13358 12880 13414 12889
rect 13464 12850 13492 13126
rect 13358 12815 13414 12824
rect 13452 12844 13504 12850
rect 13372 12782 13400 12815
rect 13452 12786 13504 12792
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13372 11762 13400 12582
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13464 11830 13492 12310
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13464 11354 13492 11766
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13266 9616 13322 9625
rect 13266 9551 13322 9560
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12900 8492 12952 8498
rect 12900 8434 12952 8440
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7274 12848 7686
rect 12912 7410 12940 8434
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13096 7274 13124 8570
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12820 7002 12848 7210
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 2922 12940 3878
rect 13004 3738 13032 4014
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 13004 2650 13032 3674
rect 13280 3058 13308 7142
rect 13358 5264 13414 5273
rect 13358 5199 13414 5208
rect 13372 5166 13400 5199
rect 13360 5160 13412 5166
rect 13556 5137 13584 13670
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 12986 13952 13330
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 12238 13952 12786
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13648 11354 13676 11630
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13648 10810 13676 11154
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13740 10674 13768 11086
rect 14108 10810 14136 11154
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10266 13768 10610
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14384 10266 14412 10542
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9654 13768 9862
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 14384 9518 14412 10202
rect 14372 9512 14424 9518
rect 14292 9472 14372 9500
rect 14292 9178 14320 9472
rect 14372 9454 14424 9460
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8498 13860 8978
rect 14372 8560 14424 8566
rect 14372 8502 14424 8508
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13832 8401 13860 8434
rect 14280 8424 14332 8430
rect 13818 8392 13874 8401
rect 14280 8366 14332 8372
rect 13818 8327 13874 8336
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13648 6186 13676 7482
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 6866 13768 7210
rect 14016 6866 14044 8298
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13740 6390 13768 6802
rect 14016 6458 14044 6802
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13360 5102 13412 5108
rect 13542 5128 13598 5137
rect 13648 5098 13676 6122
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5302 13768 5646
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 14108 5234 14136 8230
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7206 14228 7890
rect 14292 7886 14320 8366
rect 14384 8090 14412 8502
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14200 6322 14228 6734
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14200 5914 14228 6258
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14476 5778 14504 21286
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20602 15332 21422
rect 15396 21418 15424 22442
rect 16132 22114 16160 22646
rect 16212 22636 16264 22642
rect 16212 22578 16264 22584
rect 16224 22234 16252 22578
rect 16396 22500 16448 22506
rect 16396 22442 16448 22448
rect 16212 22228 16264 22234
rect 16212 22170 16264 22176
rect 15476 22092 15528 22098
rect 16132 22086 16252 22114
rect 16408 22098 16436 22442
rect 17144 22438 17172 23122
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 15476 22034 15528 22040
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15488 21350 15516 22034
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 16132 20534 16160 21082
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19242 15332 19858
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 14844 18222 14872 19178
rect 15580 18834 15608 19246
rect 15856 19174 15884 19858
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19310 15976 19790
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15580 18630 15608 18770
rect 15856 18698 15884 19110
rect 15948 18970 15976 19246
rect 16132 18970 16160 20334
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14844 18086 14872 18158
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14740 16584 14792 16590
rect 14738 16552 14740 16561
rect 14792 16552 14794 16561
rect 14738 16487 14794 16496
rect 14752 16250 14780 16487
rect 14740 16244 14792 16250
rect 14740 16186 14792 16192
rect 14844 16130 14872 18022
rect 15212 17814 15240 18090
rect 15580 18086 15608 18566
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15384 17128 15436 17134
rect 15384 17070 15436 17076
rect 15396 16726 15424 17070
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15384 16720 15436 16726
rect 15384 16662 15436 16668
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14752 16102 14872 16130
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14660 14278 14688 14894
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 13462 14688 14214
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14752 12782 14780 16102
rect 15396 15910 15424 16662
rect 15488 16250 15516 17002
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15488 15910 15516 16186
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 14890 15332 15438
rect 15396 15162 15424 15846
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13938 15332 14826
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14844 13394 14872 13806
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14844 13190 14872 13330
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14752 12442 14780 12718
rect 14844 12628 14872 13126
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15016 12640 15068 12646
rect 14844 12600 15016 12628
rect 15016 12582 15068 12588
rect 15028 12442 15056 12582
rect 14740 12436 14792 12442
rect 14660 12396 14740 12424
rect 14660 11626 14688 12396
rect 14740 12378 14792 12384
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15580 12374 15608 18022
rect 15856 17542 15884 18634
rect 15948 18290 15976 18906
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15856 16454 15884 17478
rect 16132 17338 16160 17682
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 16132 16726 16160 17274
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15856 15706 15884 16390
rect 16040 16114 16068 16526
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16040 15706 16068 16050
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 15948 15162 15976 15574
rect 16132 15570 16160 16662
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15948 14958 15976 15098
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14482 15700 14758
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 13734 15700 14418
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13394 15700 13670
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12986 15700 13330
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15672 12889 15700 12922
rect 16132 12918 16160 13126
rect 16120 12912 16172 12918
rect 15658 12880 15714 12889
rect 16120 12854 16172 12860
rect 15658 12815 15714 12824
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11880 14780 12038
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14813 11892 14865 11898
rect 14752 11852 14813 11880
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14660 10266 14688 11562
rect 14752 11354 14780 11852
rect 14813 11834 14865 11840
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15396 11558 15424 11766
rect 15580 11626 15608 12310
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11620 15620 11626
rect 15568 11562 15620 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14752 10742 14780 11290
rect 15396 11014 15424 11494
rect 15580 11286 15608 11562
rect 15672 11558 15700 12038
rect 16132 11558 16160 12854
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14752 10266 14780 10678
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 10470 14872 10610
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14752 9722 14780 10202
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14844 9654 14872 10406
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 15304 9110 15332 10066
rect 15396 9654 15424 10950
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15488 10538 15516 10610
rect 15580 10606 15608 11222
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15488 9926 15516 10474
rect 16040 10470 16068 11154
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 14752 8090 14780 9046
rect 15396 8838 15424 9590
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15488 8430 15516 9318
rect 15568 9036 15620 9042
rect 15672 9024 15700 9658
rect 15620 8996 15700 9024
rect 15568 8978 15620 8984
rect 15672 8634 15700 8996
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15672 8090 15700 8570
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15764 7954 15792 9862
rect 15948 9586 15976 9998
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9382 15976 9522
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 8974 15976 9318
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 8634 15884 8774
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15948 8566 15976 8910
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 16040 8412 16068 10406
rect 16132 8430 16160 11494
rect 15948 8384 16068 8412
rect 16120 8424 16172 8430
rect 15292 7948 15344 7954
rect 15292 7890 15344 7896
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7546 15332 7890
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15764 7342 15792 7890
rect 15948 7478 15976 8384
rect 16120 8366 16172 8372
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15396 5778 15424 6054
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 14476 5234 14504 5714
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5370 15332 5646
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 13912 5160 13964 5166
rect 13832 5120 13912 5148
rect 13542 5063 13598 5072
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 3670 13676 5034
rect 13832 4758 13860 5120
rect 13912 5102 13964 5108
rect 14108 4826 14136 5170
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 4282 13768 4558
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13832 4146 13860 4694
rect 14384 4622 14412 5034
rect 15396 5030 15424 5714
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 15292 4616 15344 4622
rect 15292 4558 15344 4564
rect 14384 4146 14412 4558
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 15304 4010 15332 4558
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 14936 3738 14964 3946
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 13636 3664 13688 3670
rect 13636 3606 13688 3612
rect 15382 3632 15438 3641
rect 15382 3567 15384 3576
rect 15436 3567 15438 3576
rect 15384 3538 15436 3544
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 3126 13400 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15396 3194 15424 3538
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13280 2378 13308 2994
rect 13372 2650 13400 3062
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 14738 2544 14794 2553
rect 14738 2479 14794 2488
rect 14752 2446 14780 2479
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 8758 0 8814 54
rect 12254 54 12572 82
rect 15488 82 15516 7142
rect 15764 7002 15792 7278
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 15948 6186 15976 6870
rect 16040 6866 16068 7822
rect 16224 7426 16252 22086
rect 16396 22092 16448 22098
rect 16396 22034 16448 22040
rect 16408 21350 16436 22034
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 21146 16436 21286
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16500 20262 16528 20470
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16592 19718 16620 20878
rect 17144 20602 17172 22374
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19514 16620 19654
rect 16580 19508 16632 19514
rect 16580 19450 16632 19456
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16316 17338 16344 17478
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16316 16998 16344 17274
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16408 16794 16436 17138
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16500 16674 16528 17478
rect 16316 16646 16528 16674
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16316 9722 16344 16646
rect 16960 16250 16988 16662
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 14958 16620 15302
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16592 14618 16620 14894
rect 16960 14822 16988 15506
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16396 14340 16448 14346
rect 16396 14282 16448 14288
rect 16408 13870 16436 14282
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13870 16528 14214
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16408 13258 16436 13806
rect 16868 13394 16896 13806
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16500 12918 16528 13126
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16500 12374 16528 12854
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16592 12646 16620 12786
rect 16684 12714 16712 13330
rect 16868 12986 16896 13330
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16500 11898 16528 12310
rect 16592 12238 16620 12582
rect 16684 12442 16712 12650
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16500 10742 16528 11834
rect 16592 11762 16620 12174
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16592 11014 16620 11698
rect 16684 11150 16712 12242
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16868 11898 16896 12106
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 9994 16620 10474
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16396 9512 16448 9518
rect 16592 9500 16620 9930
rect 16684 9926 16712 11086
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16868 10266 16896 10542
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16672 9920 16724 9926
rect 16672 9862 16724 9868
rect 16684 9654 16712 9862
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16868 9586 16896 10202
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16448 9472 16620 9500
rect 16396 9454 16448 9460
rect 16592 9178 16620 9472
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16868 8090 16896 8230
rect 17052 8090 17080 18158
rect 17420 16402 17448 20742
rect 17512 17270 17540 23446
rect 17788 23254 17816 23462
rect 18156 23322 18184 23666
rect 18800 23594 18828 24618
rect 18788 23588 18840 23594
rect 18788 23530 18840 23536
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18156 22506 18184 22918
rect 18800 22642 18828 23530
rect 18892 23225 18920 24822
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 19168 23866 19196 24210
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19156 23860 19208 23866
rect 19156 23802 19208 23808
rect 19260 23474 19288 24006
rect 19352 23798 19380 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19444 24313 19472 24686
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19430 24304 19486 24313
rect 19430 24239 19486 24248
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19260 23446 19564 23474
rect 18878 23216 18934 23225
rect 18878 23151 18934 23160
rect 19260 23118 19288 23446
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19444 22778 19472 23190
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 18156 22030 18184 22442
rect 19444 22438 19472 22714
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 18236 22160 18288 22166
rect 18236 22102 18288 22108
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17972 21554 18000 21966
rect 18248 21690 18276 22102
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 19168 21486 19196 21830
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17788 19310 17816 19858
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17880 19242 17908 20198
rect 18064 19990 18092 21422
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 21078 19380 21286
rect 19444 21146 19472 22374
rect 19536 22234 19564 23446
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 19904 22506 19932 23190
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19996 22506 20024 22578
rect 19892 22500 19944 22506
rect 19892 22442 19944 22448
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 20088 21690 20116 22374
rect 20364 22030 20392 24618
rect 20640 24342 20668 27526
rect 20902 27520 20958 27526
rect 22466 27520 22522 28000
rect 24030 27554 24086 28000
rect 23676 27526 24086 27554
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 20628 24336 20680 24342
rect 20628 24278 20680 24284
rect 21008 24206 21036 24550
rect 22480 24410 22508 27520
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20456 23594 20484 24006
rect 20444 23588 20496 23594
rect 20444 23530 20496 23536
rect 20456 23050 20484 23530
rect 20548 23322 20576 24006
rect 21008 23798 21036 24142
rect 21100 23866 21128 24278
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 21272 24200 21324 24206
rect 21272 24142 21324 24148
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 21284 23730 21312 24142
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20536 23316 20588 23322
rect 20536 23258 20588 23264
rect 21008 23186 21036 23462
rect 21376 23322 21404 23802
rect 22480 23730 22508 24210
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22008 23656 22060 23662
rect 22008 23598 22060 23604
rect 22020 23322 22048 23598
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 20444 23044 20496 23050
rect 20444 22986 20496 22992
rect 20456 22710 20484 22986
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20536 22500 20588 22506
rect 20456 22460 20536 22488
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 19708 21616 19760 21622
rect 19708 21558 19760 21564
rect 19720 21457 19748 21558
rect 19706 21448 19762 21457
rect 19706 21383 19762 21392
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 20364 21146 20392 21966
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 18616 19718 18644 20878
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20398 18736 20742
rect 19352 20534 19380 21014
rect 19800 20800 19852 20806
rect 19800 20742 19852 20748
rect 19340 20528 19392 20534
rect 19340 20470 19392 20476
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18708 19990 18736 20334
rect 19352 20262 19380 20470
rect 19812 20466 19840 20742
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 18696 19984 18748 19990
rect 18696 19926 18748 19932
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 17868 19236 17920 19242
rect 17868 19178 17920 19184
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18064 18222 18092 19110
rect 18524 18222 18552 19246
rect 18616 18290 18644 19654
rect 19168 19310 19196 19654
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18708 18834 18736 19110
rect 19168 18834 19196 19246
rect 19352 19242 19380 20198
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20088 19514 20116 19858
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 18708 18426 18736 18770
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 17512 16522 17540 17206
rect 17604 17202 17632 17614
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17500 16516 17552 16522
rect 17500 16458 17552 16464
rect 17420 16374 17540 16402
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 13938 17172 14350
rect 17420 14074 17448 14418
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17512 12442 17540 16374
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10742 17172 10950
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9518 17540 10066
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17420 8566 17448 9318
rect 17512 9178 17540 9454
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17512 8906 17540 9114
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17696 7993 17724 15846
rect 17788 15434 17816 18022
rect 18524 17542 18552 18158
rect 19168 18154 19196 18770
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18340 16046 18368 16390
rect 18328 16040 18380 16046
rect 17866 16008 17922 16017
rect 18328 15982 18380 15988
rect 17866 15943 17922 15952
rect 17880 15706 17908 15943
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17880 14958 17908 15642
rect 18524 15570 18552 15846
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18340 15434 18368 15506
rect 18328 15428 18380 15434
rect 18328 15370 18380 15376
rect 18340 15162 18368 15370
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 18156 14550 18184 15098
rect 18328 14884 18380 14890
rect 18248 14844 18328 14872
rect 18248 14618 18276 14844
rect 18328 14826 18380 14832
rect 18524 14822 18552 15506
rect 18616 15502 18644 16526
rect 18604 15496 18656 15502
rect 18604 15438 18656 15444
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18156 14074 18184 14486
rect 18248 14074 18276 14554
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13462 18092 13806
rect 18156 13802 18184 14010
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18156 13530 18184 13738
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17972 12646 18000 12718
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17788 11558 17816 11766
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17788 10810 17816 11494
rect 17880 11014 17908 11630
rect 17972 11150 18000 12582
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17880 10742 17908 10950
rect 17868 10736 17920 10742
rect 17868 10678 17920 10684
rect 17880 9994 17908 10678
rect 18064 10130 18092 12038
rect 18156 11558 18184 12242
rect 18524 11898 18552 14758
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12238 18644 12582
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18616 11830 18644 12174
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18156 11014 18184 11494
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10130 18184 10950
rect 18340 10538 18368 11154
rect 18432 10674 18460 11698
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18432 10266 18460 10610
rect 18616 10606 18644 11766
rect 18708 11014 18736 12310
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 18156 9450 18184 10066
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18604 9920 18656 9926
rect 18708 9908 18736 10950
rect 18800 10810 18828 18090
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 18892 16998 18920 17682
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19444 17134 19472 17478
rect 19996 17270 20024 17682
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18892 16697 18920 16934
rect 18878 16688 18934 16697
rect 18878 16623 18934 16632
rect 19076 16114 19104 17070
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19352 16726 19380 17002
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16794 20024 17206
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19352 16250 19380 16662
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 13462 18920 14962
rect 19064 14884 19116 14890
rect 19064 14826 19116 14832
rect 19076 13802 19104 14826
rect 19352 14550 19380 16186
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19996 15026 20024 15302
rect 20456 15026 20484 22460
rect 20536 22442 20588 22448
rect 21008 22438 21036 23122
rect 22480 22506 22508 23122
rect 22468 22500 22520 22506
rect 22468 22442 22520 22448
rect 23124 22438 23152 23122
rect 23216 22642 23244 24550
rect 23676 23866 23704 27526
rect 24030 27520 24086 27526
rect 25594 27520 25650 28000
rect 27158 27520 27214 28000
rect 24950 26888 25006 26897
rect 24950 26823 25006 26832
rect 24766 25936 24822 25945
rect 24766 25871 24822 25880
rect 24676 25356 24728 25362
rect 24676 25298 24728 25304
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24216 24744 24268 24750
rect 24216 24686 24268 24692
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23768 23474 23796 24550
rect 23848 24268 23900 24274
rect 23848 24210 23900 24216
rect 23860 23866 23888 24210
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23676 23446 23796 23474
rect 23860 23474 23888 23802
rect 23860 23446 24072 23474
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20824 21350 20852 22034
rect 21100 21690 21128 22102
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20628 19304 20680 19310
rect 20628 19246 20680 19252
rect 20640 18970 20668 19246
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20732 17338 20760 17750
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 16522 20576 16934
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20548 16046 20576 16458
rect 20536 16040 20588 16046
rect 20824 16017 20852 21286
rect 21100 21010 21128 21626
rect 22020 21554 22048 21830
rect 22572 21622 22600 21966
rect 22664 21690 22692 22102
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22664 21350 22692 21626
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 21100 20602 21128 20946
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 21008 18834 21036 19110
rect 21468 19009 21496 21286
rect 21744 21146 21772 21286
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 22480 20602 22508 21286
rect 22756 21146 22784 21830
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21560 19990 21588 20334
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 22376 19984 22428 19990
rect 22376 19926 22428 19932
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 21454 19000 21510 19009
rect 21928 18970 21956 19858
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22296 19378 22324 19790
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22296 19281 22324 19314
rect 22282 19272 22338 19281
rect 22100 19236 22152 19242
rect 22282 19207 22338 19216
rect 22100 19178 22152 19184
rect 21454 18935 21510 18944
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 21008 18426 21036 18770
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21928 18290 21956 18906
rect 22112 18884 22140 19178
rect 22388 19174 22416 19926
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22284 18896 22336 18902
rect 22112 18856 22284 18884
rect 22284 18838 22336 18844
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21928 17814 21956 18226
rect 22008 18148 22060 18154
rect 22008 18090 22060 18096
rect 22020 17814 22048 18090
rect 22296 18086 22324 18838
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22848 18426 22876 18702
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 22284 18080 22336 18086
rect 22284 18022 22336 18028
rect 21916 17808 21968 17814
rect 21916 17750 21968 17756
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21008 17202 21036 17614
rect 22296 17338 22324 18022
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22572 17338 22600 17682
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 21270 17232 21326 17241
rect 20996 17196 21048 17202
rect 21270 17167 21326 17176
rect 21640 17196 21692 17202
rect 20996 17138 21048 17144
rect 21008 16794 21036 17138
rect 21284 17066 21312 17167
rect 21640 17138 21692 17144
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21284 16794 21312 17002
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21652 16726 21680 17138
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21100 16114 21128 16662
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21376 16114 21404 16526
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 20536 15982 20588 15988
rect 20810 16008 20866 16017
rect 20810 15943 20866 15952
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20444 15020 20496 15026
rect 20444 14962 20496 14968
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19996 14618 20024 14962
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20088 14550 20116 14826
rect 19340 14544 19392 14550
rect 19340 14486 19392 14492
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18892 12986 18920 13398
rect 19352 13326 19380 13738
rect 19536 13734 19564 14214
rect 20456 14006 20484 14962
rect 21652 14958 21680 15302
rect 21640 14952 21692 14958
rect 21640 14894 21692 14900
rect 21548 14476 21600 14482
rect 21548 14418 21600 14424
rect 21560 14074 21588 14418
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 21560 13802 21588 14010
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 19076 12918 19104 13262
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 20364 12782 20392 13330
rect 20640 13326 20668 13670
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19076 11898 19104 12242
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19168 11694 19196 12038
rect 20364 11898 20392 12718
rect 20640 12102 20668 13262
rect 21192 13258 21220 13670
rect 21652 13462 21680 14894
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21640 13456 21692 13462
rect 21640 13398 21692 13404
rect 21836 13394 21864 13806
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12170 20760 12718
rect 21192 12306 21220 13194
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12850 21956 13126
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 20720 12164 20772 12170
rect 20772 12124 20852 12152
rect 20720 12106 20772 12112
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20364 11694 20392 11834
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 19168 10470 19196 11086
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19168 10062 19196 10406
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 18656 9880 18736 9908
rect 18604 9862 18656 9868
rect 18248 9654 18276 9862
rect 18616 9722 18644 9862
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18156 9178 18184 9386
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18236 9036 18288 9042
rect 18288 8996 18368 9024
rect 18236 8978 18288 8984
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17788 8294 17816 8910
rect 18340 8294 18368 8996
rect 18616 8838 18644 9658
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18800 8498 18828 9522
rect 19168 9382 19196 9998
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9518 19288 9862
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 17682 7984 17738 7993
rect 16948 7948 17000 7954
rect 17682 7919 17738 7928
rect 16948 7890 17000 7896
rect 16960 7546 16988 7890
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16224 7398 16344 7426
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 6866 16252 7210
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16040 6458 16068 6802
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 16316 6390 16344 7398
rect 17236 7206 17264 7822
rect 17788 7750 17816 8230
rect 18340 7954 18368 8230
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 19168 7886 19196 9318
rect 19260 8838 19288 9454
rect 19352 8838 19380 9590
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19260 8430 19288 8774
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19444 7954 19472 9386
rect 19536 9178 19564 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 9722 20024 10406
rect 20364 10130 20392 11630
rect 20640 11286 20668 12038
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20732 11014 20760 11630
rect 20824 11354 20852 12124
rect 21192 11898 21220 12242
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10606 20760 10950
rect 21192 10674 21220 11834
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21284 11150 21312 11562
rect 21652 11354 21680 12582
rect 22204 11762 22232 15846
rect 22296 15638 22324 17274
rect 23032 17134 23060 21286
rect 23124 19786 23152 22374
rect 23216 22166 23244 22578
rect 23204 22160 23256 22166
rect 23204 22102 23256 22108
rect 23676 21350 23704 23446
rect 23756 22500 23808 22506
rect 23756 22442 23808 22448
rect 23848 22500 23900 22506
rect 23848 22442 23900 22448
rect 23768 22234 23796 22442
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23768 21894 23796 22170
rect 23860 22166 23888 22442
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23952 20330 23980 20946
rect 24044 20942 24072 23446
rect 24136 23186 24164 24074
rect 24228 23322 24256 24686
rect 24688 24614 24716 25298
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24780 24410 24808 25871
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24964 23866 24992 26823
rect 25502 25120 25558 25129
rect 25502 25055 25558 25064
rect 25228 24880 25280 24886
rect 25228 24822 25280 24828
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25148 23866 25176 24210
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24216 23316 24268 23322
rect 24216 23258 24268 23264
rect 24412 23225 24440 23598
rect 24398 23216 24454 23225
rect 24124 23180 24176 23186
rect 24398 23151 24454 23160
rect 24676 23180 24728 23186
rect 24124 23122 24176 23128
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 24766 22944 24822 22953
rect 24766 22879 24822 22888
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 24136 21690 24164 22034
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22879
rect 24124 21684 24176 21690
rect 24124 21626 24176 21632
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24216 21480 24268 21486
rect 25148 21457 25176 23802
rect 25240 22574 25268 24822
rect 25410 24168 25466 24177
rect 25410 24103 25466 24112
rect 25424 22778 25452 24103
rect 25516 23322 25544 25055
rect 25608 24954 25636 27520
rect 27172 25498 27200 27520
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 25596 24948 25648 24954
rect 25596 24890 25648 24896
rect 25504 23316 25556 23322
rect 25504 23258 25556 23264
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 25502 21856 25558 21865
rect 25502 21791 25558 21800
rect 24216 21422 24268 21428
rect 25134 21448 25190 21457
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24044 20602 24072 20742
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 23940 20324 23992 20330
rect 23940 20266 23992 20272
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23112 19780 23164 19786
rect 23112 19722 23164 19728
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23216 19310 23244 19654
rect 23204 19304 23256 19310
rect 23204 19246 23256 19252
rect 23308 18970 23336 20198
rect 23952 19990 23980 20266
rect 24044 20262 24072 20538
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 23400 18834 23428 19110
rect 23388 18828 23440 18834
rect 23388 18770 23440 18776
rect 22560 17128 22612 17134
rect 23020 17128 23072 17134
rect 22560 17070 22612 17076
rect 22926 17096 22982 17105
rect 22468 16720 22520 16726
rect 22468 16662 22520 16668
rect 22480 16182 22508 16662
rect 22468 16176 22520 16182
rect 22468 16118 22520 16124
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22296 14890 22324 15574
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22388 14618 22416 15438
rect 22480 15162 22508 16118
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22388 14006 22416 14554
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22480 12374 22508 13262
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20456 10266 20484 10542
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19536 8362 19564 9114
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19720 8634 19748 8774
rect 20272 8634 20300 9114
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20364 8022 20392 10066
rect 20456 9722 20484 10202
rect 20732 10198 20760 10542
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 20720 10192 20772 10198
rect 20720 10134 20772 10140
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 9722 20944 10066
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20456 9518 20484 9658
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17512 7342 17540 7686
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 16486 6896 16542 6905
rect 16486 6831 16542 6840
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16500 6322 16528 6831
rect 17788 6662 17816 7686
rect 17880 7478 17908 7686
rect 19352 7546 19380 7890
rect 19444 7546 19472 7890
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 16500 5914 16528 6258
rect 16592 6186 16620 6598
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16592 5642 16620 6122
rect 17144 5846 17172 6122
rect 17972 5846 18000 7278
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18340 6186 18368 7142
rect 18800 7002 18828 7278
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 18524 5846 18552 6326
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15672 4826 15700 5034
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 17420 4690 17448 5578
rect 17880 5234 17908 5782
rect 17972 5370 18000 5782
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 4826 17816 4966
rect 18156 4826 18184 5034
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18970 4720 19026 4729
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 17408 4684 17460 4690
rect 18970 4655 18972 4664
rect 17408 4626 17460 4632
rect 19024 4655 19026 4664
rect 18972 4626 19024 4632
rect 15856 4282 15884 4626
rect 17420 4282 17448 4626
rect 18984 4282 19012 4626
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 15750 82 15806 480
rect 15488 54 15806 82
rect 19076 82 19104 6598
rect 19444 6458 19472 6802
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5778 20024 7822
rect 20824 7546 20852 9454
rect 21192 8430 21220 10406
rect 21284 10198 21312 11086
rect 21652 10470 21680 11290
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21836 10266 21864 10542
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21284 7954 21312 9522
rect 21376 9518 21404 10066
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21376 9178 21404 9454
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21468 8498 21496 9998
rect 22190 9616 22246 9625
rect 22190 9551 22246 9560
rect 22204 8974 22232 9551
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22296 9110 22324 9454
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22204 8498 22232 8910
rect 22296 8634 22324 9046
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 21468 8090 21496 8434
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 22020 8022 22048 8366
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20824 7342 20852 7482
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 21732 7268 21784 7274
rect 21732 7210 21784 7216
rect 21744 6866 21772 7210
rect 22020 7206 22048 7958
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22388 7546 22416 7890
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22020 6934 22048 7142
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 22020 6458 22048 6870
rect 22572 6458 22600 17070
rect 23020 17070 23072 17076
rect 22926 17031 22982 17040
rect 22940 16590 22968 17031
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16726 23428 16934
rect 23388 16720 23440 16726
rect 23388 16662 23440 16668
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 22940 15638 22968 16526
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22928 15632 22980 15638
rect 22928 15574 22980 15580
rect 22742 15056 22798 15065
rect 22742 14991 22798 15000
rect 22756 14414 22784 14991
rect 22928 14544 22980 14550
rect 22928 14486 22980 14492
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22756 14074 22784 14350
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22940 13814 22968 14486
rect 23124 13977 23152 15846
rect 23400 15706 23428 16662
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23676 14414 23704 19722
rect 24044 19378 24072 19790
rect 24228 19446 24256 21422
rect 25134 21383 25190 21392
rect 25516 21146 25544 21791
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24492 20324 24544 20330
rect 24492 20266 24544 20272
rect 24504 19990 24532 20266
rect 25148 20262 25176 20946
rect 27620 20936 27672 20942
rect 25410 20904 25466 20913
rect 27620 20878 27672 20884
rect 25410 20839 25466 20848
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25148 20058 25176 20198
rect 25332 20058 25360 20402
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25320 20052 25372 20058
rect 25320 19994 25372 20000
rect 24492 19984 24544 19990
rect 24492 19926 24544 19932
rect 24858 19952 24914 19961
rect 24504 19786 24532 19926
rect 24858 19887 24914 19896
rect 24492 19780 24544 19786
rect 24492 19722 24544 19728
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24216 19440 24268 19446
rect 24216 19382 24268 19388
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23768 18630 23796 19178
rect 24766 19136 24822 19145
rect 24766 19071 24822 19080
rect 24216 18828 24268 18834
rect 24216 18770 24268 18776
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 24228 18086 24256 18770
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 18426 24808 19071
rect 24872 18970 24900 19887
rect 25424 19514 25452 20839
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 24768 18420 24820 18426
rect 24768 18362 24820 18368
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24032 17672 24084 17678
rect 24032 17614 24084 17620
rect 24044 17338 24072 17614
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24044 16998 24072 17274
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24136 16794 24164 17138
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24228 16250 24256 18022
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24780 16590 24808 17206
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 23940 15972 23992 15978
rect 23940 15914 23992 15920
rect 24492 15972 24544 15978
rect 24688 15960 24716 16458
rect 24544 15932 24716 15960
rect 24492 15914 24544 15920
rect 23952 15638 23980 15914
rect 24504 15706 24532 15914
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 23940 15632 23992 15638
rect 23940 15574 23992 15580
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 24228 14958 24256 15302
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24780 15162 24808 15506
rect 24768 15156 24820 15162
rect 24768 15098 24820 15104
rect 24216 14952 24268 14958
rect 24216 14894 24268 14900
rect 24032 14544 24084 14550
rect 24032 14486 24084 14492
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23110 13968 23166 13977
rect 23584 13938 23612 14350
rect 24044 14074 24072 14486
rect 24228 14278 24256 14894
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 14550 24532 14758
rect 24688 14550 24716 14826
rect 24492 14544 24544 14550
rect 24492 14486 24544 14492
rect 24676 14544 24728 14550
rect 24676 14486 24728 14492
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23110 13903 23166 13912
rect 23572 13932 23624 13938
rect 23572 13874 23624 13880
rect 22848 13786 22968 13814
rect 24228 13814 24256 14214
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14486
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24780 14006 24808 14350
rect 24768 14000 24820 14006
rect 24768 13942 24820 13948
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24228 13802 24348 13814
rect 24228 13796 24360 13802
rect 24228 13786 24308 13796
rect 22848 13734 22876 13786
rect 24308 13738 24360 13744
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22744 13524 22796 13530
rect 22744 13466 22796 13472
rect 22756 12646 22784 13466
rect 22848 12986 22876 13670
rect 24320 13530 24348 13738
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24596 13326 24624 13874
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22848 12782 22876 12922
rect 24688 12850 24716 13398
rect 24676 12844 24728 12850
rect 24676 12786 24728 12792
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 24768 12300 24820 12306
rect 24768 12242 24820 12248
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24136 11898 24164 12038
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 23110 11656 23166 11665
rect 23110 11591 23166 11600
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23032 10810 23060 11290
rect 23124 11286 23152 11591
rect 24136 11558 24164 11834
rect 24308 11620 24360 11626
rect 24308 11562 24360 11568
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 23112 11280 23164 11286
rect 23112 11222 23164 11228
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23032 10130 23060 10746
rect 23124 10266 23152 11222
rect 23400 10742 23428 11494
rect 24320 11354 24348 11562
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24780 11286 24808 12242
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 24044 10674 24072 11086
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24780 10810 24808 11222
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23388 10464 23440 10470
rect 23388 10406 23440 10412
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23400 10198 23428 10406
rect 23768 10198 23796 10474
rect 24768 10464 24820 10470
rect 24768 10406 24820 10412
rect 24780 10198 24808 10406
rect 24872 10266 24900 18022
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24964 16726 24992 17682
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24964 16250 24992 16662
rect 25056 16250 25084 18566
rect 25240 17610 25268 19246
rect 25228 17604 25280 17610
rect 25228 17546 25280 17552
rect 27632 16425 27660 20878
rect 27618 16416 27674 16425
rect 27618 16351 27674 16360
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25228 16108 25280 16114
rect 25228 16050 25280 16056
rect 25240 15910 25268 16050
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25872 15904 25924 15910
rect 25872 15846 25924 15852
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25148 12646 25176 13194
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24964 11150 24992 11698
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 23756 10192 23808 10198
rect 23756 10134 23808 10140
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 23020 10124 23072 10130
rect 23020 10066 23072 10072
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 23032 9722 23060 10066
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 10066
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23952 9110 23980 9318
rect 23940 9104 23992 9110
rect 23940 9046 23992 9052
rect 24216 9104 24268 9110
rect 24216 9046 24268 9052
rect 23952 8634 23980 9046
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22020 5846 22048 6394
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 22020 5370 22048 5782
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 22572 5370 22600 5714
rect 22008 5364 22060 5370
rect 22008 5306 22060 5312
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19246 82 19302 480
rect 19076 54 19302 82
rect 22664 82 22692 8502
rect 24044 8498 24072 8910
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24032 8356 24084 8362
rect 24032 8298 24084 8304
rect 24044 8090 24072 8298
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24044 7750 24072 8026
rect 24228 8022 24256 9046
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24688 8498 24716 9658
rect 24964 9178 24992 9862
rect 25148 9722 25176 12582
rect 25240 12442 25268 15846
rect 25884 15065 25912 15846
rect 25870 15056 25926 15065
rect 25870 14991 25926 15000
rect 25412 12912 25464 12918
rect 25412 12854 25464 12860
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 24964 8634 24992 9114
rect 25424 8634 25452 12854
rect 27618 12472 27674 12481
rect 27618 12407 27674 12416
rect 27632 12374 27660 12407
rect 27620 12368 27672 12374
rect 27620 12310 27672 12316
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25516 11898 25544 12242
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25778 10840 25834 10849
rect 25778 10775 25834 10784
rect 25792 10742 25820 10775
rect 25780 10736 25832 10742
rect 25780 10678 25832 10684
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 26160 9897 26188 10066
rect 26146 9888 26202 9897
rect 26146 9823 26202 9832
rect 26160 9722 26188 9823
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 27620 9580 27672 9586
rect 27620 9522 27672 9528
rect 27632 9489 27660 9522
rect 27618 9480 27674 9489
rect 27618 9415 27674 9424
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 24676 8492 24728 8498
rect 24596 8452 24676 8480
rect 24216 8016 24268 8022
rect 24216 7958 24268 7964
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 7342 24072 7686
rect 24228 7546 24256 7958
rect 24596 7886 24624 8452
rect 24676 8434 24728 8440
rect 27618 8392 27674 8401
rect 27618 8327 27674 8336
rect 27632 8294 27660 8327
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 25226 7984 25282 7993
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24688 7410 24716 7958
rect 25226 7919 25282 7928
rect 25240 7546 25268 7919
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 27618 7440 27674 7449
rect 24676 7404 24728 7410
rect 27618 7375 27674 7384
rect 24676 7346 24728 7352
rect 27632 7342 27660 7375
rect 24032 7336 24084 7342
rect 24032 7278 24084 7284
rect 27620 7336 27672 7342
rect 27620 7278 27672 7284
rect 24044 7002 24072 7278
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 24216 6860 24268 6866
rect 24216 6802 24268 6808
rect 23032 6458 23060 6802
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 24136 6458 24164 6734
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 24124 6452 24176 6458
rect 24124 6394 24176 6400
rect 24136 6118 24164 6394
rect 24228 6390 24256 6802
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 6384 24268 6390
rect 24216 6326 24268 6332
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 24228 5914 24256 6326
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23492 5370 23520 5646
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 24044 5166 24072 5510
rect 24228 5370 24256 5850
rect 24596 5710 24624 6258
rect 26054 5944 26110 5953
rect 26054 5879 26110 5888
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24676 5636 24728 5642
rect 24676 5578 24728 5584
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4826 24072 5102
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24044 3942 24072 4762
rect 24412 4758 24440 4966
rect 24688 4758 24716 5578
rect 26068 5370 26096 5879
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 26068 5166 26096 5306
rect 26056 5160 26108 5166
rect 25042 5128 25098 5137
rect 26056 5102 26108 5108
rect 25042 5063 25098 5072
rect 25964 5092 26016 5098
rect 25056 5030 25084 5063
rect 25964 5034 26016 5040
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 24124 4752 24176 4758
rect 24124 4694 24176 4700
rect 24400 4752 24452 4758
rect 24400 4694 24452 4700
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 24136 4282 24164 4694
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24688 4146 24716 4694
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25240 4282 25268 4558
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24308 4004 24360 4010
rect 24308 3946 24360 3952
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24044 3738 24072 3878
rect 24320 3738 24348 3946
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 2854 24716 3334
rect 24676 2848 24728 2854
rect 24676 2790 24728 2796
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1057 24716 2790
rect 25240 2650 25268 4218
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 2310 25176 2450
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25148 2009 25176 2246
rect 25134 2000 25190 2009
rect 25134 1935 25190 1944
rect 24674 1048 24730 1057
rect 24674 983 24730 992
rect 22742 82 22798 480
rect 22664 54 22798 82
rect 25976 82 26004 5034
rect 26238 82 26294 480
rect 25976 54 26294 82
rect 12254 0 12310 54
rect 15750 0 15806 54
rect 19246 0 19302 54
rect 22742 0 22798 54
rect 26238 0 26294 54
<< via2 >>
rect 1306 25608 1362 25664
rect 1122 22072 1178 22128
rect 1122 18536 1178 18592
rect 1950 17040 2006 17096
rect 1766 15000 1822 15056
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 8482 24656 8538 24712
rect 6918 24248 6974 24304
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 9678 19216 9734 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 3882 17176 3938 17232
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 8942 16496 8998 16552
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 3238 15952 3294 16008
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5446 15136 5502 15192
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 1306 11600 1362 11656
rect 2686 11600 2742 11656
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 1214 8064 1270 8120
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 8758 8336 8814 8392
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 7746 6840 7802 6896
rect 1582 4528 1638 4584
rect 1858 2216 1914 2272
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 18602 24656 18658 24712
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 13358 12824 13414 12880
rect 13266 9560 13322 9616
rect 13358 5208 13414 5264
rect 13818 8336 13874 8392
rect 13542 5072 13598 5128
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14738 16532 14740 16552
rect 14740 16532 14792 16552
rect 14792 16532 14794 16552
rect 14738 16496 14794 16532
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15658 12824 15714 12880
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15382 3596 15438 3632
rect 15382 3576 15384 3596
rect 15384 3576 15436 3596
rect 15436 3576 15438 3596
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14738 2488 14794 2544
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19430 24248 19486 24304
rect 18878 23160 18934 23216
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19706 21392 19762 21448
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 17866 15952 17922 16008
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 18878 16632 18934 16688
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 24950 26832 25006 26888
rect 24766 25880 24822 25936
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 21454 18944 21510 19000
rect 22282 19216 22338 19272
rect 21270 17176 21326 17232
rect 20810 15952 20866 16008
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 17682 7928 17738 7984
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 25502 25064 25558 25120
rect 24398 23160 24454 23216
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22888 24822 22944
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25410 24112 25466 24168
rect 25502 21800 25558 21856
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 16486 6840 16542 6896
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 18970 4684 19026 4720
rect 18970 4664 18972 4684
rect 18972 4664 19024 4684
rect 19024 4664 19026 4684
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 22190 9560 22246 9616
rect 22926 17040 22982 17096
rect 22742 15000 22798 15056
rect 25134 21392 25190 21448
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 25410 20848 25466 20904
rect 24858 19896 24914 19952
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 19080 24822 19136
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23110 13912 23166 13968
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23110 11600 23166 11656
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 27618 16360 27674 16416
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 25870 15000 25926 15056
rect 27618 12416 27674 12472
rect 25778 10784 25834 10840
rect 26146 9832 26202 9888
rect 27618 9424 27674 9480
rect 27618 8336 27674 8392
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 25226 7928 25282 7984
rect 27618 7384 27674 7440
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 26054 5888 26110 5944
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25042 5072 25098 5128
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25134 1944 25190 2000
rect 24674 992 24730 1048
<< metal3 >>
rect 27520 27344 28000 27464
rect 24945 26890 25011 26893
rect 27662 26890 27722 27344
rect 24945 26888 27722 26890
rect 24945 26832 24950 26888
rect 25006 26832 27722 26888
rect 24945 26830 27722 26832
rect 24945 26827 25011 26830
rect 27520 26392 28000 26512
rect 0 26120 480 26240
rect 62 25666 122 26120
rect 24761 25938 24827 25941
rect 27662 25938 27722 26392
rect 24761 25936 27722 25938
rect 24761 25880 24766 25936
rect 24822 25880 27722 25936
rect 24761 25878 27722 25880
rect 24761 25875 24827 25878
rect 1301 25666 1367 25669
rect 62 25664 1367 25666
rect 62 25608 1306 25664
rect 1362 25608 1367 25664
rect 62 25606 1367 25608
rect 1301 25603 1367 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 27520 25304 28000 25424
rect 25497 25122 25563 25125
rect 27662 25122 27722 25304
rect 25497 25120 27722 25122
rect 25497 25064 25502 25120
rect 25558 25064 27722 25120
rect 25497 25062 27722 25064
rect 25497 25059 25563 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 8477 24714 8543 24717
rect 18597 24714 18663 24717
rect 8477 24712 18663 24714
rect 8477 24656 8482 24712
rect 8538 24656 18602 24712
rect 18658 24656 18663 24712
rect 8477 24654 18663 24656
rect 8477 24651 8543 24654
rect 18597 24651 18663 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 27520 24352 28000 24472
rect 6913 24306 6979 24309
rect 19425 24306 19491 24309
rect 6913 24304 19491 24306
rect 6913 24248 6918 24304
rect 6974 24248 19430 24304
rect 19486 24248 19491 24304
rect 6913 24246 19491 24248
rect 6913 24243 6979 24246
rect 19425 24243 19491 24246
rect 25405 24170 25471 24173
rect 27662 24170 27722 24352
rect 25405 24168 27722 24170
rect 25405 24112 25410 24168
rect 25466 24112 27722 24168
rect 25405 24110 27722 24112
rect 25405 24107 25471 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 27520 23400 28000 23520
rect 19610 23359 19930 23360
rect 18873 23218 18939 23221
rect 24393 23218 24459 23221
rect 18873 23216 24459 23218
rect 18873 23160 18878 23216
rect 18934 23160 24398 23216
rect 24454 23160 24459 23216
rect 18873 23158 24459 23160
rect 18873 23155 18939 23158
rect 24393 23155 24459 23158
rect 24761 22946 24827 22949
rect 27662 22946 27722 23400
rect 24761 22944 27722 22946
rect 24761 22888 24766 22944
rect 24822 22888 27722 22944
rect 24761 22886 27722 22888
rect 24761 22883 24827 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22584 480 22704
rect 62 22130 122 22584
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 27520 22312 28000 22432
rect 19610 22271 19930 22272
rect 1117 22130 1183 22133
rect 62 22128 1183 22130
rect 62 22072 1122 22128
rect 1178 22072 1183 22128
rect 62 22070 1183 22072
rect 1117 22067 1183 22070
rect 25497 21858 25563 21861
rect 27662 21858 27722 22312
rect 25497 21856 27722 21858
rect 25497 21800 25502 21856
rect 25558 21800 27722 21856
rect 25497 21798 27722 21800
rect 25497 21795 25563 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 19701 21450 19767 21453
rect 25129 21450 25195 21453
rect 19701 21448 25195 21450
rect 19701 21392 19706 21448
rect 19762 21392 25134 21448
rect 25190 21392 25195 21448
rect 19701 21390 25195 21392
rect 19701 21387 19767 21390
rect 25129 21387 25195 21390
rect 27520 21360 28000 21480
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 25405 20906 25471 20909
rect 27662 20906 27722 21360
rect 25405 20904 27722 20906
rect 25405 20848 25410 20904
rect 25466 20848 27722 20904
rect 25405 20846 27722 20848
rect 25405 20843 25471 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 27520 20408 28000 20528
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 24853 19954 24919 19957
rect 27662 19954 27722 20408
rect 24853 19952 27722 19954
rect 24853 19896 24858 19952
rect 24914 19896 27722 19952
rect 24853 19894 27722 19896
rect 24853 19891 24919 19894
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 27520 19320 28000 19440
rect 9673 19274 9739 19277
rect 22277 19274 22343 19277
rect 9673 19272 22343 19274
rect 9673 19216 9678 19272
rect 9734 19216 22282 19272
rect 22338 19216 22343 19272
rect 9673 19214 22343 19216
rect 9673 19211 9739 19214
rect 22277 19211 22343 19214
rect 0 19048 480 19168
rect 24761 19138 24827 19141
rect 27662 19138 27722 19320
rect 24761 19136 27722 19138
rect 24761 19080 24766 19136
rect 24822 19080 27722 19136
rect 24761 19078 27722 19080
rect 24761 19075 24827 19078
rect 10277 19072 10597 19073
rect 62 18594 122 19048
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 21449 19002 21515 19005
rect 21449 19000 27722 19002
rect 21449 18944 21454 19000
rect 21510 18944 27722 19000
rect 21449 18942 27722 18944
rect 21449 18939 21515 18942
rect 1117 18594 1183 18597
rect 62 18592 1183 18594
rect 62 18536 1122 18592
rect 1178 18536 1183 18592
rect 62 18534 1183 18536
rect 1117 18531 1183 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 27662 18488 27722 18942
rect 24277 18463 24597 18464
rect 27520 18368 28000 18488
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17536
rect 24277 17375 24597 17376
rect 3877 17234 3943 17237
rect 21265 17234 21331 17237
rect 3877 17232 21331 17234
rect 3877 17176 3882 17232
rect 3938 17176 21270 17232
rect 21326 17176 21331 17232
rect 3877 17174 21331 17176
rect 3877 17171 3943 17174
rect 21265 17171 21331 17174
rect 1945 17098 2011 17101
rect 22921 17098 22987 17101
rect 1945 17096 22987 17098
rect 1945 17040 1950 17096
rect 2006 17040 22926 17096
rect 22982 17040 22987 17096
rect 1945 17038 22987 17040
rect 1945 17035 2011 17038
rect 22921 17035 22987 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 18873 16690 18939 16693
rect 27662 16690 27722 17416
rect 18873 16688 27722 16690
rect 18873 16632 18878 16688
rect 18934 16632 27722 16688
rect 18873 16630 27722 16632
rect 18873 16627 18939 16630
rect 8937 16554 9003 16557
rect 14733 16554 14799 16557
rect 8937 16552 14799 16554
rect 8937 16496 8942 16552
rect 8998 16496 14738 16552
rect 14794 16496 14799 16552
rect 8937 16494 14799 16496
rect 8937 16491 9003 16494
rect 14733 16491 14799 16494
rect 27520 16416 28000 16448
rect 27520 16360 27618 16416
rect 27674 16360 28000 16416
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 27520 16328 28000 16360
rect 24277 16287 24597 16288
rect 3233 16010 3299 16013
rect 17861 16010 17927 16013
rect 3233 16008 17927 16010
rect 3233 15952 3238 16008
rect 3294 15952 17866 16008
rect 17922 15952 17927 16008
rect 3233 15950 17927 15952
rect 3233 15947 3299 15950
rect 17861 15947 17927 15950
rect 20805 16010 20871 16013
rect 20805 16008 27722 16010
rect 20805 15952 20810 16008
rect 20866 15952 27722 16008
rect 20805 15950 27722 15952
rect 20805 15947 20871 15950
rect 10277 15808 10597 15809
rect 0 15648 480 15768
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 62 15194 122 15648
rect 27662 15496 27722 15950
rect 27520 15376 28000 15496
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 5441 15194 5507 15197
rect 62 15192 5507 15194
rect 62 15136 5446 15192
rect 5502 15136 5507 15192
rect 62 15134 5507 15136
rect 5441 15131 5507 15134
rect 1761 15058 1827 15061
rect 22737 15058 22803 15061
rect 1761 15056 22803 15058
rect 1761 15000 1766 15056
rect 1822 15000 22742 15056
rect 22798 15000 22803 15056
rect 1761 14998 22803 15000
rect 1761 14995 1827 14998
rect 22737 14995 22803 14998
rect 25865 15058 25931 15061
rect 25865 15056 27722 15058
rect 25865 15000 25870 15056
rect 25926 15000 27722 15056
rect 25865 14998 27722 15000
rect 25865 14995 25931 14998
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 27662 14544 27722 14998
rect 27520 14424 28000 14544
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 23105 13970 23171 13973
rect 23105 13968 27722 13970
rect 23105 13912 23110 13968
rect 23166 13912 27722 13968
rect 23105 13910 27722 13912
rect 23105 13907 23171 13910
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 27662 13456 27722 13910
rect 27520 13336 28000 13456
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 13353 12882 13419 12885
rect 15653 12882 15719 12885
rect 13353 12880 15719 12882
rect 13353 12824 13358 12880
rect 13414 12824 15658 12880
rect 15714 12824 15719 12880
rect 13353 12822 15719 12824
rect 13353 12819 13419 12822
rect 15653 12819 15719 12822
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 27520 12472 28000 12504
rect 27520 12416 27618 12472
rect 27674 12416 28000 12472
rect 27520 12384 28000 12416
rect 0 12112 480 12232
rect 62 11658 122 12112
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 1301 11658 1367 11661
rect 62 11656 1367 11658
rect 62 11600 1306 11656
rect 1362 11600 1367 11656
rect 62 11598 1367 11600
rect 1301 11595 1367 11598
rect 2681 11658 2747 11661
rect 23105 11658 23171 11661
rect 2681 11656 23171 11658
rect 2681 11600 2686 11656
rect 2742 11600 23110 11656
rect 23166 11600 23171 11656
rect 2681 11598 23171 11600
rect 2681 11595 2747 11598
rect 23105 11595 23171 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 27520 11296 28000 11416
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 25773 10842 25839 10845
rect 27662 10842 27722 11296
rect 25773 10840 27722 10842
rect 25773 10784 25778 10840
rect 25834 10784 27722 10840
rect 25773 10782 27722 10784
rect 25773 10779 25839 10782
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 27520 10344 28000 10464
rect 19610 10303 19930 10304
rect 26141 9890 26207 9893
rect 27662 9890 27722 10344
rect 26141 9888 27722 9890
rect 26141 9832 26146 9888
rect 26202 9832 27722 9888
rect 26141 9830 27722 9832
rect 26141 9827 26207 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 13261 9618 13327 9621
rect 22185 9618 22251 9621
rect 13261 9616 22251 9618
rect 13261 9560 13266 9616
rect 13322 9560 22190 9616
rect 22246 9560 22251 9616
rect 13261 9558 22251 9560
rect 13261 9555 13327 9558
rect 22185 9555 22251 9558
rect 27520 9480 28000 9512
rect 27520 9424 27618 9480
rect 27674 9424 28000 9480
rect 27520 9392 28000 9424
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 5610 8736 5930 8737
rect 0 8576 480 8696
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 62 8122 122 8576
rect 8753 8394 8819 8397
rect 13813 8394 13879 8397
rect 8753 8392 13879 8394
rect 8753 8336 8758 8392
rect 8814 8336 13818 8392
rect 13874 8336 13879 8392
rect 8753 8334 13879 8336
rect 8753 8331 8819 8334
rect 13813 8331 13879 8334
rect 27520 8392 28000 8424
rect 27520 8336 27618 8392
rect 27674 8336 28000 8392
rect 27520 8304 28000 8336
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 1209 8122 1275 8125
rect 62 8120 1275 8122
rect 62 8064 1214 8120
rect 1270 8064 1275 8120
rect 62 8062 1275 8064
rect 1209 8059 1275 8062
rect 17677 7986 17743 7989
rect 25221 7986 25287 7989
rect 17677 7984 25287 7986
rect 17677 7928 17682 7984
rect 17738 7928 25226 7984
rect 25282 7928 25287 7984
rect 17677 7926 25287 7928
rect 17677 7923 17743 7926
rect 25221 7923 25287 7926
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7440 28000 7472
rect 27520 7384 27618 7440
rect 27674 7384 28000 7440
rect 27520 7352 28000 7384
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 7741 6898 7807 6901
rect 16481 6898 16547 6901
rect 7741 6896 16547 6898
rect 7741 6840 7746 6896
rect 7802 6840 16486 6896
rect 16542 6840 16547 6896
rect 7741 6838 16547 6840
rect 7741 6835 7807 6838
rect 16481 6835 16547 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 27520 6400 28000 6520
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 26049 5946 26115 5949
rect 27662 5946 27722 6400
rect 26049 5944 27722 5946
rect 26049 5888 26054 5944
rect 26110 5888 27722 5944
rect 26049 5886 27722 5888
rect 26049 5883 26115 5886
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 27520 5404 28000 5432
rect 27520 5340 27660 5404
rect 27724 5340 28000 5404
rect 27520 5312 28000 5340
rect 13353 5266 13419 5269
rect 13353 5264 27354 5266
rect 13353 5208 13358 5264
rect 13414 5208 27354 5264
rect 13353 5206 27354 5208
rect 13353 5203 13419 5206
rect 0 5040 480 5160
rect 13537 5130 13603 5133
rect 25037 5130 25103 5133
rect 13537 5128 25103 5130
rect 13537 5072 13542 5128
rect 13598 5072 25042 5128
rect 25098 5072 25103 5128
rect 13537 5070 25103 5072
rect 27294 5130 27354 5206
rect 27654 5130 27660 5132
rect 27294 5070 27660 5130
rect 13537 5067 13603 5070
rect 25037 5067 25103 5070
rect 27654 5068 27660 5070
rect 27724 5068 27730 5132
rect 62 4586 122 5040
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 18965 4722 19031 4725
rect 18965 4720 27722 4722
rect 18965 4664 18970 4720
rect 19026 4664 27722 4720
rect 18965 4662 27722 4664
rect 18965 4659 19031 4662
rect 1577 4586 1643 4589
rect 62 4584 1643 4586
rect 62 4528 1582 4584
rect 1638 4528 1643 4584
rect 62 4526 1643 4528
rect 1577 4523 1643 4526
rect 27662 4480 27722 4662
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4480
rect 24277 4319 24597 4320
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 27654 3770 27660 3772
rect 27294 3710 27660 3770
rect 15377 3634 15443 3637
rect 27294 3634 27354 3710
rect 27654 3708 27660 3710
rect 27724 3708 27730 3772
rect 15377 3632 27354 3634
rect 15377 3576 15382 3632
rect 15438 3576 27354 3632
rect 15377 3574 27354 3576
rect 15377 3571 15443 3574
rect 27520 3500 28000 3528
rect 27520 3436 27660 3500
rect 27724 3436 28000 3500
rect 27520 3408 28000 3436
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 27654 2682 27660 2684
rect 27294 2622 27660 2682
rect 14733 2546 14799 2549
rect 27294 2546 27354 2622
rect 27654 2620 27660 2622
rect 27724 2620 27730 2684
rect 14733 2544 27354 2546
rect 14733 2488 14738 2544
rect 14794 2488 27354 2544
rect 14733 2486 27354 2488
rect 14733 2483 14799 2486
rect 27520 2412 28000 2440
rect 27520 2348 27660 2412
rect 27724 2348 28000 2412
rect 27520 2320 28000 2348
rect 1853 2274 1919 2277
rect 62 2272 1919 2274
rect 62 2216 1858 2272
rect 1914 2216 1919 2272
rect 62 2214 1919 2216
rect 62 1760 122 2214
rect 1853 2211 1919 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 25129 2002 25195 2005
rect 25129 2000 27722 2002
rect 25129 1944 25134 2000
rect 25190 1944 27722 2000
rect 25129 1942 27722 1944
rect 25129 1939 25195 1942
rect 0 1640 480 1760
rect 27662 1488 27722 1942
rect 27520 1368 28000 1488
rect 24669 1050 24735 1053
rect 24669 1048 27722 1050
rect 24669 992 24674 1048
rect 24730 992 27722 1048
rect 24669 990 27722 992
rect 24669 987 24735 990
rect 27662 536 27722 990
rect 27520 416 28000 536
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 27660 5340 27724 5404
rect 27660 5068 27724 5132
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 27660 3708 27724 3772
rect 27660 3436 27724 3500
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 27660 2620 27724 2684
rect 27660 2348 27724 2412
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 27659 5404 27725 5405
rect 27659 5340 27660 5404
rect 27724 5340 27725 5404
rect 27659 5339 27725 5340
rect 27662 5133 27722 5339
rect 27659 5132 27725 5133
rect 27659 5068 27660 5132
rect 27724 5068 27725 5132
rect 27659 5067 27725 5068
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 27659 3772 27725 3773
rect 27659 3708 27660 3772
rect 27724 3708 27725 3772
rect 27659 3707 27725 3708
rect 27662 3501 27722 3707
rect 27659 3500 27725 3501
rect 27659 3436 27660 3500
rect 27724 3436 27725 3500
rect 27659 3435 27725 3436
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 27659 2684 27725 2685
rect 27659 2620 27660 2684
rect 27724 2620 27725 2684
rect 27659 2619 27725 2620
rect 27662 2413 27722 2619
rect 27659 2412 27725 2413
rect 27659 2348 27660 2412
rect 27724 2348 27725 2412
rect 27659 2347 27725 2348
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_0_22 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_30 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_110 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_139
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_151
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_156
timestamp 1586364061
transform 1 0 15456 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_180
timestamp 1586364061
transform 1 0 17664 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_253
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_134
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_157
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_181
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_258
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_270
timestamp 1586364061
transform 1 0 25944 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_274
timestamp 1586364061
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_55
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _173_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_192
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_195
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_239
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_260
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_264
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_3_276
timestamp 1586364061
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_18
timestamp 1586364061
transform 1 0 2760 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_6  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_163
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _177_
timestamp 1586364061
transform 1 0 17296 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_167
timestamp 1586364061
transform 1 0 16468 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_175
timestamp 1586364061
transform 1 0 17204 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_185
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_196
timestamp 1586364061
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 23920 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_2  FILLER_4_250
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_261
timestamp 1586364061
transform 1 0 25116 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_273
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_130
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_134
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_174
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_209
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22724 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_229
timestamp 1586364061
transform 1 0 22172 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_233
timestamp 1586364061
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 23920 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_241
timestamp 1586364061
transform 1 0 23276 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_261
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_268
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_272
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_127
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _222_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 774 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_161
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_165
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_172
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _223_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 590 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_242
timestamp 1586364061
transform 1 0 23368 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_250
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_260
timestamp 1586364061
transform 1 0 25024 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_82
timestamp 1586364061
transform 1 0 8648 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_nor2_4  _107_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_8_181
timestamp 1586364061
transform 1 0 17756 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_242
timestamp 1586364061
transform 1 0 23368 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_248
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_259
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 774 592
use scs8hd_inv_8  _101_
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_70
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_89
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_165
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_181
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 590 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_209
timestamp 1586364061
transform 1 0 20332 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_212
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21988 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_225
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_233
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 774 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 23736 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_241
timestamp 1586364061
transform 1 0 23276 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_255
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_259
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_270
timestamp 1586364061
transform 1 0 25944 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_276
timestamp 1586364061
transform 1 0 26496 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 774 592
use scs8hd_or2_4  _102_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 682 592
use scs8hd_fill_1  FILLER_10_76
timestamp 1586364061
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_8  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_8  _172_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_101
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_8  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _097_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__D
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_or4_4  _166_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_175
timestamp 1586364061
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_192
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_221
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_10_225
timestamp 1586364061
transform 1 0 21804 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_237
timestamp 1586364061
transform 1 0 22908 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_12  FILLER_10_259
timestamp 1586364061
transform 1 0 24932 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_271
timestamp 1586364061
transform 1 0 26036 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_nand2_4  _108_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_103
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 590 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_11_149
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_164
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _099_
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_or4_4  _143_
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_210
timestamp 1586364061
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_256
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_267
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_271
timestamp 1586364061
transform 1 0 26036 0 1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_131
timestamp 1586364061
transform 1 0 13156 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14812 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_151
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_or4_4  _104_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_168
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_172
timestamp 1586364061
transform 1 0 16928 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 222 592
use scs8hd_nand2_4  _138_
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__D
timestamp 1586364061
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_180
timestamp 1586364061
transform 1 0 17664 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__D
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_207
timestamp 1586364061
transform 1 0 20148 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22080 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_237
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_254
timestamp 1586364061
transform 1 0 24472 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_265
timestamp 1586364061
transform 1 0 25484 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_273
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_115
timestamp 1586364061
transform 1 0 11684 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_134
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_138
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_141
timestamp 1586364061
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _109_
timestamp 1586364061
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__D
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _110_
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _115_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_158
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_1  _139_
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__146__D
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_179
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 222 592
use scs8hd_or4_4  _140_
timestamp 1586364061
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use scs8hd_or4_4  _146_
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_183
timestamp 1586364061
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_196
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_194
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_206
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_202
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__C
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _145_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_221
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_228
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_232
timestamp 1586364061
transform 1 0 22448 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_225
timestamp 1586364061
transform 1 0 21804 0 1 9248
box -38 -48 774 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23552 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_241
timestamp 1586364061
transform 1 0 23276 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_242
timestamp 1586364061
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_246
timestamp 1586364061
transform 1 0 23736 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_254
timestamp 1586364061
transform 1 0 24472 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_258
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_14_250
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_256
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_265
timestamp 1586364061
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_267
timestamp 1586364061
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_19
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_31
timestamp 1586364061
transform 1 0 3956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_43
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_15_55
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_102
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 314 592
use scs8hd_or4_4  _118_
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__D
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_or4_4  _157_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__D
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_205
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_221
timestamp 1586364061
transform 1 0 21436 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_258
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_265
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_18
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_127
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__123__C
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__D
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__C
timestamp 1586364061
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__D
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_157
timestamp 1586364061
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_161
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_179
timestamp 1586364061
transform 1 0 17572 0 -1 11424
box -38 -48 222 592
use scs8hd_or4_4  _149_
timestamp 1586364061
transform 1 0 18308 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__D
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_183
timestamp 1586364061
transform 1 0 17940 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_196
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_208
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23000 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_16_247
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_253
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_264
timestamp 1586364061
transform 1 0 25392 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_272
timestamp 1586364061
transform 1 0 26128 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_102
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12604 0 1 11424
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use scs8hd_or4_4  _123_
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_143
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _134_
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__D
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_or4_4  _153_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 20516 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 22540 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_224
timestamp 1586364061
transform 1 0 21712 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 590 592
use scs8hd_decap_4  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_17_274
timestamp 1586364061
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__D
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _126_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  _114_
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_171
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_177
timestamp 1586364061
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use scs8hd_or4_4  _160_
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__C
timestamp 1586364061
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_181
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 20976 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_225
timestamp 1586364061
transform 1 0 21804 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_234
timestamp 1586364061
transform 1 0 22632 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_18_246
timestamp 1586364061
transform 1 0 23736 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_256
timestamp 1586364061
transform 1 0 24656 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_106
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 866 592
use scs8hd_conb_1  _224_
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_128
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_132
timestamp 1586364061
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_148
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__D
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _132_
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_160
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__C
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_or4_4  _130_
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_8  _121_
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_207
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_203
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_205
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_201
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_217
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_221
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_228
timestamp 1586364061
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_262
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_260
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_19_274
timestamp 1586364061
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_272
timestamp 1586364061
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_134
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_195
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_199
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 20792 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_212
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_229
timestamp 1586364061
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_233
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_238
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_242
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_267
timestamp 1586364061
transform 1 0 25668 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_1  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_8  _095_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use scs8hd_buf_1  _129_
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_168
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_174
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_195
timestamp 1586364061
transform 1 0 19044 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_230
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_233
timestamp 1586364061
transform 1 0 22540 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_245
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_249
timestamp 1586364061
transform 1 0 24012 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_262
timestamp 1586364061
transform 1 0 25208 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_45
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_162
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_194
timestamp 1586364061
transform 1 0 18952 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_23_213
timestamp 1586364061
transform 1 0 20700 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 23920 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_261
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 406 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 25484 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_268
timestamp 1586364061
transform 1 0 25760 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_276
timestamp 1586364061
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_132
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_136
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 590 592
use scs8hd_buf_1  _152_
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_165
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_169
timestamp 1586364061
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_176
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 18032 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_203
timestamp 1586364061
transform 1 0 19780 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_206
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22356 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_223
timestamp 1586364061
transform 1 0 21620 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23552 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_246
timestamp 1586364061
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 24104 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25116 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_150
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_154
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_167
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_173
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_177
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_200
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_213
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_217
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21528 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_225
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_229
timestamp 1586364061
transform 1 0 22172 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_255
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_270
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_52
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 774 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 12512 0 1 16864
box -38 -48 866 592
use scs8hd_conb_1  _225_
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_113
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_119
timestamp 1586364061
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_12  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_133
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_148
timestamp 1586364061
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_157
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_161
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_189
timestamp 1586364061
transform 1 0 18492 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_182
timestamp 1586364061
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_205
timestamp 1586364061
transform 1 0 19964 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_3  FILLER_27_194
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_214
timestamp 1586364061
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_224
timestamp 1586364061
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_228
timestamp 1586364061
transform 1 0 22080 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_227
timestamp 1586364061
transform 1 0 21988 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22816 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_245
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_262
timestamp 1586364061
transform 1 0 25208 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 774 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 25576 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_171
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_182
timestamp 1586364061
transform 1 0 17848 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_195
timestamp 1586364061
transform 1 0 19044 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 22448 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_241
timestamp 1586364061
transform 1 0 23276 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_258
timestamp 1586364061
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_270
timestamp 1586364061
transform 1 0 25944 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_274
timestamp 1586364061
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_23
timestamp 1586364061
transform 1 0 3220 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_29
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_45
timestamp 1586364061
transform 1 0 5244 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_nor3_4  _169_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_164
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 20148 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 19964 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_201
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_210
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_227
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_231
timestamp 1586364061
transform 1 0 22356 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_234
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_238
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use scs8hd_decap_8  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _234_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24564 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_259
timestamp 1586364061
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_263
timestamp 1586364061
transform 1 0 25300 0 1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_133
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use scs8hd_nor3_4  _170_
timestamp 1586364061
transform 1 0 15824 0 -1 19040
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_173
timestamp 1586364061
transform 1 0 17020 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_6  FILLER_30_185
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_12  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22448 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_243
timestamp 1586364061
transform 1 0 23460 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_248
timestamp 1586364061
transform 1 0 23920 0 -1 19040
box -38 -48 222 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 24564 0 -1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_252
timestamp 1586364061
transform 1 0 24288 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_259
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_271
timestamp 1586364061
transform 1 0 26036 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_140
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_148
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_152
timestamp 1586364061
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use scs8hd_nor3_4  _171_
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_178
timestamp 1586364061
transform 1 0 17480 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 18492 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 17664 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_182
timestamp 1586364061
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_188
timestamp 1586364061
transform 1 0 18400 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 19688 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_200
timestamp 1586364061
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_204
timestamp 1586364061
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_231
timestamp 1586364061
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_254
timestamp 1586364061
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_258
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_266
timestamp 1586364061
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_270
timestamp 1586364061
transform 1 0 25944 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_276
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_140
timestamp 1586364061
transform 1 0 13984 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_4  FILLER_32_146
timestamp 1586364061
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_150
timestamp 1586364061
transform 1 0 14904 0 -1 20128
box -38 -48 130 592
use scs8hd_nor3_4  _168_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _164_
timestamp 1586364061
transform 1 0 17296 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_167
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_185
timestamp 1586364061
transform 1 0 18124 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_189
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_32_221
timestamp 1586364061
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22172 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21620 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_225
timestamp 1586364061
transform 1 0 21804 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_238
timestamp 1586364061
transform 1 0 23000 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_242
timestamp 1586364061
transform 1 0 23368 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_255
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 774 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_266
timestamp 1586364061
transform 1 0 25576 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_6
timestamp 1586364061
transform 1 0 1656 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_19
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_18
timestamp 1586364061
transform 1 0 2760 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_50
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11776 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_113
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_136
timestamp 1586364061
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_133
timestamp 1586364061
transform 1 0 13340 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_140
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15824 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_155
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_171
timestamp 1586364061
transform 1 0 16836 0 -1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 18216 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_183
timestamp 1586364061
transform 1 0 17940 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_188
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_195
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_199
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_200
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_205
timestamp 1586364061
transform 1 0 19964 0 -1 21216
box -38 -48 590 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 21160 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_214
timestamp 1586364061
transform 1 0 20792 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_218
timestamp 1586364061
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_211
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 22724 0 -1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_33_233
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 774 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 23736 0 -1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_237
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_238
timestamp 1586364061
transform 1 0 23000 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_33_259
timestamp 1586364061
transform 1 0 24932 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_255
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 774 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25300 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_265
timestamp 1586364061
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_267
timestamp 1586364061
transform 1 0 25668 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 590 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_152
timestamp 1586364061
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_163
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_167
timestamp 1586364061
transform 1 0 16468 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_188
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_192
timestamp 1586364061
transform 1 0 18768 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_207
timestamp 1586364061
transform 1 0 20148 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_222
timestamp 1586364061
transform 1 0 21528 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_235
timestamp 1586364061
transform 1 0 22724 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22908 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 24012 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_239
timestamp 1586364061
transform 1 0 23092 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 406 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_251
timestamp 1586364061
transform 1 0 24196 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 774 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_139
timestamp 1586364061
transform 1 0 13892 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_8  _207_
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_157
timestamp 1586364061
transform 1 0 15548 0 -1 22304
box -38 -48 590 592
use scs8hd_decap_8  FILLER_36_174
timestamp 1586364061
transform 1 0 17112 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_4  FILLER_36_191
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_195
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_198
timestamp 1586364061
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_224
timestamp 1586364061
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_228
timestamp 1586364061
transform 1 0 22080 0 -1 22304
box -38 -48 406 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 24012 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_241
timestamp 1586364061
transform 1 0 23276 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_247
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_258
timestamp 1586364061
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_270
timestamp 1586364061
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_274
timestamp 1586364061
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_128
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14444 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_139
timestamp 1586364061
transform 1 0 13892 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_154
timestamp 1586364061
transform 1 0 15272 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_198
timestamp 1586364061
transform 1 0 19320 0 1 22304
box -38 -48 314 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 21160 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 20792 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_212
timestamp 1586364061
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_216
timestamp 1586364061
transform 1 0 20976 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_229
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 314 592
use scs8hd_decap_4  FILLER_37_234
timestamp 1586364061
transform 1 0 22632 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_270
timestamp 1586364061
transform 1 0 25944 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_147
timestamp 1586364061
transform 1 0 14628 0 -1 23392
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16008 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_165
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 17020 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_182
timestamp 1586364061
transform 1 0 17848 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19136 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_205
timestamp 1586364061
transform 1 0 19964 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_209
timestamp 1586364061
transform 1 0 20332 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_224
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  FILLER_38_229
timestamp 1586364061
transform 1 0 22172 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_235
timestamp 1586364061
transform 1 0 22724 0 -1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_243
timestamp 1586364061
transform 1 0 23460 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_247
timestamp 1586364061
transform 1 0 23828 0 -1 23392
box -38 -48 774 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_14
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_26
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_38
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_50
timestamp 1586364061
transform 1 0 5704 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_58
timestamp 1586364061
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_113
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_117
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_121
timestamp 1586364061
transform 1 0 12236 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 13156 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 13708 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_127
timestamp 1586364061
transform 1 0 12788 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_130
timestamp 1586364061
transform 1 0 13064 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_39_139
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_151
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_151
timestamp 1586364061
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 15180 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_155
timestamp 1586364061
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_163
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17112 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_170
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_177
timestamp 1586364061
transform 1 0 17388 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 18124 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 18676 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_189
timestamp 1586364061
transform 1 0 18492 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_193
timestamp 1586364061
transform 1 0 18860 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_199
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_200
timestamp 1586364061
transform 1 0 19504 0 -1 24480
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_218
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_208
timestamp 1586364061
transform 1 0 20240 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_211
timestamp 1586364061
transform 1 0 20516 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_226
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_231
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_235
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_224
timestamp 1586364061
transform 1 0 21712 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_249
timestamp 1586364061
transform 1 0 24012 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_243
timestamp 1586364061
transform 1 0 23460 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_247
timestamp 1586364061
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_259
timestamp 1586364061
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_271
timestamp 1586364061
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 16928 0 1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18768 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_190
timestamp 1586364061
transform 1 0 18584 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_194
timestamp 1586364061
transform 1 0 18952 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_198
timestamp 1586364061
transform 1 0 19320 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_202
timestamp 1586364061
transform 1 0 19688 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_206
timestamp 1586364061
transform 1 0 20056 0 1 24480
box -38 -48 406 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 20424 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_213
timestamp 1586364061
transform 1 0 20700 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_225
timestamp 1586364061
transform 1 0 21804 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_259
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_263
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_41_275
timestamp 1586364061
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_6  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_259
timestamp 1586364061
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_271
timestamp 1586364061
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
<< labels >>
rlabel metal2 s 5262 0 5318 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8758 0 8814 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 12254 0 12310 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15750 0 15806 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 19246 0 19302 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 22742 0 22798 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[0]
port 6 nsew default input
rlabel metal3 s 27520 2320 28000 2440 6 chanx_right_in[1]
port 7 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 chanx_right_in[2]
port 8 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[3]
port 9 nsew default input
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_in[4]
port 10 nsew default input
rlabel metal3 s 27520 6400 28000 6520 6 chanx_right_in[5]
port 11 nsew default input
rlabel metal3 s 27520 7352 28000 7472 6 chanx_right_in[6]
port 12 nsew default input
rlabel metal3 s 27520 8304 28000 8424 6 chanx_right_in[7]
port 13 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[8]
port 14 nsew default input
rlabel metal3 s 27520 19320 28000 19440 6 chanx_right_out[0]
port 15 nsew default tristate
rlabel metal3 s 27520 20408 28000 20528 6 chanx_right_out[1]
port 16 nsew default tristate
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_out[2]
port 17 nsew default tristate
rlabel metal3 s 27520 22312 28000 22432 6 chanx_right_out[3]
port 18 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chanx_right_out[4]
port 19 nsew default tristate
rlabel metal3 s 27520 24352 28000 24472 6 chanx_right_out[5]
port 20 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[6]
port 21 nsew default tristate
rlabel metal3 s 27520 26392 28000 26512 6 chanx_right_out[7]
port 22 nsew default tristate
rlabel metal3 s 27520 27344 28000 27464 6 chanx_right_out[8]
port 23 nsew default tristate
rlabel metal2 s 754 27520 810 28000 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 2226 27520 2282 28000 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal2 s 8482 27520 8538 28000 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 10046 27520 10102 28000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal2 s 11610 27520 11666 28000 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 13174 27520 13230 28000 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 14738 27520 14794 28000 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 19338 27520 19394 28000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal2 s 24030 27520 24086 28000 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal2 s 25594 27520 25650 28000 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 27158 27520 27214 28000 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 26238 0 26294 480 6 data_in
port 42 nsew default input
rlabel metal2 s 1766 0 1822 480 6 enable
port 43 nsew default input
rlabel metal3 s 27520 16328 28000 16448 6 right_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 27520 17416 28000 17536 6 right_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal3 s 27520 18368 28000 18488 6 right_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 right_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal3 s 27520 12384 28000 12504 6 right_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 right_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal3 s 27520 14424 28000 14544 6 right_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 right_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 27520 10344 28000 10464 6 right_top_grid_pin_10_
port 52 nsew default input
rlabel metal3 s 0 19048 480 19168 6 top_left_grid_pin_11_
port 53 nsew default input
rlabel metal3 s 0 22584 480 22704 6 top_left_grid_pin_13_
port 54 nsew default input
rlabel metal3 s 0 26120 480 26240 6 top_left_grid_pin_15_
port 55 nsew default input
rlabel metal3 s 0 1640 480 1760 6 top_left_grid_pin_1_
port 56 nsew default input
rlabel metal3 s 0 5040 480 5160 6 top_left_grid_pin_3_
port 57 nsew default input
rlabel metal3 s 0 8576 480 8696 6 top_left_grid_pin_5_
port 58 nsew default input
rlabel metal3 s 0 12112 480 12232 6 top_left_grid_pin_7_
port 59 nsew default input
rlabel metal3 s 0 15648 480 15768 6 top_left_grid_pin_9_
port 60 nsew default input
rlabel metal3 s 27520 416 28000 536 6 top_right_grid_pin_11_
port 61 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 62 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 63 nsew default input
<< end >>
