magic
tech EFS8A
magscale 1 2
timestamp 1602524676
<< locali >>
rect 9275 18377 9321 18411
rect 9631 17697 9758 17731
rect 7199 16983 7233 17051
rect 7199 16949 7205 16983
rect 10051 13481 10057 13515
rect 10051 13413 10085 13481
rect 9976 12325 10044 12359
rect 10051 11305 10057 11339
rect 10051 11237 10085 11305
rect 8953 10523 8987 10693
rect 11287 10081 11322 10115
rect 11563 8993 11598 9027
<< viali >>
rect 2053 34697 2087 34731
rect 10885 34697 10919 34731
rect 1593 34629 1627 34663
rect 8263 34561 8297 34595
rect 1409 34493 1443 34527
rect 8176 34493 8210 34527
rect 10701 34493 10735 34527
rect 11253 34493 11287 34527
rect 8677 34357 8711 34391
rect 5365 29801 5399 29835
rect 5181 29665 5215 29699
rect 5181 28985 5215 29019
rect 13645 28713 13679 28747
rect 13461 28577 13495 28611
rect 13461 27829 13495 27863
rect 4629 26537 4663 26571
rect 4445 26401 4479 26435
rect 4537 25653 4571 25687
rect 1409 22049 1443 22083
rect 1593 21845 1627 21879
rect 1593 21641 1627 21675
rect 6352 19873 6386 19907
rect 6423 19669 6457 19703
rect 6929 19669 6963 19703
rect 5273 19465 5307 19499
rect 6377 19465 6411 19499
rect 7205 19329 7239 19363
rect 5089 19261 5123 19295
rect 6929 19193 6963 19227
rect 7021 19193 7055 19227
rect 5641 19125 5675 19159
rect 9873 18921 9907 18955
rect 6009 18853 6043 18887
rect 6837 18853 6871 18887
rect 7573 18853 7607 18887
rect 4880 18785 4914 18819
rect 9689 18785 9723 18819
rect 5917 18717 5951 18751
rect 6193 18717 6227 18751
rect 7481 18717 7515 18751
rect 8033 18649 8067 18683
rect 4951 18581 4985 18615
rect 5365 18581 5399 18615
rect 5733 18581 5767 18615
rect 4307 18377 4341 18411
rect 9321 18377 9355 18411
rect 4721 18309 4755 18343
rect 5273 18241 5307 18275
rect 8033 18241 8067 18275
rect 8953 18241 8987 18275
rect 4236 18173 4270 18207
rect 9172 18173 9206 18207
rect 5365 18105 5399 18139
rect 5917 18105 5951 18139
rect 7021 18105 7055 18139
rect 7665 18105 7699 18139
rect 7757 18105 7791 18139
rect 5089 18037 5123 18071
rect 6193 18037 6227 18071
rect 6653 18037 6687 18071
rect 7481 18037 7515 18071
rect 9689 18037 9723 18071
rect 6009 17833 6043 17867
rect 9827 17833 9861 17867
rect 5181 17765 5215 17799
rect 6745 17765 6779 17799
rect 1409 17697 1443 17731
rect 3024 17697 3058 17731
rect 9597 17697 9631 17731
rect 11437 17697 11471 17731
rect 3111 17629 3145 17663
rect 5089 17629 5123 17663
rect 6653 17629 6687 17663
rect 6929 17629 6963 17663
rect 7941 17629 7975 17663
rect 8125 17629 8159 17663
rect 1593 17561 1627 17595
rect 5641 17561 5675 17595
rect 7665 17493 7699 17527
rect 11621 17493 11655 17527
rect 1593 17289 1627 17323
rect 2973 17289 3007 17323
rect 6193 17289 6227 17323
rect 7757 17289 7791 17323
rect 8401 17289 8435 17323
rect 11437 17289 11471 17323
rect 4307 17221 4341 17255
rect 8033 17221 8067 17255
rect 5273 17153 5307 17187
rect 5917 17153 5951 17187
rect 8677 17153 8711 17187
rect 9321 17153 9355 17187
rect 4236 17085 4270 17119
rect 6837 17085 6871 17119
rect 5089 17017 5123 17051
rect 5365 17017 5399 17051
rect 8769 17017 8803 17051
rect 4721 16949 4755 16983
rect 6653 16949 6687 16983
rect 7205 16949 7239 16983
rect 9689 16949 9723 16983
rect 4813 16745 4847 16779
rect 6285 16745 6319 16779
rect 8033 16745 8067 16779
rect 5686 16677 5720 16711
rect 7434 16677 7468 16711
rect 5365 16541 5399 16575
rect 7113 16541 7147 16575
rect 5273 16405 5307 16439
rect 6837 16405 6871 16439
rect 8585 16405 8619 16439
rect 5917 16201 5951 16235
rect 8217 16201 8251 16235
rect 4997 15997 5031 16031
rect 7297 15997 7331 16031
rect 4905 15929 4939 15963
rect 5359 15929 5393 15963
rect 6285 15929 6319 15963
rect 7618 15929 7652 15963
rect 4537 15861 4571 15895
rect 6653 15861 6687 15895
rect 7205 15861 7239 15895
rect 6377 15657 6411 15691
rect 5778 15589 5812 15623
rect 5457 15453 5491 15487
rect 8309 15453 8343 15487
rect 4997 15317 5031 15351
rect 7205 15317 7239 15351
rect 7481 15317 7515 15351
rect 5549 15113 5583 15147
rect 8309 15113 8343 15147
rect 8585 14977 8619 15011
rect 8861 14977 8895 15011
rect 8033 14841 8067 14875
rect 8677 14841 8711 14875
rect 5917 14773 5951 14807
rect 8677 14569 8711 14603
rect 13645 14569 13679 14603
rect 8119 14501 8153 14535
rect 9873 14501 9907 14535
rect 13461 14433 13495 14467
rect 7757 14365 7791 14399
rect 9781 14365 9815 14399
rect 10333 14297 10367 14331
rect 6929 14229 6963 14263
rect 7297 14229 7331 14263
rect 11253 14025 11287 14059
rect 8217 13957 8251 13991
rect 8953 13957 8987 13991
rect 9781 13889 9815 13923
rect 10241 13889 10275 13923
rect 6837 13821 6871 13855
rect 7297 13821 7331 13855
rect 7757 13821 7791 13855
rect 8033 13821 8067 13855
rect 9965 13753 9999 13787
rect 10057 13753 10091 13787
rect 13461 13753 13495 13787
rect 6193 13685 6227 13719
rect 6653 13685 6687 13719
rect 8677 13685 8711 13719
rect 9413 13685 9447 13719
rect 10977 13685 11011 13719
rect 10057 13481 10091 13515
rect 10609 13481 10643 13515
rect 6285 13413 6319 13447
rect 11621 13413 11655 13447
rect 12173 13413 12207 13447
rect 4537 13345 4571 13379
rect 5273 13345 5307 13379
rect 7021 13345 7055 13379
rect 7205 13345 7239 13379
rect 7573 13345 7607 13379
rect 7941 13345 7975 13379
rect 5917 13277 5951 13311
rect 8217 13277 8251 13311
rect 9689 13277 9723 13311
rect 11529 13277 11563 13311
rect 6653 13141 6687 13175
rect 8493 13141 8527 13175
rect 9229 13141 9263 13175
rect 10701 12937 10735 12971
rect 11713 12937 11747 12971
rect 12587 12937 12621 12971
rect 3985 12801 4019 12835
rect 11437 12801 11471 12835
rect 4629 12733 4663 12767
rect 5181 12733 5215 12767
rect 5273 12733 5307 12767
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 7297 12733 7331 12767
rect 7665 12733 7699 12767
rect 8033 12733 8067 12767
rect 9137 12733 9171 12767
rect 10057 12733 10091 12767
rect 10952 12733 10986 12767
rect 12484 12733 12518 12767
rect 12909 12733 12943 12767
rect 8585 12665 8619 12699
rect 9499 12665 9533 12699
rect 4353 12597 4387 12631
rect 4721 12597 4755 12631
rect 6193 12597 6227 12631
rect 6561 12597 6595 12631
rect 7113 12597 7147 12631
rect 9045 12597 9079 12631
rect 10333 12597 10367 12631
rect 11023 12597 11057 12631
rect 12173 12597 12207 12631
rect 6469 12393 6503 12427
rect 9137 12393 9171 12427
rect 10609 12393 10643 12427
rect 13645 12393 13679 12427
rect 9942 12325 9976 12359
rect 11529 12325 11563 12359
rect 11621 12325 11655 12359
rect 5181 12257 5215 12291
rect 6101 12257 6135 12291
rect 6469 12257 6503 12291
rect 6653 12257 6687 12291
rect 7113 12257 7147 12291
rect 7389 12257 7423 12291
rect 8620 12257 8654 12291
rect 13461 12257 13495 12291
rect 9689 12189 9723 12223
rect 4997 12121 5031 12155
rect 8723 12121 8757 12155
rect 12081 12121 12115 12155
rect 4537 12053 4571 12087
rect 5365 12053 5399 12087
rect 5733 12053 5767 12087
rect 7941 12053 7975 12087
rect 8309 12053 8343 12087
rect 11621 11849 11655 11883
rect 12173 11849 12207 11883
rect 13461 11849 13495 11883
rect 3985 11781 4019 11815
rect 6285 11713 6319 11747
rect 12817 11713 12851 11747
rect 4445 11645 4479 11679
rect 5181 11645 5215 11679
rect 5273 11645 5307 11679
rect 5641 11645 5675 11679
rect 6837 11645 6871 11679
rect 7297 11645 7331 11679
rect 7665 11645 7699 11679
rect 8033 11645 8067 11679
rect 8953 11645 8987 11679
rect 9137 11645 9171 11679
rect 9873 11645 9907 11679
rect 9965 11645 9999 11679
rect 10333 11645 10367 11679
rect 10885 11645 10919 11679
rect 11253 11577 11287 11611
rect 12541 11577 12575 11611
rect 12633 11577 12667 11611
rect 3617 11509 3651 11543
rect 4353 11509 4387 11543
rect 4537 11509 4571 11543
rect 6561 11509 6595 11543
rect 6929 11509 6963 11543
rect 8585 11509 8619 11543
rect 9413 11509 9447 11543
rect 3801 11305 3835 11339
rect 4445 11305 4479 11339
rect 5273 11305 5307 11339
rect 6837 11305 6871 11339
rect 9137 11305 9171 11339
rect 10057 11305 10091 11339
rect 11253 11305 11287 11339
rect 7481 11237 7515 11271
rect 8217 11237 8251 11271
rect 11621 11237 11655 11271
rect 4629 11169 4663 11203
rect 5641 11169 5675 11203
rect 6101 11169 6135 11203
rect 6653 11169 6687 11203
rect 7021 11169 7055 11203
rect 10609 11169 10643 11203
rect 8125 11101 8159 11135
rect 8769 11101 8803 11135
rect 9689 11101 9723 11135
rect 11529 11101 11563 11135
rect 11805 11101 11839 11135
rect 4813 11033 4847 11067
rect 7849 10965 7883 10999
rect 10885 10965 10919 10999
rect 12449 10965 12483 10999
rect 5917 10761 5951 10795
rect 6285 10761 6319 10795
rect 10149 10761 10183 10795
rect 11115 10761 11149 10795
rect 12173 10761 12207 10795
rect 8953 10693 8987 10727
rect 9045 10693 9079 10727
rect 11805 10693 11839 10727
rect 4813 10625 4847 10659
rect 8401 10625 8435 10659
rect 4905 10557 4939 10591
rect 6653 10557 6687 10591
rect 7205 10557 7239 10591
rect 7665 10557 7699 10591
rect 7757 10557 7791 10591
rect 8125 10557 8159 10591
rect 10793 10625 10827 10659
rect 9229 10557 9263 10591
rect 11044 10557 11078 10591
rect 8953 10489 8987 10523
rect 9550 10489 9584 10523
rect 10425 10489 10459 10523
rect 4261 10421 4295 10455
rect 4629 10421 4663 10455
rect 8677 10421 8711 10455
rect 11529 10421 11563 10455
rect 5641 10217 5675 10251
rect 8585 10217 8619 10251
rect 8861 10217 8895 10251
rect 11391 10217 11425 10251
rect 5365 10149 5399 10183
rect 8217 10149 8251 10183
rect 9229 10149 9263 10183
rect 9781 10149 9815 10183
rect 9873 10149 9907 10183
rect 10425 10149 10459 10183
rect 6745 10081 6779 10115
rect 7481 10081 7515 10115
rect 7573 10081 7607 10115
rect 8033 10081 8067 10115
rect 11253 10081 11287 10115
rect 4905 9877 4939 9911
rect 6285 9877 6319 9911
rect 6653 9877 6687 9911
rect 5273 9673 5307 9707
rect 5641 9673 5675 9707
rect 8953 9673 8987 9707
rect 10241 9673 10275 9707
rect 6653 9605 6687 9639
rect 10563 9605 10597 9639
rect 8309 9537 8343 9571
rect 5733 9469 5767 9503
rect 6837 9469 6871 9503
rect 7573 9469 7607 9503
rect 7757 9469 7791 9503
rect 8033 9469 8067 9503
rect 8585 9469 8619 9503
rect 9480 9469 9514 9503
rect 9873 9469 9907 9503
rect 10460 9469 10494 9503
rect 10885 9469 10919 9503
rect 5917 9333 5951 9367
rect 6193 9333 6227 9367
rect 9551 9333 9585 9367
rect 11345 9333 11379 9367
rect 6745 9129 6779 9163
rect 8585 9129 8619 9163
rect 9505 9129 9539 9163
rect 11667 9129 11701 9163
rect 12679 9129 12713 9163
rect 8309 9061 8343 9095
rect 5641 8993 5675 9027
rect 7205 8993 7239 9027
rect 7665 8993 7699 9027
rect 10333 8993 10367 9027
rect 11529 8993 11563 9027
rect 12587 8993 12621 9027
rect 6009 8925 6043 8959
rect 6377 8925 6411 8959
rect 7757 8925 7791 8959
rect 9045 8857 9079 8891
rect 4905 8789 4939 8823
rect 5273 8789 5307 8823
rect 5779 8789 5813 8823
rect 5917 8789 5951 8823
rect 9965 8789 9999 8823
rect 6653 8585 6687 8619
rect 9873 8585 9907 8619
rect 10977 8585 11011 8619
rect 13645 8585 13679 8619
rect 4353 8517 4387 8551
rect 5319 8517 5353 8551
rect 5457 8517 5491 8551
rect 5549 8449 5583 8483
rect 5917 8449 5951 8483
rect 8493 8449 8527 8483
rect 8769 8449 8803 8483
rect 9505 8449 9539 8483
rect 10057 8449 10091 8483
rect 12449 8449 12483 8483
rect 4721 8381 4755 8415
rect 6837 8381 6871 8415
rect 7297 8381 7331 8415
rect 13461 8381 13495 8415
rect 14013 8381 14047 8415
rect 5181 8313 5215 8347
rect 6193 8313 6227 8347
rect 7573 8313 7607 8347
rect 8585 8313 8619 8347
rect 10149 8313 10183 8347
rect 10701 8313 10735 8347
rect 12909 8313 12943 8347
rect 5089 8245 5123 8279
rect 7849 8245 7883 8279
rect 8309 8245 8343 8279
rect 11529 8245 11563 8279
rect 4537 8041 4571 8075
rect 7297 8041 7331 8075
rect 8769 8041 8803 8075
rect 8170 7973 8204 8007
rect 9873 7973 9907 8007
rect 10425 7973 10459 8007
rect 11437 7973 11471 8007
rect 4353 7905 4387 7939
rect 5365 7905 5399 7939
rect 5512 7837 5546 7871
rect 5733 7837 5767 7871
rect 7849 7837 7883 7871
rect 9781 7837 9815 7871
rect 11345 7837 11379 7871
rect 12817 7837 12851 7871
rect 4905 7769 4939 7803
rect 5825 7769 5859 7803
rect 6929 7769 6963 7803
rect 11897 7769 11931 7803
rect 5273 7701 5307 7735
rect 5641 7701 5675 7735
rect 6377 7701 6411 7735
rect 7665 7701 7699 7735
rect 5641 7497 5675 7531
rect 6561 7497 6595 7531
rect 9781 7497 9815 7531
rect 11805 7497 11839 7531
rect 3525 7429 3559 7463
rect 12587 7429 12621 7463
rect 4353 7361 4387 7395
rect 8493 7361 8527 7395
rect 11069 7361 11103 7395
rect 3617 7293 3651 7327
rect 4169 7293 4203 7327
rect 4721 7293 4755 7327
rect 5457 7293 5491 7327
rect 9413 7293 9447 7327
rect 10149 7293 10183 7327
rect 12516 7293 12550 7327
rect 12909 7293 12943 7327
rect 7021 7225 7055 7259
rect 7113 7225 7147 7259
rect 7665 7225 7699 7259
rect 8814 7225 8848 7259
rect 10425 7225 10459 7259
rect 10517 7225 10551 7259
rect 5089 7157 5123 7191
rect 6193 7157 6227 7191
rect 7941 7157 7975 7191
rect 8309 7157 8343 7191
rect 11437 7157 11471 7191
rect 3709 6953 3743 6987
rect 5365 6953 5399 6987
rect 7021 6953 7055 6987
rect 7389 6953 7423 6987
rect 7757 6953 7791 6987
rect 9045 6953 9079 6987
rect 11529 6953 11563 6987
rect 6193 6885 6227 6919
rect 8170 6885 8204 6919
rect 9873 6885 9907 6919
rect 10425 6885 10459 6919
rect 10701 6885 10735 6919
rect 4445 6817 4479 6851
rect 5457 6817 5491 6851
rect 8769 6817 8803 6851
rect 11345 6817 11379 6851
rect 5825 6749 5859 6783
rect 7849 6749 7883 6783
rect 9413 6749 9447 6783
rect 9781 6749 9815 6783
rect 5622 6681 5656 6715
rect 4629 6613 4663 6647
rect 5733 6613 5767 6647
rect 6561 6409 6595 6443
rect 8585 6409 8619 6443
rect 10793 6409 10827 6443
rect 11253 6409 11287 6443
rect 7021 6341 7055 6375
rect 10425 6341 10459 6375
rect 11483 6341 11517 6375
rect 5181 6273 5215 6307
rect 7665 6273 7699 6307
rect 9321 6273 9355 6307
rect 5273 6205 5307 6239
rect 6193 6205 6227 6239
rect 8861 6205 8895 6239
rect 11380 6205 11414 6239
rect 11805 6205 11839 6239
rect 4537 6137 4571 6171
rect 7573 6137 7607 6171
rect 7986 6137 8020 6171
rect 9873 6137 9907 6171
rect 9965 6137 9999 6171
rect 5089 6069 5123 6103
rect 9689 6069 9723 6103
rect 5089 5865 5123 5899
rect 6377 5865 6411 5899
rect 8309 5865 8343 5899
rect 9505 5865 9539 5899
rect 9689 5797 9723 5831
rect 4905 5729 4939 5763
rect 6561 5729 6595 5763
rect 8125 5729 8159 5763
rect 10333 5729 10367 5763
rect 5457 5525 5491 5559
rect 7297 5525 7331 5559
rect 7757 5525 7791 5559
rect 4905 5321 4939 5355
rect 7021 5321 7055 5355
rect 8217 5321 8251 5355
rect 9643 5321 9677 5355
rect 10333 5321 10367 5355
rect 6561 5185 6595 5219
rect 7849 5185 7883 5219
rect 5800 5117 5834 5151
rect 7205 5117 7239 5151
rect 7665 5117 7699 5151
rect 9572 5117 9606 5151
rect 6285 5049 6319 5083
rect 5871 4981 5905 5015
rect 10057 4981 10091 5015
rect 7297 4777 7331 4811
rect 9827 4777 9861 4811
rect 5549 4641 5583 4675
rect 6193 4641 6227 4675
rect 6377 4641 6411 4675
rect 6745 4641 6779 4675
rect 8493 4641 8527 4675
rect 9756 4641 9790 4675
rect 7021 4573 7055 4607
rect 5365 4437 5399 4471
rect 8125 4437 8159 4471
rect 4905 4233 4939 4267
rect 5181 4233 5215 4267
rect 6561 4233 6595 4267
rect 9597 4233 9631 4267
rect 10701 4233 10735 4267
rect 7113 4097 7147 4131
rect 5549 4029 5583 4063
rect 6193 4029 6227 4063
rect 10200 4029 10234 4063
rect 5365 3961 5399 3995
rect 7205 3961 7239 3995
rect 7757 3961 7791 3995
rect 8125 3961 8159 3995
rect 8677 3961 8711 3995
rect 8769 3961 8803 3995
rect 9321 3961 9355 3995
rect 9965 3961 9999 3995
rect 5641 3893 5675 3927
rect 8493 3893 8527 3927
rect 10287 3893 10321 3927
rect 7573 3689 7607 3723
rect 11253 3689 11287 3723
rect 7297 3621 7331 3655
rect 8078 3621 8112 3655
rect 9689 3621 9723 3655
rect 5457 3553 5491 3587
rect 6193 3553 6227 3587
rect 6285 3553 6319 3587
rect 6653 3553 6687 3587
rect 7757 3553 7791 3587
rect 8677 3553 8711 3587
rect 9781 3553 9815 3587
rect 8953 3485 8987 3519
rect 6837 3417 6871 3451
rect 5273 3349 5307 3383
rect 4721 3145 4755 3179
rect 5089 3145 5123 3179
rect 7757 3145 7791 3179
rect 8493 3145 8527 3179
rect 9781 3145 9815 3179
rect 10701 3145 10735 3179
rect 6561 3077 6595 3111
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 8677 3009 8711 3043
rect 9321 3009 9355 3043
rect 5273 2941 5307 2975
rect 8033 2941 8067 2975
rect 10149 2941 10183 2975
rect 13461 2941 13495 2975
rect 7158 2873 7192 2907
rect 8769 2873 8803 2907
rect 6193 2805 6227 2839
rect 10333 2805 10367 2839
rect 13645 2805 13679 2839
rect 14105 2805 14139 2839
rect 5641 2601 5675 2635
rect 7113 2601 7147 2635
rect 8861 2601 8895 2635
rect 4905 2533 4939 2567
rect 7665 2533 7699 2567
rect 7941 2533 7975 2567
rect 8493 2533 8527 2567
rect 4261 2465 4295 2499
rect 5733 2465 5767 2499
rect 6285 2465 6319 2499
rect 9781 2465 9815 2499
rect 13461 2465 13495 2499
rect 14013 2465 14047 2499
rect 7849 2397 7883 2431
rect 5917 2329 5951 2363
rect 13645 2329 13679 2363
rect 3801 2261 3835 2295
rect 5181 2261 5215 2295
rect 9965 2261 9999 2295
rect 10425 2261 10459 2295
<< metal1 >>
rect 6638 39652 6644 39704
rect 6696 39692 6702 39704
rect 9306 39692 9312 39704
rect 6696 39664 9312 39692
rect 6696 39652 6702 39664
rect 9306 39652 9312 39664
rect 9364 39652 9370 39704
rect 9858 39652 9864 39704
rect 9916 39692 9922 39704
rect 13722 39692 13728 39704
rect 9916 39664 13728 39692
rect 9916 39652 9922 39664
rect 13722 39652 13728 39664
rect 13780 39652 13786 39704
rect 14 39584 20 39636
rect 72 39624 78 39636
rect 658 39624 664 39636
rect 72 39596 664 39624
rect 72 39584 78 39596
rect 658 39584 664 39596
rect 716 39584 722 39636
rect 1486 39584 1492 39636
rect 1544 39624 1550 39636
rect 2038 39624 2044 39636
rect 1544 39596 2044 39624
rect 1544 39584 1550 39596
rect 2038 39584 2044 39596
rect 2096 39584 2102 39636
rect 5626 39584 5632 39636
rect 5684 39624 5690 39636
rect 6454 39624 6460 39636
rect 5684 39596 6460 39624
rect 5684 39584 5690 39596
rect 6454 39584 6460 39596
rect 6512 39584 6518 39636
rect 7098 39584 7104 39636
rect 7156 39624 7162 39636
rect 7926 39624 7932 39636
rect 7156 39596 7932 39624
rect 7156 39584 7162 39596
rect 7926 39584 7932 39596
rect 7984 39584 7990 39636
rect 9766 39584 9772 39636
rect 9824 39624 9830 39636
rect 10778 39624 10784 39636
rect 9824 39596 10784 39624
rect 9824 39584 9830 39596
rect 10778 39584 10784 39596
rect 10836 39584 10842 39636
rect 13814 39584 13820 39636
rect 13872 39624 13878 39636
rect 15194 39624 15200 39636
rect 13872 39596 15200 39624
rect 13872 39584 13878 39596
rect 15194 39584 15200 39596
rect 15252 39584 15258 39636
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 2041 34731 2099 34737
rect 2041 34697 2053 34731
rect 2087 34728 2099 34731
rect 3142 34728 3148 34740
rect 2087 34700 3148 34728
rect 2087 34697 2099 34700
rect 2041 34691 2099 34697
rect 1578 34660 1584 34672
rect 1539 34632 1584 34660
rect 1578 34620 1584 34632
rect 1636 34620 1642 34672
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 2056 34524 2084 34691
rect 3142 34688 3148 34700
rect 3200 34688 3206 34740
rect 10873 34731 10931 34737
rect 10873 34697 10885 34731
rect 10919 34728 10931 34731
rect 11974 34728 11980 34740
rect 10919 34700 11980 34728
rect 10919 34697 10931 34700
rect 10873 34691 10931 34697
rect 11974 34688 11980 34700
rect 12032 34688 12038 34740
rect 8018 34552 8024 34604
rect 8076 34592 8082 34604
rect 8251 34595 8309 34601
rect 8251 34592 8263 34595
rect 8076 34564 8263 34592
rect 8076 34552 8082 34564
rect 8251 34561 8263 34564
rect 8297 34561 8309 34595
rect 8251 34555 8309 34561
rect 1443 34496 2084 34524
rect 8164 34527 8222 34533
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 8164 34493 8176 34527
rect 8210 34524 8222 34527
rect 8210 34496 8708 34524
rect 8210 34493 8222 34496
rect 8164 34487 8222 34493
rect 8680 34397 8708 34496
rect 9490 34484 9496 34536
rect 9548 34524 9554 34536
rect 10689 34527 10747 34533
rect 10689 34524 10701 34527
rect 9548 34496 10701 34524
rect 9548 34484 9554 34496
rect 10689 34493 10701 34496
rect 10735 34524 10747 34527
rect 11241 34527 11299 34533
rect 11241 34524 11253 34527
rect 10735 34496 11253 34524
rect 10735 34493 10747 34496
rect 10689 34487 10747 34493
rect 11241 34493 11253 34496
rect 11287 34493 11299 34527
rect 11241 34487 11299 34493
rect 8665 34391 8723 34397
rect 8665 34357 8677 34391
rect 8711 34388 8723 34391
rect 8846 34388 8852 34400
rect 8711 34360 8852 34388
rect 8711 34357 8723 34360
rect 8665 34351 8723 34357
rect 8846 34348 8852 34360
rect 8904 34348 8910 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 5350 29832 5356 29844
rect 5311 29804 5356 29832
rect 5350 29792 5356 29804
rect 5408 29792 5414 29844
rect 5166 29696 5172 29708
rect 5127 29668 5172 29696
rect 5166 29656 5172 29668
rect 5224 29656 5230 29708
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 4062 28976 4068 29028
rect 4120 29016 4126 29028
rect 5166 29016 5172 29028
rect 4120 28988 5172 29016
rect 4120 28976 4126 28988
rect 5166 28976 5172 28988
rect 5224 28976 5230 29028
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 13630 28744 13636 28756
rect 13591 28716 13636 28744
rect 13630 28704 13636 28716
rect 13688 28704 13694 28756
rect 13446 28608 13452 28620
rect 13407 28580 13452 28608
rect 13446 28568 13452 28580
rect 13504 28568 13510 28620
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 11330 27820 11336 27872
rect 11388 27860 11394 27872
rect 13446 27860 13452 27872
rect 11388 27832 13452 27860
rect 11388 27820 11394 27832
rect 13446 27820 13452 27832
rect 13504 27820 13510 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 4614 26568 4620 26580
rect 4575 26540 4620 26568
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 4430 26432 4436 26444
rect 4391 26404 4436 26432
rect 4430 26392 4436 26404
rect 4488 26392 4494 26444
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4430 25644 4436 25696
rect 4488 25684 4494 25696
rect 4525 25687 4583 25693
rect 4525 25684 4537 25687
rect 4488 25656 4537 25684
rect 4488 25644 4494 25656
rect 4525 25653 4537 25656
rect 4571 25684 4583 25687
rect 5994 25684 6000 25696
rect 4571 25656 6000 25684
rect 4571 25653 4583 25656
rect 4525 25647 4583 25653
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 106 22040 112 22092
rect 164 22080 170 22092
rect 1397 22083 1455 22089
rect 1397 22080 1409 22083
rect 164 22052 1409 22080
rect 164 22040 170 22052
rect 1397 22049 1409 22052
rect 1443 22080 1455 22083
rect 1578 22080 1584 22092
rect 1443 22052 1584 22080
rect 1443 22049 1455 22052
rect 1397 22043 1455 22049
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 106 21836 112 21888
rect 164 21876 170 21888
rect 1581 21879 1639 21885
rect 1581 21876 1593 21879
rect 164 21848 1593 21876
rect 164 21836 170 21848
rect 1581 21845 1593 21848
rect 1627 21845 1639 21879
rect 1581 21839 1639 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 6340 19907 6398 19913
rect 6340 19873 6352 19907
rect 6386 19904 6398 19907
rect 6638 19904 6644 19916
rect 6386 19876 6644 19904
rect 6386 19873 6398 19876
rect 6340 19867 6398 19873
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6411 19703 6469 19709
rect 6411 19669 6423 19703
rect 6457 19700 6469 19703
rect 6730 19700 6736 19712
rect 6457 19672 6736 19700
rect 6457 19669 6469 19672
rect 6411 19663 6469 19669
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 6914 19700 6920 19712
rect 6875 19672 6920 19700
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 5258 19496 5264 19508
rect 5219 19468 5264 19496
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 6365 19499 6423 19505
rect 6365 19465 6377 19499
rect 6411 19496 6423 19499
rect 6638 19496 6644 19508
rect 6411 19468 6644 19496
rect 6411 19465 6423 19468
rect 6365 19459 6423 19465
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5166 19292 5172 19304
rect 5123 19264 5172 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 1394 19184 1400 19236
rect 1452 19224 1458 19236
rect 6380 19224 6408 19459
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 7064 19332 7205 19360
rect 7064 19320 7070 19332
rect 7193 19329 7205 19332
rect 7239 19329 7251 19363
rect 7193 19323 7251 19329
rect 6914 19224 6920 19236
rect 1452 19196 6408 19224
rect 6875 19196 6920 19224
rect 1452 19184 1458 19196
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 7009 19227 7067 19233
rect 7009 19193 7021 19227
rect 7055 19193 7067 19227
rect 7009 19187 7067 19193
rect 5166 19116 5172 19168
rect 5224 19156 5230 19168
rect 5629 19159 5687 19165
rect 5629 19156 5641 19159
rect 5224 19128 5641 19156
rect 5224 19116 5230 19128
rect 5629 19125 5641 19128
rect 5675 19125 5687 19159
rect 5629 19119 5687 19125
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7024 19156 7052 19187
rect 6880 19128 7052 19156
rect 6880 19116 6886 19128
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 9861 18955 9919 18961
rect 9861 18952 9873 18955
rect 9824 18924 9873 18952
rect 9824 18912 9830 18924
rect 9861 18921 9873 18924
rect 9907 18921 9919 18955
rect 9861 18915 9919 18921
rect 5997 18887 6055 18893
rect 5997 18853 6009 18887
rect 6043 18884 6055 18887
rect 6086 18884 6092 18896
rect 6043 18856 6092 18884
rect 6043 18853 6055 18856
rect 5997 18847 6055 18853
rect 6086 18844 6092 18856
rect 6144 18884 6150 18896
rect 6822 18884 6828 18896
rect 6144 18856 6828 18884
rect 6144 18844 6150 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 7561 18887 7619 18893
rect 7561 18884 7573 18887
rect 7524 18856 7573 18884
rect 7524 18844 7530 18856
rect 7561 18853 7573 18856
rect 7607 18853 7619 18887
rect 7561 18847 7619 18853
rect 4868 18819 4926 18825
rect 4868 18785 4880 18819
rect 4914 18816 4926 18819
rect 5166 18816 5172 18828
rect 4914 18788 5172 18816
rect 4914 18785 4926 18788
rect 4868 18779 4926 18785
rect 5166 18776 5172 18788
rect 5224 18776 5230 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18717 5963 18751
rect 6178 18748 6184 18760
rect 6139 18720 6184 18748
rect 5905 18711 5963 18717
rect 5920 18680 5948 18711
rect 6178 18708 6184 18720
rect 6236 18708 6242 18760
rect 7006 18708 7012 18760
rect 7064 18748 7070 18760
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 7064 18720 7481 18748
rect 7064 18708 7070 18720
rect 7469 18717 7481 18720
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 6638 18680 6644 18692
rect 5920 18652 6644 18680
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 8018 18680 8024 18692
rect 7979 18652 8024 18680
rect 8018 18640 8024 18652
rect 8076 18640 8082 18692
rect 4939 18615 4997 18621
rect 4939 18581 4951 18615
rect 4985 18612 4997 18615
rect 5074 18612 5080 18624
rect 4985 18584 5080 18612
rect 4985 18581 4997 18584
rect 4939 18575 4997 18581
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 5350 18612 5356 18624
rect 5311 18584 5356 18612
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 5718 18612 5724 18624
rect 5679 18584 5724 18612
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 4295 18411 4353 18417
rect 4295 18377 4307 18411
rect 4341 18408 4353 18411
rect 6914 18408 6920 18420
rect 4341 18380 6920 18408
rect 4341 18377 4353 18380
rect 4295 18371 4353 18377
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 9306 18408 9312 18420
rect 9267 18380 9312 18408
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 4709 18343 4767 18349
rect 4709 18309 4721 18343
rect 4755 18340 4767 18343
rect 7834 18340 7840 18352
rect 4755 18312 7840 18340
rect 4755 18309 4767 18312
rect 4709 18303 4767 18309
rect 4224 18207 4282 18213
rect 4224 18173 4236 18207
rect 4270 18204 4282 18207
rect 4724 18204 4752 18303
rect 7834 18300 7840 18312
rect 7892 18300 7898 18352
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18272 5319 18275
rect 5718 18272 5724 18284
rect 5307 18244 5724 18272
rect 5307 18241 5319 18244
rect 5261 18235 5319 18241
rect 5718 18232 5724 18244
rect 5776 18272 5782 18284
rect 6822 18272 6828 18284
rect 5776 18244 6828 18272
rect 5776 18232 5782 18244
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 8018 18272 8024 18284
rect 7979 18244 8024 18272
rect 8018 18232 8024 18244
rect 8076 18272 8082 18284
rect 8941 18275 8999 18281
rect 8941 18272 8953 18275
rect 8076 18244 8953 18272
rect 8076 18232 8082 18244
rect 8941 18241 8953 18244
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 4270 18176 4752 18204
rect 8956 18204 8984 18235
rect 9160 18207 9218 18213
rect 9160 18204 9172 18207
rect 8956 18176 9172 18204
rect 4270 18173 4282 18176
rect 4224 18167 4282 18173
rect 9160 18173 9172 18176
rect 9206 18204 9218 18207
rect 9306 18204 9312 18216
rect 9206 18176 9312 18204
rect 9206 18173 9218 18176
rect 9160 18167 9218 18173
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 5350 18096 5356 18148
rect 5408 18136 5414 18148
rect 5902 18136 5908 18148
rect 5408 18108 5453 18136
rect 5863 18108 5908 18136
rect 5408 18096 5414 18108
rect 5902 18096 5908 18108
rect 5960 18136 5966 18148
rect 7006 18136 7012 18148
rect 5960 18108 7012 18136
rect 5960 18096 5966 18108
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 7653 18139 7711 18145
rect 7653 18105 7665 18139
rect 7699 18105 7711 18139
rect 7653 18099 7711 18105
rect 5077 18071 5135 18077
rect 5077 18037 5089 18071
rect 5123 18068 5135 18071
rect 5166 18068 5172 18080
rect 5123 18040 5172 18068
rect 5123 18037 5135 18040
rect 5077 18031 5135 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 6086 18028 6092 18080
rect 6144 18068 6150 18080
rect 6181 18071 6239 18077
rect 6181 18068 6193 18071
rect 6144 18040 6193 18068
rect 6144 18028 6150 18040
rect 6181 18037 6193 18040
rect 6227 18037 6239 18071
rect 6638 18068 6644 18080
rect 6599 18040 6644 18068
rect 6181 18031 6239 18037
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7558 18028 7564 18080
rect 7616 18068 7622 18080
rect 7668 18068 7696 18099
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 7800 18108 7845 18136
rect 7800 18096 7806 18108
rect 7616 18040 7696 18068
rect 7616 18028 7622 18040
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 9674 18068 9680 18080
rect 7892 18040 9680 18068
rect 7892 18028 7898 18040
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 5074 17824 5080 17876
rect 5132 17864 5138 17876
rect 5997 17867 6055 17873
rect 5997 17864 6009 17867
rect 5132 17836 6009 17864
rect 5132 17824 5138 17836
rect 5997 17833 6009 17836
rect 6043 17833 6055 17867
rect 5997 17827 6055 17833
rect 6822 17824 6828 17876
rect 6880 17864 6886 17876
rect 9815 17867 9873 17873
rect 9815 17864 9827 17867
rect 6880 17836 9827 17864
rect 6880 17824 6886 17836
rect 9815 17833 9827 17836
rect 9861 17833 9873 17867
rect 9815 17827 9873 17833
rect 5169 17799 5227 17805
rect 5169 17765 5181 17799
rect 5215 17796 5227 17799
rect 5258 17796 5264 17808
rect 5215 17768 5264 17796
rect 5215 17765 5227 17768
rect 5169 17759 5227 17765
rect 5258 17756 5264 17768
rect 5316 17756 5322 17808
rect 5350 17756 5356 17808
rect 5408 17796 5414 17808
rect 6733 17799 6791 17805
rect 6733 17796 6745 17799
rect 5408 17768 6745 17796
rect 5408 17756 5414 17768
rect 6733 17765 6745 17768
rect 6779 17765 6791 17799
rect 6733 17759 6791 17765
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 2958 17728 2964 17740
rect 2922 17700 2964 17728
rect 2958 17688 2964 17700
rect 3016 17737 3022 17740
rect 3016 17731 3070 17737
rect 3016 17697 3024 17731
rect 3058 17728 3070 17731
rect 3510 17728 3516 17740
rect 3058 17700 3516 17728
rect 3058 17697 3070 17700
rect 3016 17691 3070 17697
rect 3016 17688 3022 17691
rect 3510 17688 3516 17700
rect 3568 17728 3574 17740
rect 4062 17728 4068 17740
rect 3568 17700 4068 17728
rect 3568 17688 3574 17700
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 9585 17731 9643 17737
rect 9585 17697 9597 17731
rect 9631 17728 9643 17731
rect 9674 17728 9680 17740
rect 9631 17700 9680 17728
rect 9631 17697 9643 17700
rect 9585 17691 9643 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 11422 17728 11428 17740
rect 11383 17700 11428 17728
rect 11422 17688 11428 17700
rect 11480 17688 11486 17740
rect 3099 17663 3157 17669
rect 3099 17629 3111 17663
rect 3145 17660 3157 17663
rect 4798 17660 4804 17672
rect 3145 17632 4804 17660
rect 3145 17629 3157 17632
rect 3099 17623 3157 17629
rect 4798 17620 4804 17632
rect 4856 17660 4862 17672
rect 5077 17663 5135 17669
rect 5077 17660 5089 17663
rect 4856 17632 5089 17660
rect 4856 17620 4862 17632
rect 5077 17629 5089 17632
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 6641 17663 6699 17669
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 6730 17660 6736 17672
rect 6687 17632 6736 17660
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17660 6975 17663
rect 7558 17660 7564 17672
rect 6963 17632 7564 17660
rect 6963 17629 6975 17632
rect 6917 17623 6975 17629
rect 1578 17592 1584 17604
rect 1539 17564 1584 17592
rect 1578 17552 1584 17564
rect 1636 17552 1642 17604
rect 5629 17595 5687 17601
rect 5629 17561 5641 17595
rect 5675 17592 5687 17595
rect 6178 17592 6184 17604
rect 5675 17564 6184 17592
rect 5675 17561 5687 17564
rect 5629 17555 5687 17561
rect 6178 17552 6184 17564
rect 6236 17592 6242 17604
rect 6932 17592 6960 17623
rect 7558 17620 7564 17632
rect 7616 17660 7622 17672
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7616 17632 7941 17660
rect 7616 17620 7622 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 8110 17660 8116 17672
rect 8071 17632 8116 17660
rect 7929 17623 7987 17629
rect 8110 17620 8116 17632
rect 8168 17620 8174 17672
rect 6236 17564 6960 17592
rect 6236 17552 6242 17564
rect 7650 17524 7656 17536
rect 7611 17496 7656 17524
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 11609 17527 11667 17533
rect 11609 17493 11621 17527
rect 11655 17524 11667 17527
rect 11974 17524 11980 17536
rect 11655 17496 11980 17524
rect 11655 17493 11667 17496
rect 11609 17487 11667 17493
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1452 17292 1593 17320
rect 1452 17280 1458 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 2958 17320 2964 17332
rect 2919 17292 2964 17320
rect 1581 17283 1639 17289
rect 2958 17280 2964 17292
rect 3016 17280 3022 17332
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 6178 17320 6184 17332
rect 5408 17292 6184 17320
rect 5408 17280 5414 17292
rect 6178 17280 6184 17292
rect 6236 17280 6242 17332
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 7745 17323 7803 17329
rect 7745 17320 7757 17323
rect 7524 17292 7757 17320
rect 7524 17280 7530 17292
rect 7745 17289 7757 17292
rect 7791 17289 7803 17323
rect 7745 17283 7803 17289
rect 8110 17280 8116 17332
rect 8168 17320 8174 17332
rect 8389 17323 8447 17329
rect 8389 17320 8401 17323
rect 8168 17292 8401 17320
rect 8168 17280 8174 17292
rect 8389 17289 8401 17292
rect 8435 17289 8447 17323
rect 11422 17320 11428 17332
rect 11383 17292 11428 17320
rect 8389 17283 8447 17289
rect 4295 17255 4353 17261
rect 4295 17221 4307 17255
rect 4341 17252 4353 17255
rect 6638 17252 6644 17264
rect 4341 17224 6644 17252
rect 4341 17221 4353 17224
rect 4295 17215 4353 17221
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 6730 17212 6736 17264
rect 6788 17252 6794 17264
rect 8021 17255 8079 17261
rect 8021 17252 8033 17255
rect 6788 17224 8033 17252
rect 6788 17212 6794 17224
rect 8021 17221 8033 17224
rect 8067 17221 8079 17255
rect 8021 17215 8079 17221
rect 5074 17144 5080 17196
rect 5132 17184 5138 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 5132 17156 5273 17184
rect 5132 17144 5138 17156
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 5902 17184 5908 17196
rect 5863 17156 5908 17184
rect 5261 17147 5319 17153
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 8404 17184 8432 17283
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8404 17156 8677 17184
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 9306 17184 9312 17196
rect 9267 17156 9312 17184
rect 8665 17147 8723 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 4224 17119 4282 17125
rect 4224 17085 4236 17119
rect 4270 17116 4282 17119
rect 6822 17116 6828 17128
rect 4270 17088 4752 17116
rect 6783 17088 6828 17116
rect 4270 17085 4282 17088
rect 4224 17079 4282 17085
rect 4724 16989 4752 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 5077 17051 5135 17057
rect 5077 17017 5089 17051
rect 5123 17048 5135 17051
rect 5258 17048 5264 17060
rect 5123 17020 5264 17048
rect 5123 17017 5135 17020
rect 5077 17011 5135 17017
rect 5258 17008 5264 17020
rect 5316 17048 5322 17060
rect 5353 17051 5411 17057
rect 5353 17048 5365 17051
rect 5316 17020 5365 17048
rect 5316 17008 5322 17020
rect 5353 17017 5365 17020
rect 5399 17017 5411 17051
rect 8754 17048 8760 17060
rect 8715 17020 8760 17048
rect 5353 17011 5411 17017
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 4709 16983 4767 16989
rect 4709 16949 4721 16983
rect 4755 16980 4767 16983
rect 5626 16980 5632 16992
rect 4755 16952 5632 16980
rect 4755 16949 4767 16952
rect 4709 16943 4767 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 6641 16983 6699 16989
rect 6641 16949 6653 16983
rect 6687 16980 6699 16983
rect 7190 16980 7196 16992
rect 6687 16952 7196 16980
rect 6687 16949 6699 16952
rect 6641 16943 6699 16949
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 9674 16980 9680 16992
rect 9635 16952 9680 16980
rect 9674 16940 9680 16952
rect 9732 16980 9738 16992
rect 10870 16980 10876 16992
rect 9732 16952 10876 16980
rect 9732 16940 9738 16952
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 4798 16776 4804 16788
rect 4759 16748 4804 16776
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 6236 16748 6285 16776
rect 6236 16736 6242 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 7708 16748 8033 16776
rect 7708 16736 7714 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 5534 16668 5540 16720
rect 5592 16708 5598 16720
rect 5674 16711 5732 16717
rect 5674 16708 5686 16711
rect 5592 16680 5686 16708
rect 5592 16668 5598 16680
rect 5674 16677 5686 16680
rect 5720 16677 5732 16711
rect 5674 16671 5732 16677
rect 7190 16668 7196 16720
rect 7248 16708 7254 16720
rect 7422 16711 7480 16717
rect 7422 16708 7434 16711
rect 7248 16680 7434 16708
rect 7248 16668 7254 16680
rect 7422 16677 7434 16680
rect 7468 16677 7480 16711
rect 7422 16671 7480 16677
rect 5166 16600 5172 16652
rect 5224 16640 5230 16652
rect 10594 16640 10600 16652
rect 5224 16612 10600 16640
rect 5224 16600 5230 16612
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 5353 16575 5411 16581
rect 5353 16572 5365 16575
rect 4580 16544 5365 16572
rect 4580 16532 4586 16544
rect 5353 16541 5365 16544
rect 5399 16541 5411 16575
rect 5353 16535 5411 16541
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6696 16544 7113 16572
rect 6696 16532 6702 16544
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 5258 16436 5264 16448
rect 5219 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 8573 16439 8631 16445
rect 8573 16436 8585 16439
rect 8260 16408 8585 16436
rect 8260 16396 8266 16408
rect 8573 16405 8585 16408
rect 8619 16436 8631 16439
rect 8754 16436 8760 16448
rect 8619 16408 8760 16436
rect 8619 16405 8631 16408
rect 8573 16399 8631 16405
rect 8754 16396 8760 16408
rect 8812 16396 8818 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 6086 16232 6092 16244
rect 5951 16204 6092 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 8202 16232 8208 16244
rect 8163 16204 8208 16232
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 6086 16096 6092 16108
rect 5684 16068 6092 16096
rect 5684 16056 5690 16068
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 4706 15988 4712 16040
rect 4764 16028 4770 16040
rect 4985 16031 5043 16037
rect 4985 16028 4997 16031
rect 4764 16000 4997 16028
rect 4764 15988 4770 16000
rect 4985 15997 4997 16000
rect 5031 15997 5043 16031
rect 4985 15991 5043 15997
rect 7285 16031 7343 16037
rect 7285 15997 7297 16031
rect 7331 16028 7343 16031
rect 7466 16028 7472 16040
rect 7331 16000 7472 16028
rect 7331 15997 7343 16000
rect 7285 15991 7343 15997
rect 7466 15988 7472 16000
rect 7524 15988 7530 16040
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15960 4951 15963
rect 5347 15963 5405 15969
rect 5347 15960 5359 15963
rect 4939 15932 5359 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 5347 15929 5359 15932
rect 5393 15960 5405 15963
rect 5534 15960 5540 15972
rect 5393 15932 5540 15960
rect 5393 15929 5405 15932
rect 5347 15923 5405 15929
rect 5534 15920 5540 15932
rect 5592 15960 5598 15972
rect 6273 15963 6331 15969
rect 6273 15960 6285 15963
rect 5592 15932 6285 15960
rect 5592 15920 5598 15932
rect 6273 15929 6285 15932
rect 6319 15960 6331 15963
rect 7606 15963 7664 15969
rect 6319 15932 7236 15960
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 7208 15904 7236 15932
rect 7606 15929 7618 15963
rect 7652 15929 7664 15963
rect 7606 15923 7664 15929
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 6638 15892 6644 15904
rect 6599 15864 6644 15892
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15892 7254 15904
rect 7621 15892 7649 15923
rect 7248 15864 7649 15892
rect 7248 15852 7254 15864
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 6365 15691 6423 15697
rect 6365 15688 6377 15691
rect 5316 15660 6377 15688
rect 5316 15648 5322 15660
rect 6365 15657 6377 15660
rect 6411 15657 6423 15691
rect 6365 15651 6423 15657
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 5766 15623 5824 15629
rect 5766 15620 5778 15623
rect 5592 15592 5778 15620
rect 5592 15580 5598 15592
rect 5766 15589 5778 15592
rect 5812 15589 5824 15623
rect 5766 15583 5824 15589
rect 5445 15487 5503 15493
rect 5445 15453 5457 15487
rect 5491 15484 5503 15487
rect 5902 15484 5908 15496
rect 5491 15456 5908 15484
rect 5491 15453 5503 15456
rect 5445 15447 5503 15453
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 8294 15484 8300 15496
rect 8255 15456 8300 15484
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 4985 15351 5043 15357
rect 4985 15348 4997 15351
rect 4764 15320 4997 15348
rect 4764 15308 4770 15320
rect 4985 15317 4997 15320
rect 5031 15317 5043 15351
rect 7190 15348 7196 15360
rect 7151 15320 7196 15348
rect 4985 15311 5043 15317
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 7466 15348 7472 15360
rect 7427 15320 7472 15348
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 8312 15008 8340 15104
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8312 14980 8585 15008
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 8846 15008 8852 15020
rect 8807 14980 8852 15008
rect 8573 14971 8631 14977
rect 8846 14968 8852 14980
rect 8904 14968 8910 15020
rect 8021 14875 8079 14881
rect 8021 14841 8033 14875
rect 8067 14872 8079 14875
rect 8662 14872 8668 14884
rect 8067 14844 8668 14872
rect 8067 14841 8079 14844
rect 8021 14835 8079 14841
rect 8662 14832 8668 14844
rect 8720 14832 8726 14884
rect 5902 14804 5908 14816
rect 5815 14776 5908 14804
rect 5902 14764 5908 14776
rect 5960 14804 5966 14816
rect 6914 14804 6920 14816
rect 5960 14776 6920 14804
rect 5960 14764 5966 14776
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 8662 14600 8668 14612
rect 8623 14572 8668 14600
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 13630 14600 13636 14612
rect 13591 14572 13636 14600
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 7190 14492 7196 14544
rect 7248 14532 7254 14544
rect 8107 14535 8165 14541
rect 8107 14532 8119 14535
rect 7248 14504 8119 14532
rect 7248 14492 7254 14504
rect 8107 14501 8119 14504
rect 8153 14501 8165 14535
rect 8107 14495 8165 14501
rect 8122 14464 8150 14495
rect 9766 14492 9772 14544
rect 9824 14532 9830 14544
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9824 14504 9873 14532
rect 9824 14492 9830 14504
rect 9861 14501 9873 14504
rect 9907 14501 9919 14535
rect 9861 14495 9919 14501
rect 8662 14464 8668 14476
rect 8122 14436 8668 14464
rect 8662 14424 8668 14436
rect 8720 14424 8726 14476
rect 13446 14464 13452 14476
rect 13407 14436 13452 14464
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14396 7803 14399
rect 8202 14396 8208 14408
rect 7791 14368 8208 14396
rect 7791 14365 7803 14368
rect 7745 14359 7803 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 11238 14396 11244 14408
rect 9815 14368 11244 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 8846 14288 8852 14340
rect 8904 14328 8910 14340
rect 10321 14331 10379 14337
rect 10321 14328 10333 14331
rect 8904 14300 10333 14328
rect 8904 14288 8910 14300
rect 10321 14297 10333 14300
rect 10367 14328 10379 14331
rect 12158 14328 12164 14340
rect 10367 14300 12164 14328
rect 10367 14297 10379 14300
rect 10321 14291 10379 14297
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7006 14260 7012 14272
rect 6963 14232 7012 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7285 14263 7343 14269
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 8018 14260 8024 14272
rect 7331 14232 8024 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 11238 14056 11244 14068
rect 11199 14028 11244 14056
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 8202 13988 8208 14000
rect 8163 13960 8208 13988
rect 8202 13948 8208 13960
rect 8260 13988 8266 14000
rect 8941 13991 8999 13997
rect 8941 13988 8953 13991
rect 8260 13960 8953 13988
rect 8260 13948 8266 13960
rect 8941 13957 8953 13960
rect 8987 13957 8999 13991
rect 8941 13951 8999 13957
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10008 13960 11008 13988
rect 10008 13948 10014 13960
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10042 13920 10048 13932
rect 9815 13892 10048 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10226 13920 10232 13932
rect 10187 13892 10232 13920
rect 10226 13880 10232 13892
rect 10284 13880 10290 13932
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6178 13716 6184 13728
rect 6139 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6840 13716 6868 13815
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 7282 13852 7288 13864
rect 7064 13824 7288 13852
rect 7064 13812 7070 13824
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7708 13824 7757 13852
rect 7708 13812 7714 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 8018 13852 8024 13864
rect 7979 13824 8024 13852
rect 7745 13815 7803 13821
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 9950 13784 9956 13796
rect 9911 13756 9956 13784
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10042 13744 10048 13796
rect 10100 13784 10106 13796
rect 10100 13756 10145 13784
rect 10100 13744 10106 13756
rect 7006 13716 7012 13728
rect 6687 13688 7012 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 8662 13716 8668 13728
rect 8623 13688 8668 13716
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 9398 13716 9404 13728
rect 9359 13688 9404 13716
rect 9398 13676 9404 13688
rect 9456 13716 9462 13728
rect 9674 13716 9680 13728
rect 9456 13688 9680 13716
rect 9456 13676 9462 13688
rect 9674 13676 9680 13688
rect 9732 13676 9738 13728
rect 10980 13725 11008 13960
rect 11054 13744 11060 13796
rect 11112 13784 11118 13796
rect 13446 13784 13452 13796
rect 11112 13756 13452 13784
rect 11112 13744 11118 13756
rect 13446 13744 13452 13756
rect 13504 13744 13510 13796
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 12250 13716 12256 13728
rect 11011 13688 12256 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 12250 13676 12256 13688
rect 12308 13676 12314 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 14 13472 20 13524
rect 72 13512 78 13524
rect 10042 13512 10048 13524
rect 72 13484 4154 13512
rect 10003 13484 10048 13512
rect 72 13472 78 13484
rect 4126 13376 4154 13484
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10597 13515 10655 13521
rect 10597 13481 10609 13515
rect 10643 13512 10655 13515
rect 10643 13484 11652 13512
rect 10643 13481 10655 13484
rect 10597 13475 10655 13481
rect 6178 13404 6184 13456
rect 6236 13444 6242 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 6236 13416 6285 13444
rect 6236 13404 6242 13416
rect 6273 13413 6285 13416
rect 6319 13444 6331 13447
rect 7650 13444 7656 13456
rect 6319 13416 7656 13444
rect 6319 13413 6331 13416
rect 6273 13407 6331 13413
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 11624 13453 11652 13484
rect 11609 13447 11667 13453
rect 11609 13413 11621 13447
rect 11655 13444 11667 13447
rect 11698 13444 11704 13456
rect 11655 13416 11704 13444
rect 11655 13413 11667 13416
rect 11609 13407 11667 13413
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 12158 13444 12164 13456
rect 12119 13416 12164 13444
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4126 13348 4537 13376
rect 4525 13345 4537 13348
rect 4571 13376 4583 13379
rect 5166 13376 5172 13388
rect 4571 13348 5172 13376
rect 4571 13345 4583 13348
rect 4525 13339 4583 13345
rect 5166 13336 5172 13348
rect 5224 13376 5230 13388
rect 5261 13379 5319 13385
rect 5261 13376 5273 13379
rect 5224 13348 5273 13376
rect 5224 13336 5230 13348
rect 5261 13345 5273 13348
rect 5307 13345 5319 13379
rect 7006 13376 7012 13388
rect 6967 13348 7012 13376
rect 5261 13339 5319 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 7282 13376 7288 13388
rect 7239 13348 7288 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 7208 13308 7236 13339
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 7558 13376 7564 13388
rect 7519 13348 7564 13376
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7926 13376 7932 13388
rect 7887 13348 7932 13376
rect 7926 13336 7932 13348
rect 7984 13336 7990 13388
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 10284 13348 10824 13376
rect 10284 13336 10290 13348
rect 5951 13280 7236 13308
rect 8205 13311 8263 13317
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6656 13181 6684 13280
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 8251 13280 9689 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 9677 13277 9689 13280
rect 9723 13308 9735 13311
rect 10686 13308 10692 13320
rect 9723 13280 10692 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10796 13308 10824 13348
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 10796 13280 11529 13308
rect 11517 13277 11529 13280
rect 11563 13308 11575 13311
rect 12158 13308 12164 13320
rect 11563 13280 12164 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 6641 13175 6699 13181
rect 6641 13141 6653 13175
rect 6687 13172 6699 13175
rect 6730 13172 6736 13184
rect 6687 13144 6736 13172
rect 6687 13141 6699 13144
rect 6641 13135 6699 13141
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8076 13144 8493 13172
rect 8076 13132 8082 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 9306 13172 9312 13184
rect 9263 13144 9312 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 10686 12968 10692 12980
rect 10647 12940 10692 12968
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11698 12968 11704 12980
rect 11659 12940 11704 12968
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12250 12928 12256 12980
rect 12308 12968 12314 12980
rect 12575 12971 12633 12977
rect 12575 12968 12587 12971
rect 12308 12940 12587 12968
rect 12308 12928 12314 12940
rect 12575 12937 12587 12940
rect 12621 12937 12633 12971
rect 12575 12931 12633 12937
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12832 4031 12835
rect 4154 12832 4160 12844
rect 4019 12804 4160 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 4154 12792 4160 12804
rect 4212 12792 4218 12844
rect 5074 12792 5080 12844
rect 5132 12832 5138 12844
rect 8386 12832 8392 12844
rect 5132 12804 8392 12832
rect 5132 12792 5138 12804
rect 8386 12792 8392 12804
rect 8444 12832 8450 12844
rect 11054 12832 11060 12844
rect 8444 12804 11060 12832
rect 8444 12792 8450 12804
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11425 12835 11483 12841
rect 11425 12801 11437 12835
rect 11471 12832 11483 12835
rect 13722 12832 13728 12844
rect 11471 12804 13728 12832
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 4614 12764 4620 12776
rect 4575 12736 4620 12764
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5166 12764 5172 12776
rect 5127 12736 5172 12764
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12733 5319 12767
rect 5626 12764 5632 12776
rect 5587 12736 5632 12764
rect 5261 12727 5319 12733
rect 5276 12696 5304 12727
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6564 12736 6837 12764
rect 4356 12668 5304 12696
rect 4356 12640 4384 12668
rect 4338 12628 4344 12640
rect 4299 12600 4344 12628
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 4706 12628 4712 12640
rect 4667 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 6178 12588 6184 12600
rect 6236 12628 6242 12640
rect 6564 12637 6592 12736
rect 6825 12733 6837 12736
rect 6871 12764 6883 12767
rect 7006 12764 7012 12776
rect 6871 12736 7012 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7650 12764 7656 12776
rect 7611 12736 7656 12764
rect 7285 12727 7343 12733
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 7300 12696 7328 12727
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 8018 12764 8024 12776
rect 7979 12736 8024 12764
rect 8018 12724 8024 12736
rect 8076 12724 8082 12776
rect 9125 12767 9183 12773
rect 9125 12733 9137 12767
rect 9171 12764 9183 12767
rect 9306 12764 9312 12776
rect 9171 12736 9312 12764
rect 9171 12733 9183 12736
rect 9125 12727 9183 12733
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 10778 12764 10784 12776
rect 10091 12736 10784 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 10940 12767 10998 12773
rect 10940 12733 10952 12767
rect 10986 12764 10998 12767
rect 11440 12764 11468 12795
rect 13722 12792 13728 12804
rect 13780 12832 13786 12844
rect 14734 12832 14740 12844
rect 13780 12804 14740 12832
rect 13780 12792 13786 12804
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 10986 12736 11468 12764
rect 10986 12733 10998 12736
rect 10940 12727 10998 12733
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12472 12767 12530 12773
rect 12472 12764 12484 12767
rect 12124 12736 12484 12764
rect 12124 12724 12130 12736
rect 12472 12733 12484 12736
rect 12518 12764 12530 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12518 12736 12909 12764
rect 12518 12733 12530 12736
rect 12472 12727 12530 12733
rect 12897 12733 12909 12736
rect 12943 12764 12955 12767
rect 13446 12764 13452 12776
rect 12943 12736 13452 12764
rect 12943 12733 12955 12736
rect 12897 12727 12955 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 8573 12699 8631 12705
rect 8573 12696 8585 12699
rect 6788 12668 8585 12696
rect 6788 12656 6794 12668
rect 8573 12665 8585 12668
rect 8619 12665 8631 12699
rect 8573 12659 8631 12665
rect 9487 12699 9545 12705
rect 9487 12665 9499 12699
rect 9533 12665 9545 12699
rect 9487 12659 9545 12665
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6236 12600 6561 12628
rect 6236 12588 6242 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 7466 12628 7472 12640
rect 7147 12600 7472 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 9033 12631 9091 12637
rect 9033 12628 9045 12631
rect 8720 12600 9045 12628
rect 8720 12588 8726 12600
rect 9033 12597 9045 12600
rect 9079 12628 9091 12631
rect 9508 12628 9536 12659
rect 10042 12628 10048 12640
rect 9079 12600 10048 12628
rect 9079 12597 9091 12600
rect 9033 12591 9091 12597
rect 10042 12588 10048 12600
rect 10100 12628 10106 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 10100 12600 10333 12628
rect 10100 12588 10106 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10321 12591 10379 12597
rect 11011 12631 11069 12637
rect 11011 12597 11023 12631
rect 11057 12628 11069 12631
rect 11238 12628 11244 12640
rect 11057 12600 11244 12628
rect 11057 12597 11069 12600
rect 11011 12591 11069 12597
rect 11238 12588 11244 12600
rect 11296 12588 11302 12640
rect 12158 12628 12164 12640
rect 12119 12600 12164 12628
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 6457 12427 6515 12433
rect 6457 12393 6469 12427
rect 6503 12424 6515 12427
rect 6638 12424 6644 12436
rect 6503 12396 6644 12424
rect 6503 12393 6515 12396
rect 6457 12387 6515 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 7708 12396 9137 12424
rect 7708 12384 7714 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 7558 12356 7564 12368
rect 7116 12328 7564 12356
rect 5166 12288 5172 12300
rect 5079 12260 5172 12288
rect 5166 12248 5172 12260
rect 5224 12288 5230 12300
rect 5718 12288 5724 12300
rect 5224 12260 5724 12288
rect 5224 12248 5230 12260
rect 5718 12248 5724 12260
rect 5776 12248 5782 12300
rect 6089 12291 6147 12297
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6178 12288 6184 12300
rect 6135 12260 6184 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 6178 12248 6184 12260
rect 6236 12288 6242 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6236 12260 6469 12288
rect 6236 12248 6242 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6638 12288 6644 12300
rect 6599 12260 6644 12288
rect 6457 12251 6515 12257
rect 6472 12220 6500 12251
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 7116 12297 7144 12328
rect 7558 12316 7564 12328
rect 7616 12356 7622 12368
rect 8294 12356 8300 12368
rect 7616 12328 8300 12356
rect 7616 12316 7622 12328
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 9140 12356 9168 12387
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 9456 12396 10609 12424
rect 9456 12384 9462 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 13630 12424 13636 12436
rect 10836 12396 11652 12424
rect 13591 12396 13636 12424
rect 10836 12384 10842 12396
rect 11624 12368 11652 12396
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 9490 12356 9496 12368
rect 9140 12328 9496 12356
rect 9490 12316 9496 12328
rect 9548 12316 9554 12368
rect 9930 12359 9988 12365
rect 9930 12325 9942 12359
rect 9976 12356 9988 12359
rect 10042 12356 10048 12368
rect 9976 12328 10048 12356
rect 9976 12325 9988 12328
rect 9930 12319 9988 12325
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 11238 12316 11244 12368
rect 11296 12356 11302 12368
rect 11517 12359 11575 12365
rect 11517 12356 11529 12359
rect 11296 12328 11529 12356
rect 11296 12316 11302 12328
rect 11517 12325 11529 12328
rect 11563 12325 11575 12359
rect 11517 12319 11575 12325
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 11664 12328 11757 12356
rect 11664 12316 11670 12328
rect 7101 12291 7159 12297
rect 7101 12257 7113 12291
rect 7147 12257 7159 12291
rect 7101 12251 7159 12257
rect 7377 12291 7435 12297
rect 7377 12257 7389 12291
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 7190 12220 7196 12232
rect 6472 12192 7196 12220
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4212 12124 4997 12152
rect 4212 12112 4218 12124
rect 4985 12121 4997 12124
rect 5031 12152 5043 12155
rect 5626 12152 5632 12164
rect 5031 12124 5632 12152
rect 5031 12121 5043 12124
rect 4985 12115 5043 12121
rect 5626 12112 5632 12124
rect 5684 12152 5690 12164
rect 7006 12152 7012 12164
rect 5684 12124 7012 12152
rect 5684 12112 5690 12124
rect 7006 12112 7012 12124
rect 7064 12152 7070 12164
rect 7392 12152 7420 12251
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 8608 12291 8666 12297
rect 8608 12288 8620 12291
rect 8444 12260 8620 12288
rect 8444 12248 8450 12260
rect 8608 12257 8620 12260
rect 8654 12257 8666 12291
rect 13446 12288 13452 12300
rect 13407 12260 13452 12288
rect 8608 12251 8666 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12220 9735 12223
rect 10778 12220 10784 12232
rect 9723 12192 10784 12220
rect 9723 12189 9735 12192
rect 9677 12183 9735 12189
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 7064 12124 7420 12152
rect 8711 12155 8769 12161
rect 7064 12112 7070 12124
rect 8711 12121 8723 12155
rect 8757 12152 8769 12155
rect 9766 12152 9772 12164
rect 8757 12124 9772 12152
rect 8757 12121 8769 12124
rect 8711 12115 8769 12121
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 12066 12152 12072 12164
rect 11204 12124 12072 12152
rect 11204 12112 11210 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 4525 12087 4583 12093
rect 4525 12053 4537 12087
rect 4571 12084 4583 12087
rect 4614 12084 4620 12096
rect 4571 12056 4620 12084
rect 4571 12053 4583 12056
rect 4525 12047 4583 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5353 12087 5411 12093
rect 5353 12084 5365 12087
rect 5224 12056 5365 12084
rect 5224 12044 5230 12056
rect 5353 12053 5365 12056
rect 5399 12053 5411 12087
rect 5718 12084 5724 12096
rect 5679 12056 5724 12084
rect 5353 12047 5411 12053
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 7926 12084 7932 12096
rect 7887 12056 7932 12084
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 9950 11880 9956 11892
rect 9548 11852 9956 11880
rect 9548 11840 9554 11852
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 11606 11880 11612 11892
rect 11567 11852 11612 11880
rect 11606 11840 11612 11852
rect 11664 11880 11670 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 11664 11852 12173 11880
rect 11664 11840 11670 11852
rect 12161 11849 12173 11852
rect 12207 11880 12219 11883
rect 12618 11880 12624 11892
rect 12207 11852 12624 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 3973 11815 4031 11821
rect 3973 11781 3985 11815
rect 4019 11812 4031 11815
rect 5166 11812 5172 11824
rect 4019 11784 5172 11812
rect 4019 11781 4031 11784
rect 3973 11775 4031 11781
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 7926 11772 7932 11824
rect 7984 11812 7990 11824
rect 10318 11812 10324 11824
rect 7984 11784 10324 11812
rect 7984 11772 7990 11784
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 6273 11747 6331 11753
rect 6273 11744 6285 11747
rect 5776 11716 6285 11744
rect 5776 11704 5782 11716
rect 6273 11713 6285 11716
rect 6319 11744 6331 11747
rect 6319 11716 7144 11744
rect 6319 11713 6331 11716
rect 6273 11707 6331 11713
rect 4430 11676 4436 11688
rect 4391 11648 4436 11676
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 5166 11676 5172 11688
rect 5127 11648 5172 11676
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 5261 11679 5319 11685
rect 5261 11645 5273 11679
rect 5307 11645 5319 11679
rect 5626 11676 5632 11688
rect 5587 11648 5632 11676
rect 5261 11639 5319 11645
rect 5276 11608 5304 11639
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6564 11648 6837 11676
rect 4356 11580 5304 11608
rect 4356 11552 4384 11580
rect 3602 11540 3608 11552
rect 3563 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 4522 11540 4528 11552
rect 4483 11512 4528 11540
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 6564 11549 6592 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 7116 11676 7144 11716
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 12158 11744 12164 11756
rect 8812 11716 12164 11744
rect 8812 11704 8818 11716
rect 12158 11704 12164 11716
rect 12216 11744 12222 11756
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12216 11716 12817 11744
rect 12216 11704 12222 11716
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 7116 11648 7297 11676
rect 6825 11639 6883 11645
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 7524 11648 7665 11676
rect 7524 11636 7530 11648
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 8018 11676 8024 11688
rect 7931 11648 8024 11676
rect 7653 11639 7711 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8570 11636 8576 11688
rect 8628 11676 8634 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 8628 11648 8953 11676
rect 8628 11636 8634 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 9122 11676 9128 11688
rect 9083 11648 9128 11676
rect 8941 11639 8999 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 7006 11568 7012 11620
rect 7064 11608 7070 11620
rect 8036 11608 8064 11636
rect 7064 11580 8064 11608
rect 7064 11568 7070 11580
rect 8662 11568 8668 11620
rect 8720 11608 8726 11620
rect 9876 11608 9904 11639
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10318 11676 10324 11688
rect 10008 11648 10053 11676
rect 10279 11648 10324 11676
rect 10008 11636 10014 11648
rect 10318 11636 10324 11648
rect 10376 11676 10382 11688
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10376 11648 10885 11676
rect 10376 11636 10382 11648
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11241 11611 11299 11617
rect 11241 11608 11253 11611
rect 8720 11580 11253 11608
rect 8720 11568 8726 11580
rect 11241 11577 11253 11580
rect 11287 11577 11299 11611
rect 11241 11571 11299 11577
rect 12529 11611 12587 11617
rect 12529 11577 12541 11611
rect 12575 11577 12587 11611
rect 12529 11571 12587 11577
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 4672 11512 6561 11540
rect 4672 11500 4678 11512
rect 6549 11509 6561 11512
rect 6595 11509 6607 11543
rect 6914 11540 6920 11552
rect 6875 11512 6920 11540
rect 6549 11503 6607 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8444 11512 8585 11540
rect 8444 11500 8450 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9364 11512 9413 11540
rect 9364 11500 9370 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12544 11540 12572 11571
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 12676 11580 12721 11608
rect 12676 11568 12682 11580
rect 12492 11512 12572 11540
rect 12492 11500 12498 11512
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3660 11308 3801 11336
rect 3660 11296 3666 11308
rect 3789 11305 3801 11308
rect 3835 11336 3847 11339
rect 4154 11336 4160 11348
rect 3835 11308 4160 11336
rect 3835 11305 3847 11308
rect 3789 11299 3847 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4430 11336 4436 11348
rect 4391 11308 4436 11336
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5718 11336 5724 11348
rect 5307 11308 5724 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7190 11296 7196 11348
rect 7248 11336 7254 11348
rect 9122 11336 9128 11348
rect 7248 11308 9128 11336
rect 7248 11296 7254 11308
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 10042 11336 10048 11348
rect 10003 11308 10048 11336
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 4448 11268 4476 11296
rect 6730 11268 6736 11280
rect 4448 11240 5672 11268
rect 6643 11240 6736 11268
rect 5644 11212 5672 11240
rect 4614 11200 4620 11212
rect 4575 11172 4620 11200
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5626 11200 5632 11212
rect 5539 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 6104 11132 6132 11163
rect 6178 11160 6184 11212
rect 6236 11200 6242 11212
rect 6656 11209 6684 11240
rect 6730 11228 6736 11240
rect 6788 11268 6794 11280
rect 7466 11268 7472 11280
rect 6788 11240 7472 11268
rect 6788 11228 6794 11240
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 8205 11271 8263 11277
rect 8205 11237 8217 11271
rect 8251 11268 8263 11271
rect 8846 11268 8852 11280
rect 8251 11240 8852 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 11609 11271 11667 11277
rect 11609 11268 11621 11271
rect 10612 11240 11621 11268
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6236 11172 6653 11200
rect 6236 11160 6242 11172
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 7006 11200 7012 11212
rect 6967 11172 7012 11200
rect 6641 11163 6699 11169
rect 7006 11160 7012 11172
rect 7064 11160 7070 11212
rect 8864 11200 8892 11228
rect 10612 11209 10640 11240
rect 11609 11237 11621 11240
rect 11655 11268 11667 11271
rect 11790 11268 11796 11280
rect 11655 11240 11796 11268
rect 11655 11237 11667 11240
rect 11609 11231 11667 11237
rect 11790 11228 11796 11240
rect 11848 11228 11854 11280
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 8864 11172 10609 11200
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 7466 11132 7472 11144
rect 5224 11104 7472 11132
rect 5224 11092 5230 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 8110 11132 8116 11144
rect 8071 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11092 8174 11144
rect 8754 11132 8760 11144
rect 8715 11104 8760 11132
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 9674 11132 9680 11144
rect 9635 11104 9680 11132
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 11514 11132 11520 11144
rect 11475 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 4801 11067 4859 11073
rect 4801 11033 4813 11067
rect 4847 11064 4859 11067
rect 7190 11064 7196 11076
rect 4847 11036 7196 11064
rect 4847 11033 4859 11036
rect 4801 11027 4859 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 10410 11024 10416 11076
rect 10468 11064 10474 11076
rect 11808 11064 11836 11095
rect 12066 11064 12072 11076
rect 10468 11036 12072 11064
rect 10468 11024 10474 11036
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 7837 10999 7895 11005
rect 7837 10965 7849 10999
rect 7883 10996 7895 10999
rect 8018 10996 8024 11008
rect 7883 10968 8024 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 8018 10956 8024 10968
rect 8076 10956 8082 11008
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 10873 10999 10931 11005
rect 10873 10996 10885 10999
rect 10836 10968 10885 10996
rect 10836 10956 10842 10968
rect 10873 10965 10885 10968
rect 10919 10965 10931 10999
rect 12434 10996 12440 11008
rect 12395 10968 12440 10996
rect 10873 10959 10931 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6178 10792 6184 10804
rect 5951 10764 6184 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6638 10792 6644 10804
rect 6319 10764 6644 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 10134 10792 10140 10804
rect 10095 10764 10140 10792
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11103 10795 11161 10801
rect 11103 10761 11115 10795
rect 11149 10792 11161 10795
rect 11514 10792 11520 10804
rect 11149 10764 11520 10792
rect 11149 10761 11161 10764
rect 11103 10755 11161 10761
rect 11514 10752 11520 10764
rect 11572 10792 11578 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11572 10764 12173 10792
rect 11572 10752 11578 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 8570 10724 8576 10736
rect 7984 10696 8576 10724
rect 7984 10684 7990 10696
rect 8570 10684 8576 10696
rect 8628 10724 8634 10736
rect 8941 10727 8999 10733
rect 8941 10724 8953 10727
rect 8628 10696 8953 10724
rect 8628 10684 8634 10696
rect 8941 10693 8953 10696
rect 8987 10724 8999 10727
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 8987 10696 9045 10724
rect 8987 10693 8999 10696
rect 8941 10687 8999 10693
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 11790 10724 11796 10736
rect 11751 10696 11796 10724
rect 9033 10687 9091 10693
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 4430 10616 4436 10668
rect 4488 10656 4494 10668
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 4488 10628 4813 10656
rect 4488 10616 4494 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 9674 10656 9680 10668
rect 8435 10628 9680 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 9674 10616 9680 10628
rect 9732 10656 9738 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 9732 10628 10793 10656
rect 9732 10616 9738 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 10781 10619 10839 10625
rect 4614 10588 4620 10600
rect 4527 10560 4620 10588
rect 4614 10548 4620 10560
rect 4672 10588 4678 10600
rect 4893 10591 4951 10597
rect 4893 10588 4905 10591
rect 4672 10560 4905 10588
rect 4672 10548 4678 10560
rect 4893 10557 4905 10560
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7190 10588 7196 10600
rect 6687 10560 7196 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 4246 10452 4252 10464
rect 4207 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10452 4310 10464
rect 4632 10461 4660 10548
rect 7466 10480 7472 10532
rect 7524 10520 7530 10532
rect 7668 10520 7696 10551
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 7800 10560 7845 10588
rect 7800 10548 7806 10560
rect 8018 10548 8024 10600
rect 8076 10588 8082 10600
rect 8113 10591 8171 10597
rect 8113 10588 8125 10591
rect 8076 10560 8125 10588
rect 8076 10548 8082 10560
rect 8113 10557 8125 10560
rect 8159 10557 8171 10591
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 8113 10551 8171 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 11032 10591 11090 10597
rect 11032 10557 11044 10591
rect 11078 10588 11090 10591
rect 11078 10560 11560 10588
rect 11078 10557 11090 10560
rect 11032 10551 11090 10557
rect 8570 10520 8576 10532
rect 7524 10492 8576 10520
rect 7524 10480 7530 10492
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 8941 10523 8999 10529
rect 8941 10489 8953 10523
rect 8987 10520 8999 10523
rect 9538 10523 9596 10529
rect 9538 10520 9550 10523
rect 8987 10492 9550 10520
rect 8987 10489 8999 10492
rect 8941 10483 8999 10489
rect 9538 10489 9550 10492
rect 9584 10520 9596 10523
rect 10042 10520 10048 10532
rect 9584 10492 10048 10520
rect 9584 10489 9596 10492
rect 9538 10483 9596 10489
rect 10042 10480 10048 10492
rect 10100 10520 10106 10532
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 10100 10492 10425 10520
rect 10100 10480 10106 10492
rect 10413 10489 10425 10492
rect 10459 10489 10471 10523
rect 10413 10483 10471 10489
rect 4617 10455 4675 10461
rect 4617 10452 4629 10455
rect 4304 10424 4629 10452
rect 4304 10412 4310 10424
rect 4617 10421 4629 10424
rect 4663 10421 4675 10455
rect 4617 10415 4675 10421
rect 7742 10412 7748 10464
rect 7800 10452 7806 10464
rect 8294 10452 8300 10464
rect 7800 10424 8300 10452
rect 7800 10412 7806 10424
rect 8294 10412 8300 10424
rect 8352 10452 8358 10464
rect 11532 10461 11560 10560
rect 8665 10455 8723 10461
rect 8665 10452 8677 10455
rect 8352 10424 8677 10452
rect 8352 10412 8358 10424
rect 8665 10421 8677 10424
rect 8711 10421 8723 10455
rect 8665 10415 8723 10421
rect 11517 10455 11575 10461
rect 11517 10421 11529 10455
rect 11563 10452 11575 10455
rect 13446 10452 13452 10464
rect 11563 10424 13452 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 5626 10248 5632 10260
rect 5587 10220 5632 10248
rect 5626 10208 5632 10220
rect 5684 10208 5690 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 8662 10248 8668 10260
rect 8619 10220 8668 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 8846 10248 8852 10260
rect 8807 10220 8852 10248
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 11379 10251 11437 10257
rect 11379 10217 11391 10251
rect 11425 10248 11437 10251
rect 12434 10248 12440 10260
rect 11425 10220 12440 10248
rect 11425 10217 11437 10220
rect 11379 10211 11437 10217
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 5353 10183 5411 10189
rect 5353 10149 5365 10183
rect 5399 10180 5411 10183
rect 8205 10183 8263 10189
rect 5399 10152 7512 10180
rect 5399 10149 5411 10152
rect 5353 10143 5411 10149
rect 7484 10124 7512 10152
rect 8205 10149 8217 10183
rect 8251 10180 8263 10183
rect 9214 10180 9220 10192
rect 8251 10152 9220 10180
rect 8251 10149 8263 10152
rect 8205 10143 8263 10149
rect 9214 10140 9220 10152
rect 9272 10140 9278 10192
rect 9766 10180 9772 10192
rect 9727 10152 9772 10180
rect 9766 10140 9772 10152
rect 9824 10140 9830 10192
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 10134 10180 10140 10192
rect 9907 10152 10140 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 10410 10180 10416 10192
rect 10371 10152 10416 10180
rect 10410 10140 10416 10152
rect 10468 10140 10474 10192
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 5684 10084 6745 10112
rect 5684 10072 5690 10084
rect 6733 10081 6745 10084
rect 6779 10112 6791 10115
rect 6822 10112 6828 10124
rect 6779 10084 6828 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7466 10112 7472 10124
rect 7427 10084 7472 10112
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10112 7619 10115
rect 7742 10112 7748 10124
rect 7607 10084 7748 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 7576 10044 7604 10075
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8018 10112 8024 10124
rect 7979 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10112 11299 10115
rect 11330 10112 11336 10124
rect 11287 10084 11336 10112
rect 11287 10081 11299 10084
rect 11241 10075 11299 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 7024 10016 7604 10044
rect 7024 9920 7052 10016
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4522 9908 4528 9920
rect 4212 9880 4528 9908
rect 4212 9868 4218 9880
rect 4522 9868 4528 9880
rect 4580 9908 4586 9920
rect 4893 9911 4951 9917
rect 4893 9908 4905 9911
rect 4580 9880 4905 9908
rect 4580 9868 4586 9880
rect 4893 9877 4905 9880
rect 4939 9877 4951 9911
rect 4893 9871 4951 9877
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 6641 9911 6699 9917
rect 6641 9908 6653 9911
rect 6319 9880 6653 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 6641 9877 6653 9880
rect 6687 9908 6699 9911
rect 7006 9908 7012 9920
rect 6687 9880 7012 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 5261 9707 5319 9713
rect 5261 9673 5273 9707
rect 5307 9704 5319 9707
rect 5626 9704 5632 9716
rect 5307 9676 5632 9704
rect 5307 9673 5319 9676
rect 5261 9667 5319 9673
rect 5626 9664 5632 9676
rect 5684 9664 5690 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8720 9676 8953 9704
rect 8720 9664 8726 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 8941 9667 8999 9673
rect 10134 9664 10140 9716
rect 10192 9704 10198 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 10192 9676 10241 9704
rect 10192 9664 10198 9676
rect 10229 9673 10241 9676
rect 10275 9673 10287 9707
rect 10229 9667 10287 9673
rect 6638 9636 6644 9648
rect 6551 9608 6644 9636
rect 6638 9596 6644 9608
rect 6696 9636 6702 9648
rect 7650 9636 7656 9648
rect 6696 9608 7656 9636
rect 6696 9596 6702 9608
rect 7650 9596 7656 9608
rect 7708 9596 7714 9648
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 10551 9639 10609 9645
rect 10551 9636 10563 9639
rect 8168 9608 10563 9636
rect 8168 9596 8174 9608
rect 10551 9605 10563 9608
rect 10597 9605 10609 9639
rect 10551 9599 10609 9605
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 10778 9568 10784 9580
rect 8343 9540 10784 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 6822 9500 6828 9512
rect 5767 9472 6224 9500
rect 6783 9472 6828 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 6196 9376 6224 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7576 9432 7604 9463
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7708 9472 7757 9500
rect 7708 9460 7714 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 8018 9500 8024 9512
rect 7979 9472 8024 9500
rect 7745 9463 7803 9469
rect 8018 9460 8024 9472
rect 8076 9500 8082 9512
rect 9490 9509 9496 9512
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 8076 9472 8585 9500
rect 8076 9460 8082 9472
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 9468 9503 9496 9509
rect 9468 9500 9480 9503
rect 9403 9472 9480 9500
rect 8573 9463 8631 9469
rect 9468 9469 9480 9472
rect 9548 9500 9554 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9548 9472 9873 9500
rect 9468 9463 9496 9469
rect 9490 9460 9496 9463
rect 9548 9460 9554 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 10448 9503 10506 9509
rect 10448 9500 10460 9503
rect 9861 9463 9919 9469
rect 9968 9472 10460 9500
rect 8662 9432 8668 9444
rect 7576 9404 8668 9432
rect 8662 9392 8668 9404
rect 8720 9392 8726 9444
rect 9968 9432 9996 9472
rect 10448 9469 10460 9472
rect 10494 9500 10506 9503
rect 10686 9500 10692 9512
rect 10494 9472 10692 9500
rect 10494 9469 10506 9472
rect 10448 9463 10506 9469
rect 10686 9460 10692 9472
rect 10744 9500 10750 9512
rect 10873 9503 10931 9509
rect 10873 9500 10885 9503
rect 10744 9472 10885 9500
rect 10744 9460 10750 9472
rect 10873 9469 10885 9472
rect 10919 9469 10931 9503
rect 10873 9463 10931 9469
rect 8817 9404 9996 9432
rect 5902 9364 5908 9376
rect 5863 9336 5908 9364
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 8817 9364 8845 9404
rect 7156 9336 8845 9364
rect 9539 9367 9597 9373
rect 7156 9324 7162 9336
rect 9539 9333 9551 9367
rect 9585 9364 9597 9367
rect 9674 9364 9680 9376
rect 9585 9336 9680 9364
rect 9585 9333 9597 9336
rect 9539 9327 9597 9333
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 11330 9364 11336 9376
rect 11243 9336 11336 9364
rect 11330 9324 11336 9336
rect 11388 9364 11394 9376
rect 12066 9364 12072 9376
rect 11388 9336 12072 9364
rect 11388 9324 11394 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 6733 9163 6791 9169
rect 6733 9160 6745 9163
rect 5960 9132 6745 9160
rect 5960 9120 5966 9132
rect 6733 9129 6745 9132
rect 6779 9160 6791 9163
rect 8018 9160 8024 9172
rect 6779 9132 8024 9160
rect 6779 9129 6791 9132
rect 6733 9123 6791 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 8168 9132 8585 9160
rect 8168 9120 8174 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9766 9160 9772 9172
rect 9539 9132 9772 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 11422 9120 11428 9172
rect 11480 9160 11486 9172
rect 11655 9163 11713 9169
rect 11655 9160 11667 9163
rect 11480 9132 11667 9160
rect 11480 9120 11486 9132
rect 11655 9129 11667 9132
rect 11701 9129 11713 9163
rect 11655 9123 11713 9129
rect 12667 9163 12725 9169
rect 12667 9129 12679 9163
rect 12713 9160 12725 9163
rect 13814 9160 13820 9172
rect 12713 9132 13820 9160
rect 12713 9129 12725 9132
rect 12667 9123 12725 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 8297 9095 8355 9101
rect 8297 9061 8309 9095
rect 8343 9092 8355 9095
rect 8662 9092 8668 9104
rect 8343 9064 8668 9092
rect 8343 9061 8355 9064
rect 8297 9055 8355 9061
rect 8662 9052 8668 9064
rect 8720 9052 8726 9104
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5316 8996 5641 9024
rect 5316 8984 5322 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 7006 8984 7012 9036
rect 7064 9024 7070 9036
rect 7193 9027 7251 9033
rect 7193 9024 7205 9027
rect 7064 8996 7205 9024
rect 7064 8984 7070 8996
rect 7193 8993 7205 8996
rect 7239 8993 7251 9027
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 7193 8987 7251 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 10318 9024 10324 9036
rect 10279 8996 10324 9024
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 11514 9024 11520 9036
rect 11475 8996 11520 9024
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 12575 9027 12633 9033
rect 12575 8993 12587 9027
rect 12621 8993 12633 9027
rect 12575 8987 12633 8993
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5776 8928 6009 8956
rect 5776 8916 5782 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8956 6423 8959
rect 7282 8956 7288 8968
rect 6411 8928 7288 8956
rect 6411 8925 6423 8928
rect 6365 8919 6423 8925
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7742 8956 7748 8968
rect 7703 8928 7748 8956
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 12590 8900 12618 8987
rect 4908 8860 5810 8888
rect 4908 8832 4936 8860
rect 4890 8820 4896 8832
rect 4851 8792 4896 8820
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 5258 8820 5264 8832
rect 5219 8792 5264 8820
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5782 8829 5810 8860
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 8536 8860 9045 8888
rect 8536 8848 8542 8860
rect 9033 8857 9045 8860
rect 9079 8888 9091 8891
rect 10502 8888 10508 8900
rect 9079 8860 10508 8888
rect 9079 8857 9091 8860
rect 9033 8851 9091 8857
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 12590 8860 12624 8900
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 5767 8823 5825 8829
rect 5767 8789 5779 8823
rect 5813 8789 5825 8823
rect 5902 8820 5908 8832
rect 5863 8792 5908 8820
rect 5767 8783 5825 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 9950 8820 9956 8832
rect 9911 8792 9956 8820
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 6638 8616 6644 8628
rect 6599 8588 6644 8616
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 9861 8619 9919 8625
rect 9861 8585 9873 8619
rect 9907 8616 9919 8619
rect 9950 8616 9956 8628
rect 9907 8588 9956 8616
rect 9907 8585 9919 8588
rect 9861 8579 9919 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10376 8588 10977 8616
rect 10376 8576 10382 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 13630 8616 13636 8628
rect 13591 8588 13636 8616
rect 10965 8579 11023 8585
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 4341 8551 4399 8557
rect 4341 8517 4353 8551
rect 4387 8548 4399 8551
rect 4890 8548 4896 8560
rect 4387 8520 4896 8548
rect 4387 8517 4399 8520
rect 4341 8511 4399 8517
rect 4890 8508 4896 8520
rect 4948 8548 4954 8560
rect 5307 8551 5365 8557
rect 5307 8548 5319 8551
rect 4948 8520 5319 8548
rect 4948 8508 4954 8520
rect 5307 8517 5319 8520
rect 5353 8517 5365 8551
rect 5442 8548 5448 8560
rect 5403 8520 5448 8548
rect 5307 8511 5365 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5132 8452 5549 8480
rect 5132 8440 5138 8452
rect 5537 8449 5549 8452
rect 5583 8449 5595 8483
rect 5537 8443 5595 8449
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5868 8452 5917 8480
rect 5868 8440 5874 8452
rect 5905 8449 5917 8452
rect 5951 8480 5963 8483
rect 7650 8480 7656 8492
rect 5951 8452 7656 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 8478 8480 8484 8492
rect 8439 8452 8484 8480
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8720 8452 8769 8480
rect 8720 8440 8726 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 9539 8452 10057 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 10045 8449 10057 8452
rect 10091 8480 10103 8483
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 10091 8452 12449 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 5718 8412 5724 8424
rect 4755 8384 5724 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6696 8384 6837 8412
rect 6696 8372 6702 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 7282 8412 7288 8424
rect 7243 8384 7288 8412
rect 6825 8375 6883 8381
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8412 13507 8415
rect 13722 8412 13728 8424
rect 13495 8384 13728 8412
rect 13495 8381 13507 8384
rect 13449 8375 13507 8381
rect 13722 8372 13728 8384
rect 13780 8412 13786 8424
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13780 8384 14013 8412
rect 13780 8372 13786 8384
rect 14001 8381 14013 8384
rect 14047 8381 14059 8415
rect 14001 8375 14059 8381
rect 5166 8344 5172 8356
rect 5127 8316 5172 8344
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 5442 8344 5448 8356
rect 5316 8316 5448 8344
rect 5316 8304 5322 8316
rect 5442 8304 5448 8316
rect 5500 8344 5506 8356
rect 5902 8344 5908 8356
rect 5500 8316 5908 8344
rect 5500 8304 5506 8316
rect 5902 8304 5908 8316
rect 5960 8344 5966 8356
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 5960 8316 6193 8344
rect 5960 8304 5966 8316
rect 6181 8313 6193 8316
rect 6227 8313 6239 8347
rect 6181 8307 6239 8313
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8344 7619 8347
rect 8202 8344 8208 8356
rect 7607 8316 8208 8344
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 8573 8347 8631 8353
rect 8573 8313 8585 8347
rect 8619 8313 8631 8347
rect 8573 8307 8631 8313
rect 10137 8347 10195 8353
rect 10137 8313 10149 8347
rect 10183 8313 10195 8347
rect 10137 8307 10195 8313
rect 5074 8276 5080 8288
rect 5035 8248 5080 8276
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7064 8248 7849 8276
rect 7064 8236 7070 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 8294 8276 8300 8288
rect 8255 8248 8300 8276
rect 7837 8239 7895 8245
rect 8294 8236 8300 8248
rect 8352 8276 8358 8288
rect 8588 8276 8616 8307
rect 8352 8248 8616 8276
rect 8352 8236 8358 8248
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10152 8276 10180 8307
rect 10410 8304 10416 8356
rect 10468 8344 10474 8356
rect 10689 8347 10747 8353
rect 10689 8344 10701 8347
rect 10468 8316 10701 8344
rect 10468 8304 10474 8316
rect 10689 8313 10701 8316
rect 10735 8344 10747 8347
rect 12618 8344 12624 8356
rect 10735 8316 12624 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 12618 8304 12624 8316
rect 12676 8344 12682 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12676 8316 12909 8344
rect 12676 8304 12682 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 10008 8248 10180 8276
rect 10008 8236 10014 8248
rect 11054 8236 11060 8288
rect 11112 8276 11118 8288
rect 11514 8276 11520 8288
rect 11112 8248 11520 8276
rect 11112 8236 11118 8248
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 4522 8072 4528 8084
rect 4483 8044 4528 8072
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7650 8072 7656 8084
rect 7331 8044 7656 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 10318 8072 10324 8084
rect 8803 8044 10324 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8158 8007 8216 8013
rect 8158 8004 8170 8007
rect 7984 7976 8170 8004
rect 7984 7964 7990 7976
rect 8158 7973 8170 7976
rect 8204 7973 8216 8007
rect 8158 7967 8216 7973
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 9876 8013 9904 8044
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 9861 8007 9919 8013
rect 9861 8004 9873 8007
rect 9824 7976 9873 8004
rect 9824 7964 9830 7976
rect 9861 7973 9873 7976
rect 9907 7973 9919 8007
rect 10410 8004 10416 8016
rect 10371 7976 10416 8004
rect 9861 7967 9919 7973
rect 10410 7964 10416 7976
rect 10468 7964 10474 8016
rect 11425 8007 11483 8013
rect 11425 7973 11437 8007
rect 11471 8004 11483 8007
rect 11514 8004 11520 8016
rect 11471 7976 11520 8004
rect 11471 7973 11483 7976
rect 11425 7967 11483 7973
rect 11514 7964 11520 7976
rect 11572 7964 11578 8016
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 4387 7908 4936 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4908 7809 4936 7908
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 5316 7908 5365 7936
rect 5316 7896 5322 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5500 7871 5558 7877
rect 5500 7837 5512 7871
rect 5546 7868 5558 7871
rect 5626 7868 5632 7880
rect 5546 7840 5632 7868
rect 5546 7837 5558 7840
rect 5500 7831 5558 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 5902 7868 5908 7880
rect 5767 7840 5908 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 4939 7772 5825 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 5813 7769 5825 7772
rect 5859 7769 5871 7803
rect 5813 7763 5871 7769
rect 6917 7803 6975 7809
rect 6917 7769 6929 7803
rect 6963 7800 6975 7803
rect 7282 7800 7288 7812
rect 6963 7772 7288 7800
rect 6963 7769 6975 7772
rect 6917 7763 6975 7769
rect 7282 7760 7288 7772
rect 7340 7760 7346 7812
rect 5258 7732 5264 7744
rect 5219 7704 5264 7732
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5350 7692 5356 7744
rect 5408 7732 5414 7744
rect 5629 7735 5687 7741
rect 5629 7732 5641 7735
rect 5408 7704 5641 7732
rect 5408 7692 5414 7704
rect 5629 7701 5641 7704
rect 5675 7732 5687 7735
rect 6365 7735 6423 7741
rect 6365 7732 6377 7735
rect 5675 7704 6377 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 6365 7701 6377 7704
rect 6411 7732 6423 7735
rect 6546 7732 6552 7744
rect 6411 7704 6552 7732
rect 6411 7701 6423 7704
rect 6365 7695 6423 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7650 7732 7656 7744
rect 7611 7704 7656 7732
rect 7650 7692 7656 7704
rect 7708 7732 7714 7744
rect 7852 7732 7880 7831
rect 8662 7828 8668 7880
rect 8720 7868 8726 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 8720 7840 9781 7868
rect 8720 7828 8726 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 11790 7868 11796 7880
rect 11379 7840 11796 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11790 7828 11796 7840
rect 11848 7868 11854 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 11848 7840 12817 7868
rect 11848 7828 11854 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 11885 7803 11943 7809
rect 11885 7800 11897 7803
rect 11112 7772 11897 7800
rect 11112 7760 11118 7772
rect 11885 7769 11897 7772
rect 11931 7769 11943 7803
rect 11885 7763 11943 7769
rect 7708 7704 7880 7732
rect 7708 7692 7714 7704
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 5718 7528 5724 7540
rect 5675 7500 5724 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6546 7528 6552 7540
rect 6507 7500 6552 7528
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 4798 7460 4804 7472
rect 3559 7432 4804 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 3620 7333 3648 7432
rect 4798 7420 4804 7432
rect 4856 7460 4862 7472
rect 6638 7460 6644 7472
rect 4856 7432 6644 7460
rect 4856 7420 4862 7432
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 7374 7420 7380 7472
rect 7432 7460 7438 7472
rect 12575 7463 12633 7469
rect 12575 7460 12587 7463
rect 7432 7432 12587 7460
rect 7432 7420 7438 7432
rect 12575 7429 12587 7432
rect 12621 7429 12633 7463
rect 12575 7423 12633 7429
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 7650 7392 7656 7404
rect 4387 7364 7656 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8260 7364 8493 7392
rect 8260 7352 8266 7364
rect 8481 7361 8493 7364
rect 8527 7392 8539 7395
rect 9030 7392 9036 7404
rect 8527 7364 9036 7392
rect 8527 7361 8539 7364
rect 8481 7355 8539 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 11054 7392 11060 7404
rect 11015 7364 11060 7392
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 3752 7296 4169 7324
rect 3752 7284 3758 7296
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 5258 7324 5264 7336
rect 4755 7296 5264 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 4172 7256 4200 7287
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5442 7324 5448 7336
rect 5403 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9447 7296 10149 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 12504 7327 12562 7333
rect 12504 7293 12516 7327
rect 12550 7324 12562 7327
rect 12894 7324 12900 7336
rect 12550 7296 12900 7324
rect 12550 7293 12562 7296
rect 12504 7287 12562 7293
rect 5810 7256 5816 7268
rect 4172 7228 5816 7256
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7225 7067 7259
rect 7009 7219 7067 7225
rect 5074 7188 5080 7200
rect 4987 7160 5080 7188
rect 5074 7148 5080 7160
rect 5132 7188 5138 7200
rect 5442 7188 5448 7200
rect 5132 7160 5448 7188
rect 5132 7148 5138 7160
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5902 7148 5908 7200
rect 5960 7188 5966 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 5960 7160 6193 7188
rect 5960 7148 5966 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 7024 7188 7052 7219
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 7653 7259 7711 7265
rect 7156 7228 7201 7256
rect 7156 7216 7162 7228
rect 7653 7225 7665 7259
rect 7699 7256 7711 7259
rect 8662 7256 8668 7268
rect 7699 7228 8668 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 8802 7259 8860 7265
rect 8802 7225 8814 7259
rect 8848 7225 8860 7259
rect 8802 7219 8860 7225
rect 7374 7188 7380 7200
rect 7024 7160 7380 7188
rect 6181 7151 6239 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7926 7188 7932 7200
rect 7887 7160 7932 7188
rect 7926 7148 7932 7160
rect 7984 7188 7990 7200
rect 8297 7191 8355 7197
rect 8297 7188 8309 7191
rect 7984 7160 8309 7188
rect 7984 7148 7990 7160
rect 8297 7157 8309 7160
rect 8343 7188 8355 7191
rect 8817 7188 8845 7219
rect 8343 7160 8845 7188
rect 10152 7188 10180 7287
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 10410 7256 10416 7268
rect 10371 7228 10416 7256
rect 10410 7216 10416 7228
rect 10468 7216 10474 7268
rect 10505 7259 10563 7265
rect 10505 7225 10517 7259
rect 10551 7225 10563 7259
rect 10505 7219 10563 7225
rect 10520 7188 10548 7219
rect 11330 7188 11336 7200
rect 10152 7160 11336 7188
rect 8343 7157 8355 7160
rect 8297 7151 8355 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11425 7191 11483 7197
rect 11425 7157 11437 7191
rect 11471 7188 11483 7191
rect 11514 7188 11520 7200
rect 11471 7160 11520 7188
rect 11471 7157 11483 7160
rect 11425 7151 11483 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 3694 6984 3700 6996
rect 3655 6956 3700 6984
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 5353 6987 5411 6993
rect 5353 6953 5365 6987
rect 5399 6984 5411 6987
rect 5718 6984 5724 6996
rect 5399 6956 5724 6984
rect 5399 6953 5411 6956
rect 5353 6947 5411 6953
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 7009 6987 7067 6993
rect 7009 6953 7021 6987
rect 7055 6984 7067 6987
rect 7098 6984 7104 6996
rect 7055 6956 7104 6984
rect 7055 6953 7067 6956
rect 7009 6947 7067 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 7374 6984 7380 6996
rect 7335 6956 7380 6984
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 9030 6984 9036 6996
rect 8991 6956 9036 6984
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 11514 6984 11520 6996
rect 11475 6956 11520 6984
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 6178 6916 6184 6928
rect 6139 6888 6184 6916
rect 6178 6876 6184 6888
rect 6236 6876 6242 6928
rect 7926 6876 7932 6928
rect 7984 6916 7990 6928
rect 8158 6919 8216 6925
rect 8158 6916 8170 6919
rect 7984 6888 8170 6916
rect 7984 6876 7990 6888
rect 8158 6885 8170 6888
rect 8204 6885 8216 6919
rect 9861 6919 9919 6925
rect 9861 6916 9873 6919
rect 8158 6879 8216 6885
rect 8772 6888 9873 6916
rect 4430 6848 4436 6860
rect 4391 6820 4436 6848
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 8772 6857 8800 6888
rect 9861 6885 9873 6888
rect 9907 6916 9919 6919
rect 9950 6916 9956 6928
rect 9907 6888 9956 6916
rect 9907 6885 9919 6888
rect 9861 6879 9919 6885
rect 9950 6876 9956 6888
rect 10008 6876 10014 6928
rect 10410 6916 10416 6928
rect 10371 6888 10416 6916
rect 10410 6876 10416 6888
rect 10468 6916 10474 6928
rect 10689 6919 10747 6925
rect 10689 6916 10701 6919
rect 10468 6888 10701 6916
rect 10468 6876 10474 6888
rect 10689 6885 10701 6888
rect 10735 6885 10747 6919
rect 10689 6879 10747 6885
rect 5445 6851 5503 6857
rect 5445 6848 5457 6851
rect 5408 6820 5457 6848
rect 5408 6808 5414 6820
rect 5445 6817 5457 6820
rect 5491 6817 5503 6851
rect 5445 6811 5503 6817
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6817 8815 6851
rect 11330 6848 11336 6860
rect 11291 6820 11336 6848
rect 8757 6811 8815 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5552 6752 5825 6780
rect 5442 6672 5448 6724
rect 5500 6712 5506 6724
rect 5552 6712 5580 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 5813 6743 5871 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 8720 6752 9413 6780
rect 8720 6740 8726 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9401 6743 9459 6749
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 5500 6684 5580 6712
rect 5610 6715 5668 6721
rect 5500 6672 5506 6684
rect 5610 6681 5622 6715
rect 5656 6712 5668 6715
rect 5902 6712 5908 6724
rect 5656 6684 5908 6712
rect 5656 6681 5668 6684
rect 5610 6675 5668 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6644 4675 6647
rect 5166 6644 5172 6656
rect 4663 6616 5172 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5718 6644 5724 6656
rect 5316 6616 5724 6644
rect 5316 6604 5322 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 5776 6412 6561 6440
rect 5776 6400 5782 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 8110 6440 8116 6452
rect 7156 6412 8116 6440
rect 7156 6400 7162 6412
rect 8110 6400 8116 6412
rect 8168 6440 8174 6452
rect 8573 6443 8631 6449
rect 8573 6440 8585 6443
rect 8168 6412 8585 6440
rect 8168 6400 8174 6412
rect 8573 6409 8585 6412
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 10781 6443 10839 6449
rect 10781 6440 10793 6443
rect 9824 6412 10793 6440
rect 9824 6400 9830 6412
rect 10781 6409 10793 6412
rect 10827 6409 10839 6443
rect 10781 6403 10839 6409
rect 11241 6443 11299 6449
rect 11241 6409 11253 6443
rect 11287 6440 11299 6443
rect 11330 6440 11336 6452
rect 11287 6412 11336 6440
rect 11287 6409 11299 6412
rect 11241 6403 11299 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 7009 6375 7067 6381
rect 7009 6372 7021 6375
rect 5408 6344 7021 6372
rect 5408 6332 5414 6344
rect 7009 6341 7021 6344
rect 7055 6341 7067 6375
rect 10410 6372 10416 6384
rect 10371 6344 10416 6372
rect 7009 6335 7067 6341
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 10502 6332 10508 6384
rect 10560 6372 10566 6384
rect 11471 6375 11529 6381
rect 11471 6372 11483 6375
rect 10560 6344 11483 6372
rect 10560 6332 10566 6344
rect 11471 6341 11483 6344
rect 11517 6341 11529 6375
rect 11471 6335 11529 6341
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 5169 6307 5227 6313
rect 5169 6304 5181 6307
rect 4948 6276 5181 6304
rect 4948 6264 4954 6276
rect 5169 6273 5181 6276
rect 5215 6273 5227 6307
rect 5169 6267 5227 6273
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7742 6304 7748 6316
rect 7699 6276 7748 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9950 6304 9956 6316
rect 9355 6276 9956 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9950 6264 9956 6276
rect 10008 6304 10014 6316
rect 10318 6304 10324 6316
rect 10008 6276 10324 6304
rect 10008 6264 10014 6276
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5092 6208 5273 6236
rect 4430 6128 4436 6180
rect 4488 6168 4494 6180
rect 4525 6171 4583 6177
rect 4525 6168 4537 6171
rect 4488 6140 4537 6168
rect 4488 6128 4494 6140
rect 4525 6137 4537 6140
rect 4571 6168 4583 6171
rect 4982 6168 4988 6180
rect 4571 6140 4988 6168
rect 4571 6137 4583 6140
rect 4525 6131 4583 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 5092 6112 5120 6208
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 5902 6236 5908 6248
rect 5307 6208 5908 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5902 6196 5908 6208
rect 5960 6236 5966 6248
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 5960 6208 6193 6236
rect 5960 6196 5966 6208
rect 6181 6205 6193 6208
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 7892 6208 8861 6236
rect 7892 6196 7898 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 11368 6239 11426 6245
rect 11368 6236 11380 6239
rect 10652 6208 11380 6236
rect 10652 6196 10658 6208
rect 11368 6205 11380 6208
rect 11414 6236 11426 6239
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 11414 6208 11805 6236
rect 11414 6205 11426 6208
rect 11368 6199 11426 6205
rect 11793 6205 11805 6208
rect 11839 6236 11851 6239
rect 12250 6236 12256 6248
rect 11839 6208 12256 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 7561 6171 7619 6177
rect 7561 6137 7573 6171
rect 7607 6168 7619 6171
rect 7926 6168 7932 6180
rect 7607 6140 7932 6168
rect 7607 6137 7619 6140
rect 7561 6131 7619 6137
rect 7926 6128 7932 6140
rect 7984 6177 7990 6180
rect 7984 6171 8032 6177
rect 7984 6137 7986 6171
rect 8020 6137 8032 6171
rect 9858 6168 9864 6180
rect 9819 6140 9864 6168
rect 7984 6131 8032 6137
rect 7984 6128 7990 6131
rect 9858 6128 9864 6140
rect 9916 6128 9922 6180
rect 9953 6171 10011 6177
rect 9953 6137 9965 6171
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 5074 6100 5080 6112
rect 5035 6072 5080 6100
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 9674 6100 9680 6112
rect 9635 6072 9680 6100
rect 9674 6060 9680 6072
rect 9732 6100 9738 6112
rect 9968 6100 9996 6131
rect 9732 6072 9996 6100
rect 9732 6060 9738 6072
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4856 5868 5089 5896
rect 4856 5856 4862 5868
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 5077 5859 5135 5865
rect 6365 5899 6423 5905
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 6730 5896 6736 5908
rect 6411 5868 6736 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 6380 5828 6408 5859
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9858 5896 9864 5908
rect 9539 5868 9864 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 9674 5828 9680 5840
rect 4908 5800 6408 5828
rect 9635 5800 9680 5828
rect 4908 5772 4936 5800
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 4890 5760 4896 5772
rect 4803 5732 4896 5760
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 4982 5720 4988 5772
rect 5040 5760 5046 5772
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 5040 5732 6561 5760
rect 5040 5720 5046 5732
rect 6549 5729 6561 5732
rect 6595 5760 6607 5763
rect 6638 5760 6644 5772
rect 6595 5732 6644 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 10318 5760 10324 5772
rect 10279 5732 10324 5760
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7745 5559 7803 5565
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 7926 5556 7932 5568
rect 7791 5528 7932 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 4890 5352 4896 5364
rect 4851 5324 4896 5352
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 5166 5312 5172 5364
rect 5224 5352 5230 5364
rect 7006 5352 7012 5364
rect 5224 5324 7012 5352
rect 5224 5312 5230 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 8168 5324 8217 5352
rect 8168 5312 8174 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 9631 5355 9689 5361
rect 9631 5321 9643 5355
rect 9677 5352 9689 5355
rect 9858 5352 9864 5364
rect 9677 5324 9864 5352
rect 9677 5321 9689 5324
rect 9631 5315 9689 5321
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 10318 5352 10324 5364
rect 10279 5324 10324 5352
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 5803 5188 6561 5216
rect 5803 5157 5831 5188
rect 6549 5185 6561 5188
rect 6595 5216 6607 5219
rect 6595 5188 6960 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 5788 5151 5846 5157
rect 5788 5117 5800 5151
rect 5834 5117 5846 5151
rect 5788 5111 5846 5117
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6086 5148 6092 5160
rect 5960 5120 6092 5148
rect 5960 5108 5966 5120
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6273 5083 6331 5089
rect 6273 5049 6285 5083
rect 6319 5080 6331 5083
rect 6638 5080 6644 5092
rect 6319 5052 6644 5080
rect 6319 5049 6331 5052
rect 6273 5043 6331 5049
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 6932 5080 6960 5188
rect 7024 5148 7052 5312
rect 7834 5216 7840 5228
rect 7795 5188 7840 5216
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 7024 5120 7205 5148
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 7193 5111 7251 5117
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7340 5120 7665 5148
rect 7340 5108 7346 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 9560 5151 9618 5157
rect 9560 5117 9572 5151
rect 9606 5148 9618 5151
rect 9606 5120 10088 5148
rect 9606 5117 9618 5120
rect 9560 5111 9618 5117
rect 8386 5080 8392 5092
rect 6932 5052 8392 5080
rect 8386 5040 8392 5052
rect 8444 5040 8450 5092
rect 10060 5024 10088 5120
rect 5859 5015 5917 5021
rect 5859 4981 5871 5015
rect 5905 5012 5917 5015
rect 6086 5012 6092 5024
rect 5905 4984 6092 5012
rect 5905 4981 5917 4984
rect 5859 4975 5917 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 7098 4808 7104 4820
rect 6144 4780 7104 4808
rect 6144 4768 6150 4780
rect 7098 4768 7104 4780
rect 7156 4808 7162 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 7156 4780 7297 4808
rect 7156 4768 7162 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 9766 4768 9772 4820
rect 9824 4817 9830 4820
rect 9824 4811 9873 4817
rect 9824 4777 9827 4811
rect 9861 4777 9873 4811
rect 9824 4771 9873 4777
rect 9824 4768 9830 4771
rect 106 4632 112 4684
rect 164 4672 170 4684
rect 5166 4672 5172 4684
rect 164 4644 5172 4672
rect 164 4632 170 4644
rect 5166 4632 5172 4644
rect 5224 4672 5230 4684
rect 5442 4672 5448 4684
rect 5224 4644 5448 4672
rect 5224 4632 5230 4644
rect 5442 4632 5448 4644
rect 5500 4672 5506 4684
rect 5537 4675 5595 4681
rect 5537 4672 5549 4675
rect 5500 4644 5549 4672
rect 5500 4632 5506 4644
rect 5537 4641 5549 4644
rect 5583 4641 5595 4675
rect 6178 4672 6184 4684
rect 6139 4644 6184 4672
rect 5537 4635 5595 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6730 4672 6736 4684
rect 6691 4644 6736 4672
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 8478 4672 8484 4684
rect 8439 4644 8484 4672
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 9744 4675 9802 4681
rect 9744 4641 9756 4675
rect 9790 4672 9802 4675
rect 9950 4672 9956 4684
rect 9790 4644 9956 4672
rect 9790 4641 9802 4644
rect 9744 4635 9802 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 7006 4604 7012 4616
rect 6967 4576 7012 4604
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 5350 4468 5356 4480
rect 5311 4440 5356 4468
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 8110 4468 8116 4480
rect 8071 4440 8116 4468
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5166 4264 5172 4276
rect 5127 4236 5172 4264
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6236 4236 6561 4264
rect 6236 4224 6242 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 8536 4236 9597 4264
rect 8536 4224 8542 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 9585 4227 9643 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 7098 4128 7104 4140
rect 7059 4100 7104 4128
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 10594 4128 10600 4140
rect 10203 4100 10600 4128
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 5074 4060 5080 4072
rect 3568 4032 5080 4060
rect 3568 4020 3574 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 10203 4069 10231 4100
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5132 4032 5549 4060
rect 5132 4020 5138 4032
rect 5537 4029 5549 4032
rect 5583 4060 5595 4063
rect 6181 4063 6239 4069
rect 6181 4060 6193 4063
rect 5583 4032 6193 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 6181 4029 6193 4032
rect 6227 4029 6239 4063
rect 10188 4063 10246 4069
rect 10188 4060 10200 4063
rect 10166 4032 10200 4060
rect 6181 4023 6239 4029
rect 10188 4029 10200 4032
rect 10234 4029 10246 4063
rect 10188 4023 10246 4029
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 5350 3992 5356 4004
rect 4948 3964 5356 3992
rect 4948 3952 4954 3964
rect 5350 3952 5356 3964
rect 5408 3952 5414 4004
rect 6362 3952 6368 4004
rect 6420 3952 6426 4004
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3961 7251 3995
rect 7193 3955 7251 3961
rect 7745 3995 7803 4001
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 8018 3992 8024 4004
rect 7791 3964 8024 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 5626 3924 5632 3936
rect 5587 3896 5632 3924
rect 5626 3884 5632 3896
rect 5684 3924 5690 3936
rect 6380 3924 6408 3952
rect 7208 3924 7236 3955
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 8113 3995 8171 4001
rect 8113 3961 8125 3995
rect 8159 3992 8171 3995
rect 8662 3992 8668 4004
rect 8159 3964 8668 3992
rect 8159 3961 8171 3964
rect 8113 3955 8171 3961
rect 8662 3952 8668 3964
rect 8720 3952 8726 4004
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 9306 3992 9312 4004
rect 8812 3964 8857 3992
rect 9267 3964 9312 3992
rect 8812 3952 8818 3964
rect 9306 3952 9312 3964
rect 9364 3992 9370 4004
rect 9950 3992 9956 4004
rect 9364 3964 9956 3992
rect 9364 3952 9370 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 7282 3924 7288 3936
rect 5684 3896 6408 3924
rect 7195 3896 7288 3924
rect 5684 3884 5690 3896
rect 7282 3884 7288 3896
rect 7340 3924 7346 3936
rect 8386 3924 8392 3936
rect 7340 3896 8392 3924
rect 7340 3884 7346 3896
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8772 3924 8800 3952
rect 8527 3896 8800 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 10275 3927 10333 3933
rect 10275 3924 10287 3927
rect 8904 3896 10287 3924
rect 8904 3884 8910 3896
rect 10275 3893 10287 3896
rect 10321 3893 10333 3927
rect 10275 3887 10333 3893
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 7064 3692 7573 3720
rect 7064 3680 7070 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 7282 3652 7288 3664
rect 5684 3624 6316 3652
rect 7243 3624 7288 3652
rect 5684 3612 5690 3624
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5224 3556 5457 3584
rect 5224 3544 5230 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 6178 3584 6184 3596
rect 6139 3556 6184 3584
rect 5445 3547 5503 3553
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 6288 3593 6316 3624
rect 7282 3612 7288 3624
rect 7340 3612 7346 3664
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3553 6331 3587
rect 6638 3584 6644 3596
rect 6599 3556 6644 3584
rect 6273 3547 6331 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7576 3584 7604 3683
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 8720 3692 11253 3720
rect 8720 3680 8726 3692
rect 11241 3689 11253 3692
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 7926 3612 7932 3664
rect 7984 3652 7990 3664
rect 8066 3655 8124 3661
rect 8066 3652 8078 3655
rect 7984 3624 8078 3652
rect 7984 3612 7990 3624
rect 8066 3621 8078 3624
rect 8112 3621 8124 3655
rect 8066 3615 8124 3621
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 9677 3655 9735 3661
rect 9677 3652 9689 3655
rect 8812 3624 9689 3652
rect 8812 3612 8818 3624
rect 9677 3621 9689 3624
rect 9723 3621 9735 3655
rect 9677 3615 9735 3621
rect 7745 3587 7803 3593
rect 7745 3584 7757 3587
rect 7576 3556 7757 3584
rect 7745 3553 7757 3556
rect 7791 3553 7803 3587
rect 7745 3547 7803 3553
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 9766 3584 9772 3596
rect 8711 3556 9772 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 8018 3476 8024 3528
rect 8076 3516 8082 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8076 3488 8953 3516
rect 8076 3476 8082 3488
rect 8680 3460 8708 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 8941 3479 8999 3485
rect 6822 3448 6828 3460
rect 6783 3420 6828 3448
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 8662 3408 8668 3460
rect 8720 3408 8726 3460
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 5261 3383 5319 3389
rect 5261 3380 5273 3383
rect 4764 3352 5273 3380
rect 4764 3340 4770 3352
rect 5261 3349 5273 3352
rect 5307 3380 5319 3383
rect 5626 3380 5632 3392
rect 5307 3352 5632 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 4706 3176 4712 3188
rect 4667 3148 4712 3176
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5166 3176 5172 3188
rect 5123 3148 5172 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7340 3148 7757 3176
rect 7340 3136 7346 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 8481 3179 8539 3185
rect 8481 3145 8493 3179
rect 8527 3176 8539 3179
rect 8754 3176 8760 3188
rect 8527 3148 8760 3176
rect 8527 3145 8539 3148
rect 8481 3139 8539 3145
rect 8754 3136 8760 3148
rect 8812 3176 8818 3188
rect 9766 3176 9772 3188
rect 8812 3148 9772 3176
rect 8812 3136 8818 3148
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 10652 3148 10701 3176
rect 10652 3136 10658 3148
rect 10689 3145 10701 3148
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 1762 3068 1768 3120
rect 1820 3108 1826 3120
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 1820 3080 6561 3108
rect 1820 3068 1826 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 5905 3043 5963 3049
rect 5905 3009 5917 3043
rect 5951 3040 5963 3043
rect 6178 3040 6184 3052
rect 5951 3012 6184 3040
rect 5951 3009 5963 3012
rect 5905 3003 5963 3009
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 5261 2975 5319 2981
rect 5261 2972 5273 2975
rect 5132 2944 5273 2972
rect 5132 2932 5138 2944
rect 5261 2941 5273 2944
rect 5307 2972 5319 2975
rect 5718 2972 5724 2984
rect 5307 2944 5724 2972
rect 5307 2941 5319 2944
rect 5261 2935 5319 2941
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 6564 2972 6592 3071
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8662 3040 8668 3052
rect 8623 3012 8668 3040
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 9306 3040 9312 3052
rect 9267 3012 9312 3040
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 7926 2972 7932 2984
rect 6564 2944 7932 2972
rect 6638 2904 6644 2916
rect 6196 2876 6644 2904
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 6196 2845 6224 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 7161 2913 7189 2944
rect 7926 2932 7932 2944
rect 7984 2972 7990 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 7984 2944 8033 2972
rect 7984 2932 7990 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10594 2972 10600 2984
rect 10183 2944 10600 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 13446 2972 13452 2984
rect 13407 2944 13452 2972
rect 13446 2932 13452 2944
rect 13504 2972 13510 2984
rect 13504 2944 14136 2972
rect 13504 2932 13510 2944
rect 7146 2907 7204 2913
rect 7146 2873 7158 2907
rect 7192 2873 7204 2907
rect 7146 2867 7204 2873
rect 8754 2864 8760 2916
rect 8812 2904 8818 2916
rect 8812 2876 8857 2904
rect 8812 2864 8818 2876
rect 14108 2848 14136 2944
rect 6181 2839 6239 2845
rect 6181 2836 6193 2839
rect 2924 2808 6193 2836
rect 2924 2796 2930 2808
rect 6181 2805 6193 2808
rect 6227 2805 6239 2839
rect 6181 2799 6239 2805
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 10321 2839 10379 2845
rect 10321 2836 10333 2839
rect 10008 2808 10333 2836
rect 10008 2796 10014 2808
rect 10321 2805 10333 2808
rect 10367 2805 10379 2839
rect 10321 2799 10379 2805
rect 13633 2839 13691 2845
rect 13633 2805 13645 2839
rect 13679 2836 13691 2839
rect 13906 2836 13912 2848
rect 13679 2808 13912 2836
rect 13679 2805 13691 2808
rect 13633 2799 13691 2805
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14090 2836 14096 2848
rect 14051 2808 14096 2836
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 6178 2632 6184 2644
rect 5675 2604 6184 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 6822 2592 6828 2644
rect 6880 2632 6886 2644
rect 7101 2635 7159 2641
rect 7101 2632 7113 2635
rect 6880 2604 7113 2632
rect 6880 2592 6886 2604
rect 7101 2601 7113 2604
rect 7147 2601 7159 2635
rect 8846 2632 8852 2644
rect 8807 2604 8852 2632
rect 7101 2595 7159 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 4890 2564 4896 2576
rect 4851 2536 4896 2564
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 7653 2567 7711 2573
rect 7653 2533 7665 2567
rect 7699 2564 7711 2567
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 7699 2536 7941 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 7929 2533 7941 2536
rect 7975 2564 7987 2567
rect 8110 2564 8116 2576
rect 7975 2536 8116 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 8481 2567 8539 2573
rect 8481 2533 8493 2567
rect 8527 2564 8539 2567
rect 8662 2564 8668 2576
rect 8527 2536 8668 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4126 2468 4261 2496
rect 842 2252 848 2304
rect 900 2292 906 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 900 2264 3801 2292
rect 900 2252 906 2264
rect 3789 2261 3801 2264
rect 3835 2292 3847 2295
rect 4126 2292 4154 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 4249 2459 4307 2465
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 5902 2496 5908 2508
rect 5767 2468 5908 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 5902 2456 5908 2468
rect 5960 2496 5966 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5960 2468 6285 2496
rect 5960 2456 5966 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10042 2496 10048 2508
rect 9815 2468 10048 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10042 2456 10048 2468
rect 10100 2496 10106 2508
rect 10100 2468 10456 2496
rect 10100 2456 10106 2468
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8846 2428 8852 2440
rect 7883 2400 8852 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 5905 2363 5963 2369
rect 5905 2329 5917 2363
rect 5951 2360 5963 2363
rect 8018 2360 8024 2372
rect 5951 2332 8024 2360
rect 5951 2329 5963 2332
rect 5905 2323 5963 2329
rect 8018 2320 8024 2332
rect 8076 2320 8082 2372
rect 3835 2264 4154 2292
rect 3835 2261 3847 2264
rect 3789 2255 3847 2261
rect 5074 2252 5080 2304
rect 5132 2292 5138 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 5132 2264 5181 2292
rect 5132 2252 5138 2264
rect 5169 2261 5181 2264
rect 5215 2261 5227 2295
rect 5169 2255 5227 2261
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 10428 2301 10456 2468
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 10928 2468 13461 2496
rect 10928 2456 10934 2468
rect 13449 2465 13461 2468
rect 13495 2496 13507 2499
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13495 2468 14013 2496
rect 13495 2465 13507 2468
rect 13449 2459 13507 2465
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 14001 2459 14059 2465
rect 13633 2363 13691 2369
rect 13633 2329 13645 2363
rect 13679 2360 13691 2363
rect 15194 2360 15200 2372
rect 13679 2332 15200 2360
rect 13679 2329 13691 2332
rect 13633 2323 13691 2329
rect 15194 2320 15200 2332
rect 15252 2320 15258 2372
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 8904 2264 9965 2292
rect 8904 2252 8910 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 10413 2295 10471 2301
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 12894 2292 12900 2304
rect 10459 2264 12900 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 3418 76 3424 128
rect 3476 116 3482 128
rect 6822 116 6828 128
rect 3476 88 6828 116
rect 3476 76 3482 88
rect 6822 76 6828 88
rect 6880 76 6886 128
rect 11146 76 11152 128
rect 11204 116 11210 128
rect 12066 116 12072 128
rect 11204 88 12072 116
rect 11204 76 11210 88
rect 12066 76 12072 88
rect 12124 76 12130 128
<< via1 >>
rect 6644 39652 6696 39704
rect 9312 39652 9364 39704
rect 9864 39652 9916 39704
rect 13728 39652 13780 39704
rect 20 39584 72 39636
rect 664 39584 716 39636
rect 1492 39584 1544 39636
rect 2044 39584 2096 39636
rect 5632 39584 5684 39636
rect 6460 39584 6512 39636
rect 7104 39584 7156 39636
rect 7932 39584 7984 39636
rect 9772 39584 9824 39636
rect 10784 39584 10836 39636
rect 13820 39584 13872 39636
rect 15200 39584 15252 39636
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 1584 34663 1636 34672
rect 1584 34629 1593 34663
rect 1593 34629 1627 34663
rect 1627 34629 1636 34663
rect 1584 34620 1636 34629
rect 3148 34688 3200 34740
rect 11980 34688 12032 34740
rect 8024 34552 8076 34604
rect 9496 34484 9548 34536
rect 8852 34348 8904 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 5356 29835 5408 29844
rect 5356 29801 5365 29835
rect 5365 29801 5399 29835
rect 5399 29801 5408 29835
rect 5356 29792 5408 29801
rect 5172 29699 5224 29708
rect 5172 29665 5181 29699
rect 5181 29665 5215 29699
rect 5215 29665 5224 29699
rect 5172 29656 5224 29665
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 4068 28976 4120 29028
rect 5172 29019 5224 29028
rect 5172 28985 5181 29019
rect 5181 28985 5215 29019
rect 5215 28985 5224 29019
rect 5172 28976 5224 28985
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 13636 28747 13688 28756
rect 13636 28713 13645 28747
rect 13645 28713 13679 28747
rect 13679 28713 13688 28747
rect 13636 28704 13688 28713
rect 13452 28611 13504 28620
rect 13452 28577 13461 28611
rect 13461 28577 13495 28611
rect 13495 28577 13504 28611
rect 13452 28568 13504 28577
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 11336 27820 11388 27872
rect 13452 27863 13504 27872
rect 13452 27829 13461 27863
rect 13461 27829 13495 27863
rect 13495 27829 13504 27863
rect 13452 27820 13504 27829
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 4620 26571 4672 26580
rect 4620 26537 4629 26571
rect 4629 26537 4663 26571
rect 4663 26537 4672 26571
rect 4620 26528 4672 26537
rect 4436 26435 4488 26444
rect 4436 26401 4445 26435
rect 4445 26401 4479 26435
rect 4479 26401 4488 26435
rect 4436 26392 4488 26401
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4436 25644 4488 25696
rect 6000 25644 6052 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 112 22040 164 22092
rect 1584 22040 1636 22092
rect 112 21836 164 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 6644 19864 6696 19916
rect 6736 19660 6788 19712
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 5172 19252 5224 19304
rect 1400 19184 1452 19236
rect 6644 19456 6696 19508
rect 7012 19320 7064 19372
rect 6920 19227 6972 19236
rect 6920 19193 6929 19227
rect 6929 19193 6963 19227
rect 6963 19193 6972 19227
rect 6920 19184 6972 19193
rect 5172 19116 5224 19168
rect 6828 19116 6880 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 9772 18912 9824 18964
rect 6092 18844 6144 18896
rect 6828 18887 6880 18896
rect 6828 18853 6837 18887
rect 6837 18853 6871 18887
rect 6871 18853 6880 18887
rect 6828 18844 6880 18853
rect 7472 18844 7524 18896
rect 5172 18776 5224 18828
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 7012 18708 7064 18760
rect 6644 18640 6696 18692
rect 8024 18683 8076 18692
rect 8024 18649 8033 18683
rect 8033 18649 8067 18683
rect 8067 18649 8076 18683
rect 8024 18640 8076 18649
rect 5080 18572 5132 18624
rect 5356 18615 5408 18624
rect 5356 18581 5365 18615
rect 5365 18581 5399 18615
rect 5399 18581 5408 18615
rect 5356 18572 5408 18581
rect 5724 18615 5776 18624
rect 5724 18581 5733 18615
rect 5733 18581 5767 18615
rect 5767 18581 5776 18615
rect 5724 18572 5776 18581
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 6920 18368 6972 18420
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 7840 18300 7892 18352
rect 5724 18232 5776 18284
rect 6828 18232 6880 18284
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 8024 18232 8076 18241
rect 9312 18164 9364 18216
rect 5356 18139 5408 18148
rect 5356 18105 5365 18139
rect 5365 18105 5399 18139
rect 5399 18105 5408 18139
rect 5908 18139 5960 18148
rect 5356 18096 5408 18105
rect 5908 18105 5917 18139
rect 5917 18105 5951 18139
rect 5951 18105 5960 18139
rect 7012 18139 7064 18148
rect 5908 18096 5960 18105
rect 7012 18105 7021 18139
rect 7021 18105 7055 18139
rect 7055 18105 7064 18139
rect 7012 18096 7064 18105
rect 5172 18028 5224 18080
rect 6092 18028 6144 18080
rect 6644 18071 6696 18080
rect 6644 18037 6653 18071
rect 6653 18037 6687 18071
rect 6687 18037 6696 18071
rect 6644 18028 6696 18037
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 7564 18028 7616 18080
rect 7748 18139 7800 18148
rect 7748 18105 7757 18139
rect 7757 18105 7791 18139
rect 7791 18105 7800 18139
rect 7748 18096 7800 18105
rect 7840 18028 7892 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 5080 17824 5132 17876
rect 6828 17824 6880 17876
rect 5264 17756 5316 17808
rect 5356 17756 5408 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2964 17688 3016 17740
rect 3516 17688 3568 17740
rect 4068 17688 4120 17740
rect 9680 17688 9732 17740
rect 11428 17731 11480 17740
rect 11428 17697 11437 17731
rect 11437 17697 11471 17731
rect 11471 17697 11480 17731
rect 11428 17688 11480 17697
rect 4804 17620 4856 17672
rect 6736 17620 6788 17672
rect 1584 17595 1636 17604
rect 1584 17561 1593 17595
rect 1593 17561 1627 17595
rect 1627 17561 1636 17595
rect 1584 17552 1636 17561
rect 6184 17552 6236 17604
rect 7564 17620 7616 17672
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 7656 17527 7708 17536
rect 7656 17493 7665 17527
rect 7665 17493 7699 17527
rect 7699 17493 7708 17527
rect 7656 17484 7708 17493
rect 11980 17484 12032 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 1400 17280 1452 17332
rect 2964 17323 3016 17332
rect 2964 17289 2973 17323
rect 2973 17289 3007 17323
rect 3007 17289 3016 17323
rect 2964 17280 3016 17289
rect 5356 17280 5408 17332
rect 6184 17323 6236 17332
rect 6184 17289 6193 17323
rect 6193 17289 6227 17323
rect 6227 17289 6236 17323
rect 6184 17280 6236 17289
rect 7472 17280 7524 17332
rect 8116 17280 8168 17332
rect 11428 17323 11480 17332
rect 6644 17212 6696 17264
rect 6736 17212 6788 17264
rect 5080 17144 5132 17196
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 11428 17289 11437 17323
rect 11437 17289 11471 17323
rect 11471 17289 11480 17323
rect 11428 17280 11480 17289
rect 9312 17187 9364 17196
rect 9312 17153 9321 17187
rect 9321 17153 9355 17187
rect 9355 17153 9364 17187
rect 9312 17144 9364 17153
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 5264 17008 5316 17060
rect 8760 17051 8812 17060
rect 8760 17017 8769 17051
rect 8769 17017 8803 17051
rect 8803 17017 8812 17051
rect 8760 17008 8812 17017
rect 5632 16940 5684 16992
rect 7196 16983 7248 16992
rect 7196 16949 7205 16983
rect 7205 16949 7239 16983
rect 7239 16949 7248 16983
rect 7196 16940 7248 16949
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 10876 16940 10928 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 4804 16779 4856 16788
rect 4804 16745 4813 16779
rect 4813 16745 4847 16779
rect 4847 16745 4856 16779
rect 4804 16736 4856 16745
rect 6184 16736 6236 16788
rect 7656 16736 7708 16788
rect 5540 16668 5592 16720
rect 7196 16668 7248 16720
rect 5172 16600 5224 16652
rect 10600 16600 10652 16652
rect 4528 16532 4580 16584
rect 6644 16532 6696 16584
rect 5264 16439 5316 16448
rect 5264 16405 5273 16439
rect 5273 16405 5307 16439
rect 5307 16405 5316 16439
rect 5264 16396 5316 16405
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 8208 16396 8260 16448
rect 8760 16396 8812 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 6092 16192 6144 16244
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 5632 16056 5684 16108
rect 6092 16056 6144 16108
rect 4712 15988 4764 16040
rect 7472 15988 7524 16040
rect 5540 15920 5592 15972
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 5264 15648 5316 15700
rect 5540 15580 5592 15632
rect 5908 15444 5960 15496
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 4712 15308 4764 15360
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 7472 15351 7524 15360
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 8852 15011 8904 15020
rect 8852 14977 8861 15011
rect 8861 14977 8895 15011
rect 8895 14977 8904 15011
rect 8852 14968 8904 14977
rect 8668 14875 8720 14884
rect 8668 14841 8677 14875
rect 8677 14841 8711 14875
rect 8711 14841 8720 14875
rect 8668 14832 8720 14841
rect 5908 14807 5960 14816
rect 5908 14773 5917 14807
rect 5917 14773 5951 14807
rect 5951 14773 5960 14807
rect 5908 14764 5960 14773
rect 6920 14764 6972 14816
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 7196 14492 7248 14544
rect 9772 14492 9824 14544
rect 8668 14424 8720 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 8208 14356 8260 14408
rect 11244 14356 11296 14408
rect 8852 14288 8904 14340
rect 12164 14288 12216 14340
rect 7012 14220 7064 14272
rect 8024 14220 8076 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 8208 13991 8260 14000
rect 8208 13957 8217 13991
rect 8217 13957 8251 13991
rect 8251 13957 8260 13991
rect 8208 13948 8260 13957
rect 9956 13948 10008 14000
rect 10048 13880 10100 13932
rect 10232 13923 10284 13932
rect 10232 13889 10241 13923
rect 10241 13889 10275 13923
rect 10275 13889 10284 13923
rect 10232 13880 10284 13889
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 7012 13812 7064 13864
rect 7288 13855 7340 13864
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 7656 13812 7708 13864
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 9956 13787 10008 13796
rect 9956 13753 9965 13787
rect 9965 13753 9999 13787
rect 9999 13753 10008 13787
rect 9956 13744 10008 13753
rect 10048 13787 10100 13796
rect 10048 13753 10057 13787
rect 10057 13753 10091 13787
rect 10091 13753 10100 13787
rect 10048 13744 10100 13753
rect 7012 13676 7064 13728
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 9404 13719 9456 13728
rect 9404 13685 9413 13719
rect 9413 13685 9447 13719
rect 9447 13685 9456 13719
rect 9404 13676 9456 13685
rect 9680 13676 9732 13728
rect 11060 13744 11112 13796
rect 13452 13787 13504 13796
rect 13452 13753 13461 13787
rect 13461 13753 13495 13787
rect 13495 13753 13504 13787
rect 13452 13744 13504 13753
rect 12256 13676 12308 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 20 13472 72 13524
rect 10048 13515 10100 13524
rect 10048 13481 10057 13515
rect 10057 13481 10091 13515
rect 10091 13481 10100 13515
rect 10048 13472 10100 13481
rect 6184 13404 6236 13456
rect 7656 13404 7708 13456
rect 11704 13404 11756 13456
rect 12164 13447 12216 13456
rect 12164 13413 12173 13447
rect 12173 13413 12207 13447
rect 12207 13413 12216 13447
rect 12164 13404 12216 13413
rect 5172 13336 5224 13388
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 7288 13336 7340 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 10232 13336 10284 13388
rect 10692 13268 10744 13320
rect 12164 13268 12216 13320
rect 6736 13132 6788 13184
rect 8024 13132 8076 13184
rect 9312 13132 9364 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 10692 12971 10744 12980
rect 10692 12937 10701 12971
rect 10701 12937 10735 12971
rect 10735 12937 10744 12971
rect 10692 12928 10744 12937
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 12256 12928 12308 12980
rect 4160 12792 4212 12844
rect 5080 12792 5132 12844
rect 8392 12792 8444 12844
rect 11060 12792 11112 12844
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5172 12767 5224 12776
rect 5172 12733 5181 12767
rect 5181 12733 5215 12767
rect 5215 12733 5224 12767
rect 5172 12724 5224 12733
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 4344 12631 4396 12640
rect 4344 12597 4353 12631
rect 4353 12597 4387 12631
rect 4387 12597 4396 12631
rect 4344 12588 4396 12597
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 7012 12724 7064 12776
rect 7656 12767 7708 12776
rect 6736 12656 6788 12708
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 9312 12724 9364 12776
rect 10784 12724 10836 12776
rect 13728 12792 13780 12844
rect 14740 12792 14792 12844
rect 12072 12724 12124 12776
rect 13452 12724 13504 12776
rect 6184 12588 6236 12597
rect 7472 12588 7524 12640
rect 8668 12588 8720 12640
rect 10048 12588 10100 12640
rect 11244 12588 11296 12640
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 6644 12384 6696 12436
rect 7656 12384 7708 12436
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5172 12248 5224 12257
rect 5724 12248 5776 12300
rect 6184 12248 6236 12300
rect 6644 12291 6696 12300
rect 6644 12257 6653 12291
rect 6653 12257 6687 12291
rect 6687 12257 6696 12291
rect 6644 12248 6696 12257
rect 7564 12316 7616 12368
rect 8300 12316 8352 12368
rect 9404 12384 9456 12436
rect 10784 12384 10836 12436
rect 13636 12427 13688 12436
rect 13636 12393 13645 12427
rect 13645 12393 13679 12427
rect 13679 12393 13688 12427
rect 13636 12384 13688 12393
rect 9496 12316 9548 12368
rect 10048 12316 10100 12368
rect 11244 12316 11296 12368
rect 11612 12359 11664 12368
rect 11612 12325 11621 12359
rect 11621 12325 11655 12359
rect 11655 12325 11664 12359
rect 11612 12316 11664 12325
rect 7196 12180 7248 12232
rect 4160 12112 4212 12164
rect 5632 12112 5684 12164
rect 7012 12112 7064 12164
rect 8392 12248 8444 12300
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 10784 12180 10836 12232
rect 9772 12112 9824 12164
rect 11152 12112 11204 12164
rect 12072 12155 12124 12164
rect 12072 12121 12081 12155
rect 12081 12121 12115 12155
rect 12115 12121 12124 12155
rect 12072 12112 12124 12121
rect 4620 12044 4672 12096
rect 5172 12044 5224 12096
rect 5724 12087 5776 12096
rect 5724 12053 5733 12087
rect 5733 12053 5767 12087
rect 5767 12053 5776 12087
rect 5724 12044 5776 12053
rect 7932 12087 7984 12096
rect 7932 12053 7941 12087
rect 7941 12053 7975 12087
rect 7975 12053 7984 12087
rect 7932 12044 7984 12053
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 9496 11840 9548 11892
rect 9956 11840 10008 11892
rect 11612 11883 11664 11892
rect 11612 11849 11621 11883
rect 11621 11849 11655 11883
rect 11655 11849 11664 11883
rect 11612 11840 11664 11849
rect 12624 11840 12676 11892
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 5172 11772 5224 11824
rect 7932 11772 7984 11824
rect 10324 11772 10376 11824
rect 5724 11704 5776 11756
rect 4436 11679 4488 11688
rect 4436 11645 4445 11679
rect 4445 11645 4479 11679
rect 4479 11645 4488 11679
rect 4436 11636 4488 11645
rect 5172 11679 5224 11688
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 4528 11543 4580 11552
rect 4528 11509 4537 11543
rect 4537 11509 4571 11543
rect 4571 11509 4580 11543
rect 4528 11500 4580 11509
rect 4620 11500 4672 11552
rect 8760 11704 8812 11756
rect 12164 11704 12216 11756
rect 7472 11636 7524 11688
rect 8024 11679 8076 11688
rect 8024 11645 8033 11679
rect 8033 11645 8067 11679
rect 8067 11645 8076 11679
rect 8024 11636 8076 11645
rect 8576 11636 8628 11688
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 7012 11568 7064 11620
rect 8668 11568 8720 11620
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 10324 11679 10376 11688
rect 9956 11636 10008 11645
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 8392 11500 8444 11552
rect 9312 11500 9364 11552
rect 12440 11500 12492 11552
rect 12624 11611 12676 11620
rect 12624 11577 12633 11611
rect 12633 11577 12667 11611
rect 12667 11577 12676 11611
rect 12624 11568 12676 11577
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 3608 11296 3660 11348
rect 4160 11296 4212 11348
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 5724 11296 5776 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 7196 11296 7248 11348
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 5172 11092 5224 11144
rect 6184 11160 6236 11212
rect 6736 11228 6788 11280
rect 7472 11271 7524 11280
rect 7472 11237 7481 11271
rect 7481 11237 7515 11271
rect 7515 11237 7524 11271
rect 7472 11228 7524 11237
rect 8852 11228 8904 11280
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 11796 11228 11848 11280
rect 7472 11092 7524 11144
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8760 11135 8812 11144
rect 8760 11101 8769 11135
rect 8769 11101 8803 11135
rect 8803 11101 8812 11135
rect 8760 11092 8812 11101
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 11520 11135 11572 11144
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 7196 11024 7248 11076
rect 10416 11024 10468 11076
rect 12072 11024 12124 11076
rect 8024 10956 8076 11008
rect 10784 10956 10836 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 6184 10752 6236 10804
rect 6644 10752 6696 10804
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 11520 10752 11572 10804
rect 7932 10684 7984 10736
rect 8576 10684 8628 10736
rect 11796 10727 11848 10736
rect 11796 10693 11805 10727
rect 11805 10693 11839 10727
rect 11839 10693 11848 10727
rect 11796 10684 11848 10693
rect 4436 10616 4488 10668
rect 9680 10616 9732 10668
rect 4620 10548 4672 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 7472 10480 7524 10532
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 8024 10548 8076 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 8576 10480 8628 10532
rect 10048 10480 10100 10532
rect 4252 10412 4304 10421
rect 7748 10412 7800 10464
rect 8300 10412 8352 10464
rect 13452 10412 13504 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 5632 10251 5684 10260
rect 5632 10217 5641 10251
rect 5641 10217 5675 10251
rect 5675 10217 5684 10251
rect 5632 10208 5684 10217
rect 8668 10208 8720 10260
rect 8852 10251 8904 10260
rect 8852 10217 8861 10251
rect 8861 10217 8895 10251
rect 8895 10217 8904 10251
rect 8852 10208 8904 10217
rect 12440 10208 12492 10260
rect 9220 10183 9272 10192
rect 9220 10149 9229 10183
rect 9229 10149 9263 10183
rect 9263 10149 9272 10183
rect 9220 10140 9272 10149
rect 9772 10183 9824 10192
rect 9772 10149 9781 10183
rect 9781 10149 9815 10183
rect 9815 10149 9824 10183
rect 9772 10140 9824 10149
rect 10140 10140 10192 10192
rect 10416 10183 10468 10192
rect 10416 10149 10425 10183
rect 10425 10149 10459 10183
rect 10459 10149 10468 10183
rect 10416 10140 10468 10149
rect 5632 10072 5684 10124
rect 6828 10072 6880 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 7748 10072 7800 10124
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 11336 10072 11388 10124
rect 4160 9868 4212 9920
rect 4528 9868 4580 9920
rect 7012 9868 7064 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 5632 9707 5684 9716
rect 5632 9673 5641 9707
rect 5641 9673 5675 9707
rect 5675 9673 5684 9707
rect 5632 9664 5684 9673
rect 8668 9664 8720 9716
rect 10140 9664 10192 9716
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 7656 9596 7708 9648
rect 8116 9596 8168 9648
rect 10784 9528 10836 9580
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7656 9460 7708 9512
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 9496 9503 9548 9512
rect 9496 9469 9514 9503
rect 9514 9469 9548 9503
rect 9496 9460 9548 9469
rect 8668 9392 8720 9444
rect 10692 9460 10744 9512
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 7104 9324 7156 9376
rect 9680 9324 9732 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 12072 9324 12124 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 5908 9120 5960 9172
rect 8024 9120 8076 9172
rect 8116 9120 8168 9172
rect 9772 9120 9824 9172
rect 11428 9120 11480 9172
rect 13820 9120 13872 9172
rect 8668 9052 8720 9104
rect 5264 8984 5316 9036
rect 7012 8984 7064 9036
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 10324 9027 10376 9036
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 11520 9027 11572 9036
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 5724 8916 5776 8968
rect 7288 8916 7340 8968
rect 7748 8959 7800 8968
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 8484 8848 8536 8900
rect 10508 8848 10560 8900
rect 12624 8848 12676 8900
rect 5908 8823 5960 8832
rect 5908 8789 5917 8823
rect 5917 8789 5951 8823
rect 5951 8789 5960 8823
rect 5908 8780 5960 8789
rect 9956 8823 10008 8832
rect 9956 8789 9965 8823
rect 9965 8789 9999 8823
rect 9999 8789 10008 8823
rect 9956 8780 10008 8789
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 9956 8576 10008 8628
rect 10324 8576 10376 8628
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 4896 8508 4948 8560
rect 5448 8551 5500 8560
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 5080 8440 5132 8492
rect 5816 8440 5868 8492
rect 7656 8440 7708 8492
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 8668 8440 8720 8492
rect 5724 8372 5776 8424
rect 6644 8372 6696 8424
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 13728 8372 13780 8424
rect 5172 8347 5224 8356
rect 5172 8313 5181 8347
rect 5181 8313 5215 8347
rect 5215 8313 5224 8347
rect 5172 8304 5224 8313
rect 5264 8304 5316 8356
rect 5448 8304 5500 8356
rect 5908 8304 5960 8356
rect 8208 8304 8260 8356
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 7012 8236 7064 8288
rect 8300 8279 8352 8288
rect 8300 8245 8309 8279
rect 8309 8245 8343 8279
rect 8343 8245 8352 8279
rect 8300 8236 8352 8245
rect 9956 8236 10008 8288
rect 10416 8304 10468 8356
rect 12624 8304 12676 8356
rect 11060 8236 11112 8288
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 4528 8075 4580 8084
rect 4528 8041 4537 8075
rect 4537 8041 4571 8075
rect 4571 8041 4580 8075
rect 4528 8032 4580 8041
rect 7656 8032 7708 8084
rect 7932 7964 7984 8016
rect 9772 7964 9824 8016
rect 10324 8032 10376 8084
rect 10416 8007 10468 8016
rect 10416 7973 10425 8007
rect 10425 7973 10459 8007
rect 10459 7973 10468 8007
rect 10416 7964 10468 7973
rect 11520 7964 11572 8016
rect 5264 7896 5316 7948
rect 5632 7828 5684 7880
rect 5908 7828 5960 7880
rect 7288 7760 7340 7812
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 5356 7692 5408 7744
rect 6552 7692 6604 7744
rect 7656 7735 7708 7744
rect 7656 7701 7665 7735
rect 7665 7701 7699 7735
rect 7699 7701 7708 7735
rect 8668 7828 8720 7880
rect 11796 7828 11848 7880
rect 11060 7760 11112 7812
rect 7656 7692 7708 7701
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 5724 7488 5776 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 4804 7420 4856 7472
rect 6644 7420 6696 7472
rect 7380 7420 7432 7472
rect 7656 7352 7708 7404
rect 8208 7352 8260 7404
rect 9036 7352 9088 7404
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 3700 7284 3752 7336
rect 5264 7284 5316 7336
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 12900 7327 12952 7336
rect 5816 7216 5868 7268
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 5448 7148 5500 7200
rect 5908 7148 5960 7200
rect 7104 7259 7156 7268
rect 7104 7225 7113 7259
rect 7113 7225 7147 7259
rect 7147 7225 7156 7259
rect 7104 7216 7156 7225
rect 8668 7216 8720 7268
rect 7380 7148 7432 7200
rect 7932 7191 7984 7200
rect 7932 7157 7941 7191
rect 7941 7157 7975 7191
rect 7975 7157 7984 7191
rect 7932 7148 7984 7157
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 10416 7259 10468 7268
rect 10416 7225 10425 7259
rect 10425 7225 10459 7259
rect 10459 7225 10468 7259
rect 10416 7216 10468 7225
rect 11336 7148 11388 7200
rect 11520 7148 11572 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 3700 6987 3752 6996
rect 3700 6953 3709 6987
rect 3709 6953 3743 6987
rect 3743 6953 3752 6987
rect 3700 6944 3752 6953
rect 5724 6944 5776 6996
rect 7104 6944 7156 6996
rect 7380 6987 7432 6996
rect 7380 6953 7389 6987
rect 7389 6953 7423 6987
rect 7423 6953 7432 6987
rect 7380 6944 7432 6953
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 9036 6987 9088 6996
rect 9036 6953 9045 6987
rect 9045 6953 9079 6987
rect 9079 6953 9088 6987
rect 9036 6944 9088 6953
rect 11520 6987 11572 6996
rect 11520 6953 11529 6987
rect 11529 6953 11563 6987
rect 11563 6953 11572 6987
rect 11520 6944 11572 6953
rect 6184 6919 6236 6928
rect 6184 6885 6193 6919
rect 6193 6885 6227 6919
rect 6227 6885 6236 6919
rect 6184 6876 6236 6885
rect 7932 6876 7984 6928
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 5356 6808 5408 6860
rect 9956 6876 10008 6928
rect 10416 6919 10468 6928
rect 10416 6885 10425 6919
rect 10425 6885 10459 6919
rect 10459 6885 10468 6919
rect 10416 6876 10468 6885
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 5448 6672 5500 6724
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8668 6740 8720 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 5908 6672 5960 6724
rect 5172 6604 5224 6656
rect 5264 6604 5316 6656
rect 5724 6647 5776 6656
rect 5724 6613 5733 6647
rect 5733 6613 5767 6647
rect 5767 6613 5776 6647
rect 5724 6604 5776 6613
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 5724 6400 5776 6452
rect 7104 6400 7156 6452
rect 8116 6400 8168 6452
rect 9772 6400 9824 6452
rect 11336 6400 11388 6452
rect 5356 6332 5408 6384
rect 10416 6375 10468 6384
rect 10416 6341 10425 6375
rect 10425 6341 10459 6375
rect 10459 6341 10468 6375
rect 10416 6332 10468 6341
rect 10508 6332 10560 6384
rect 4896 6264 4948 6316
rect 7748 6264 7800 6316
rect 9956 6264 10008 6316
rect 10324 6264 10376 6316
rect 4436 6128 4488 6180
rect 4988 6128 5040 6180
rect 5908 6196 5960 6248
rect 7840 6196 7892 6248
rect 10600 6196 10652 6248
rect 12256 6196 12308 6248
rect 7932 6128 7984 6180
rect 9864 6171 9916 6180
rect 9864 6137 9873 6171
rect 9873 6137 9907 6171
rect 9907 6137 9916 6171
rect 9864 6128 9916 6137
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 9680 6103 9732 6112
rect 9680 6069 9689 6103
rect 9689 6069 9723 6103
rect 9723 6069 9732 6103
rect 9680 6060 9732 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 4804 5856 4856 5908
rect 6736 5856 6788 5908
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 9864 5856 9916 5908
rect 9680 5831 9732 5840
rect 9680 5797 9689 5831
rect 9689 5797 9723 5831
rect 9723 5797 9732 5831
rect 9680 5788 9732 5797
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 4988 5720 5040 5772
rect 6644 5720 6696 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 7932 5516 7984 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 5172 5312 5224 5364
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 8116 5312 8168 5364
rect 9864 5312 9916 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 5908 5108 5960 5160
rect 6092 5108 6144 5160
rect 6644 5040 6696 5092
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 7288 5108 7340 5160
rect 8392 5040 8444 5092
rect 6092 4972 6144 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 6092 4768 6144 4820
rect 7104 4768 7156 4820
rect 9772 4768 9824 4820
rect 112 4632 164 4684
rect 5172 4632 5224 4684
rect 5448 4632 5500 4684
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 9956 4632 10008 4684
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 5356 4471 5408 4480
rect 5356 4437 5365 4471
rect 5365 4437 5399 4471
rect 5399 4437 5408 4471
rect 5356 4428 5408 4437
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 6184 4224 6236 4276
rect 8484 4224 8536 4276
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 7104 4131 7156 4140
rect 7104 4097 7113 4131
rect 7113 4097 7147 4131
rect 7147 4097 7156 4131
rect 7104 4088 7156 4097
rect 3516 4020 3568 4072
rect 5080 4020 5132 4072
rect 10600 4088 10652 4140
rect 4896 3952 4948 4004
rect 5356 3995 5408 4004
rect 5356 3961 5365 3995
rect 5365 3961 5399 3995
rect 5399 3961 5408 3995
rect 5356 3952 5408 3961
rect 6368 3952 6420 4004
rect 5632 3927 5684 3936
rect 5632 3893 5641 3927
rect 5641 3893 5675 3927
rect 5675 3893 5684 3927
rect 8024 3952 8076 4004
rect 8668 3995 8720 4004
rect 8668 3961 8677 3995
rect 8677 3961 8711 3995
rect 8711 3961 8720 3995
rect 8668 3952 8720 3961
rect 8760 3995 8812 4004
rect 8760 3961 8769 3995
rect 8769 3961 8803 3995
rect 8803 3961 8812 3995
rect 9312 3995 9364 4004
rect 8760 3952 8812 3961
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9956 3995 10008 4004
rect 9312 3952 9364 3961
rect 9956 3961 9965 3995
rect 9965 3961 9999 3995
rect 9999 3961 10008 3995
rect 9956 3952 10008 3961
rect 5632 3884 5684 3893
rect 7288 3884 7340 3936
rect 8392 3884 8444 3936
rect 8852 3884 8904 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 7012 3680 7064 3732
rect 5632 3612 5684 3664
rect 7288 3655 7340 3664
rect 5172 3544 5224 3596
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 7288 3621 7297 3655
rect 7297 3621 7331 3655
rect 7331 3621 7340 3655
rect 7288 3612 7340 3621
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 8668 3680 8720 3732
rect 7932 3612 7984 3664
rect 8760 3612 8812 3664
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 8024 3476 8076 3528
rect 6828 3451 6880 3460
rect 6828 3417 6837 3451
rect 6837 3417 6871 3451
rect 6871 3417 6880 3451
rect 6828 3408 6880 3417
rect 8668 3408 8720 3460
rect 4712 3340 4764 3392
rect 5632 3340 5684 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 4712 3179 4764 3188
rect 4712 3145 4721 3179
rect 4721 3145 4755 3179
rect 4755 3145 4764 3179
rect 4712 3136 4764 3145
rect 5172 3136 5224 3188
rect 7288 3136 7340 3188
rect 8760 3136 8812 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10600 3136 10652 3188
rect 1768 3068 1820 3120
rect 6184 3000 6236 3052
rect 5080 2932 5132 2984
rect 5724 2932 5776 2984
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 2872 2796 2924 2848
rect 6644 2864 6696 2916
rect 7932 2932 7984 2984
rect 10600 2932 10652 2984
rect 13452 2975 13504 2984
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 9956 2796 10008 2848
rect 13912 2796 13964 2848
rect 14096 2839 14148 2848
rect 14096 2805 14105 2839
rect 14105 2805 14139 2839
rect 14139 2805 14148 2839
rect 14096 2796 14148 2805
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 6184 2592 6236 2644
rect 6828 2592 6880 2644
rect 8852 2635 8904 2644
rect 8852 2601 8861 2635
rect 8861 2601 8895 2635
rect 8895 2601 8904 2635
rect 8852 2592 8904 2601
rect 4896 2567 4948 2576
rect 4896 2533 4905 2567
rect 4905 2533 4939 2567
rect 4939 2533 4948 2567
rect 4896 2524 4948 2533
rect 8116 2524 8168 2576
rect 8668 2524 8720 2576
rect 848 2252 900 2304
rect 5908 2456 5960 2508
rect 10048 2456 10100 2508
rect 8852 2388 8904 2440
rect 8024 2320 8076 2372
rect 5080 2252 5132 2304
rect 8852 2252 8904 2304
rect 10876 2456 10928 2508
rect 15200 2320 15252 2372
rect 12900 2252 12952 2304
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 3424 76 3476 128
rect 6828 76 6880 128
rect 11152 76 11204 128
rect 12072 76 12124 128
<< metal2 >>
rect 20 39636 72 39642
rect 20 39578 72 39584
rect 662 39636 718 40000
rect 662 39584 664 39636
rect 716 39584 718 39636
rect 32 13530 60 39578
rect 662 39520 718 39584
rect 1492 39636 1544 39642
rect 1492 39578 1544 39584
rect 2042 39636 2098 40000
rect 3514 39658 3570 40000
rect 2042 39584 2044 39636
rect 2096 39584 2098 39636
rect 110 24984 166 24993
rect 110 24919 166 24928
rect 124 22098 152 24919
rect 112 22092 164 22098
rect 112 22034 164 22040
rect 112 21888 164 21894
rect 112 21830 164 21836
rect 124 21729 152 21830
rect 110 21720 166 21729
rect 110 21655 166 21664
rect 1400 19236 1452 19242
rect 1400 19178 1452 19184
rect 1412 17746 1440 19178
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1412 17338 1440 17682
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1504 17105 1532 39578
rect 2042 39520 2098 39584
rect 3160 39630 3570 39658
rect 1582 34776 1638 34785
rect 3160 34746 3188 39630
rect 3514 39520 3570 39630
rect 4986 39658 5042 40000
rect 4986 39630 5304 39658
rect 4986 39520 5042 39630
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 1582 34711 1638 34720
rect 3148 34740 3200 34746
rect 1596 34678 1624 34711
rect 3148 34682 3200 34688
rect 1584 34672 1636 34678
rect 1584 34614 1636 34620
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 5172 29708 5224 29714
rect 5172 29650 5224 29656
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 5184 29034 5212 29650
rect 4068 29028 4120 29034
rect 4068 28970 4120 28976
rect 5172 29028 5224 29034
rect 5172 28970 5224 28976
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 1596 21690 1624 22034
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1596 17610 1624 17847
rect 4080 17746 4108 28970
rect 4618 27840 4674 27849
rect 4618 27775 4674 27784
rect 4632 26586 4660 27775
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4436 26444 4488 26450
rect 4436 26386 4488 26392
rect 4448 25702 4476 26386
rect 4436 25696 4488 25702
rect 4436 25638 4488 25644
rect 5276 19514 5304 39630
rect 5632 39636 5684 39642
rect 5632 39578 5684 39584
rect 6458 39636 6514 40000
rect 6644 39704 6696 39710
rect 6644 39646 6696 39652
rect 6458 39584 6460 39636
rect 6512 39584 6514 39636
rect 5354 31104 5410 31113
rect 5354 31039 5410 31048
rect 5368 29850 5396 31039
rect 5356 29844 5408 29850
rect 5356 29786 5408 29792
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 19174 5212 19246
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5184 18834 5212 19110
rect 5172 18828 5224 18834
rect 5172 18770 5224 18776
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 17882 5120 18566
rect 5184 18086 5212 18770
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18154 5396 18566
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 1584 17604 1636 17610
rect 1584 17546 1636 17552
rect 2976 17338 3004 17682
rect 2964 17332 3016 17338
rect 2964 17274 3016 17280
rect 1490 17096 1546 17105
rect 1490 17031 1546 17040
rect 20 13524 72 13530
rect 20 13466 72 13472
rect 110 4992 166 5001
rect 110 4927 166 4936
rect 124 4690 152 4927
rect 112 4684 164 4690
rect 112 4626 164 4632
rect 3528 4154 3556 17682
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 4816 16794 4844 17614
rect 5092 17202 5120 17818
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 5184 16658 5212 18022
rect 5368 17814 5396 18090
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5276 17066 5304 17750
rect 5368 17338 5396 17750
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5264 17060 5316 17066
rect 5264 17002 5316 17008
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 4540 15910 4568 16526
rect 5276 16454 5304 17002
rect 5644 16998 5672 39578
rect 6458 39520 6514 39584
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 18290 5764 18566
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 5920 17202 5948 18090
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4172 12170 4200 12786
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11354 3648 11494
rect 4172 11354 4200 12106
rect 4356 11558 4384 12582
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 4172 9926 4200 11290
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3712 7002 3740 7278
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3436 4126 3556 4154
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 848 2304 900 2310
rect 848 2246 900 2252
rect 478 82 534 480
rect 860 82 888 2246
rect 478 54 888 82
rect 1490 82 1546 480
rect 1780 82 1808 3062
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 1490 54 1808 82
rect 2594 82 2650 480
rect 2884 82 2912 2790
rect 3436 134 3464 4126
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2594 54 2912 82
rect 3424 128 3476 134
rect 3424 70 3476 76
rect 3528 82 3556 4014
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 4264 2009 4292 10406
rect 4356 6848 4384 11494
rect 4448 11354 4476 11630
rect 4540 11558 4568 15846
rect 4724 15366 4752 15982
rect 5276 15706 5304 16390
rect 5552 15978 5580 16662
rect 5644 16114 5672 16934
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5552 15638 5580 15914
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4632 12102 4660 12718
rect 4724 12646 4752 15302
rect 5552 15162 5580 15574
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5920 14822 5948 15438
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5078 14512 5134 14521
rect 5078 14447 5134 14456
rect 5092 12850 5120 14447
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5184 12782 5212 13330
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 5184 12306 5212 12718
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5644 12170 5672 12718
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4632 11558 4660 12038
rect 5184 11830 5212 12038
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5184 11694 5212 11766
rect 5644 11694 5672 12106
rect 5736 12102 5764 12242
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5736 11762 5764 12038
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4448 10674 4476 11290
rect 4632 11218 4660 11494
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4632 10606 4660 11154
rect 5184 11150 5212 11630
rect 5736 11354 5764 11698
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 5644 10266 5672 11154
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 5644 10130 5672 10202
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 8090 4568 9862
rect 5644 9722 5672 10066
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9178 5948 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5276 8838 5304 8978
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4908 8566 4936 8774
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4436 6860 4488 6866
rect 4356 6820 4436 6848
rect 4436 6802 4488 6808
rect 4448 6186 4476 6802
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4816 5914 4844 7414
rect 4908 6322 4936 8502
rect 5080 8492 5132 8498
rect 5276 8480 5304 8774
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5080 8434 5132 8440
rect 5184 8452 5396 8480
rect 5092 8294 5120 8434
rect 5184 8362 5212 8452
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7206 5120 8230
rect 5276 7954 5304 8298
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5276 7750 5304 7890
rect 5368 7750 5396 8452
rect 5460 8362 5488 8502
rect 5736 8430 5764 8910
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5632 7880 5684 7886
rect 5736 7868 5764 8366
rect 5684 7840 5764 7868
rect 5632 7822 5684 7828
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5276 7342 5304 7686
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5276 6662 5304 7278
rect 5368 6866 5396 7686
rect 5736 7546 5764 7840
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5460 7206 5488 7278
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4988 6180 5040 6186
rect 4988 6122 5040 6128
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5000 5778 5028 6122
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4988 5772 5040 5778
rect 4988 5714 5040 5720
rect 4908 5370 4936 5714
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 4282 4936 5306
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5092 4078 5120 6054
rect 5184 5370 5212 6598
rect 5368 6390 5396 6802
rect 5460 6730 5488 7142
rect 5736 7002 5764 7482
rect 5828 7274 5856 8434
rect 5920 8362 5948 8774
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5920 7206 5948 7822
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5920 6730 5948 7142
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 4282 5212 4626
rect 5368 4486 5396 6326
rect 5460 5574 5488 6666
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5736 6458 5764 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 4690 5488 5510
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3194 4752 3334
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4908 2582 4936 3946
rect 5184 3602 5212 4218
rect 5368 4010 5396 4422
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3670 5672 3878
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3194 5212 3538
rect 5644 3398 5672 3606
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5736 2990 5764 6394
rect 5920 6254 5948 6666
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 5092 2310 5120 2926
rect 5920 2514 5948 5102
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4250 2000 4306 2009
rect 4250 1935 4306 1944
rect 3606 82 3662 480
rect 3528 54 3662 82
rect 478 0 534 54
rect 1490 0 1546 54
rect 2594 0 2650 54
rect 3606 0 3662 54
rect 4710 82 4766 480
rect 5092 82 5120 2246
rect 4710 54 5120 82
rect 5814 82 5870 480
rect 6012 82 6040 25638
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6656 19922 6684 39646
rect 7104 39636 7156 39642
rect 7104 39578 7156 39584
rect 7930 39636 7986 40000
rect 7930 39584 7932 39636
rect 7984 39584 7986 39636
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6656 19514 6684 19858
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6092 18896 6144 18902
rect 6092 18838 6144 18844
rect 6104 18086 6132 18838
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6104 16250 6132 18022
rect 6196 17610 6224 18702
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18086 6684 18634
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6184 17604 6236 17610
rect 6184 17546 6236 17552
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6196 16794 6224 17274
rect 6656 17270 6684 18022
rect 6748 17678 6776 19654
rect 6932 19242 6960 19654
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6840 18902 6868 19110
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6932 18426 6960 19178
rect 7024 18766 7052 19314
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6840 17882 6868 18226
rect 7024 18154 7052 18702
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 6748 17270 6776 17614
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6736 17264 6788 17270
rect 6736 17206 6788 17212
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6104 5166 6132 16050
rect 6656 15910 6684 16526
rect 6840 16454 6868 17070
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13462 6224 13670
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12306 6224 12582
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6656 12442 6684 15846
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6748 12714 6776 13126
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6644 12300 6696 12306
rect 6748 12288 6776 12650
rect 6696 12260 6776 12288
rect 6644 12242 6696 12248
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6184 11212 6236 11218
rect 6184 11154 6236 11160
rect 6196 10810 6224 11154
rect 6656 10810 6684 12242
rect 6840 11354 6868 16390
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6932 11558 6960 14758
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13870 7052 14214
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7024 13394 7052 13670
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7024 12782 7052 13330
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7012 12164 7064 12170
rect 7012 12106 7064 12112
rect 7024 11626 7052 12106
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 6934 6224 9318
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6656 8634 6684 9590
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6656 8430 6684 8570
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7546 6592 7686
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6656 7478 6684 8366
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6748 5914 6776 11222
rect 7024 11218 7052 11562
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9518 6868 10066
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 7024 9042 7052 9862
rect 7116 9382 7144 39578
rect 7930 39520 7986 39584
rect 9310 39704 9366 40000
rect 9310 39652 9312 39704
rect 9364 39652 9366 39704
rect 9310 39520 9366 39652
rect 9864 39704 9916 39710
rect 9864 39646 9916 39652
rect 9772 39636 9824 39642
rect 9772 39578 9824 39584
rect 8022 37768 8078 37777
rect 8022 37703 8078 37712
rect 8036 34610 8064 37703
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8024 34604 8076 34610
rect 8024 34546 8076 34552
rect 9496 34536 9548 34542
rect 9496 34478 9548 34484
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7484 18086 7512 18838
rect 8024 18692 8076 18698
rect 8024 18634 8076 18640
rect 7840 18352 7892 18358
rect 7840 18294 7892 18300
rect 7748 18148 7800 18154
rect 7668 18108 7748 18136
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7484 17338 7512 18022
rect 7576 17678 7604 18022
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7668 17542 7696 18108
rect 7748 18090 7800 18096
rect 7852 18086 7880 18294
rect 8036 18290 8064 18634
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7472 17332 7524 17338
rect 7472 17274 7524 17280
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7208 16726 7236 16934
rect 7668 16794 7696 17478
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7196 16720 7248 16726
rect 7196 16662 7248 16668
rect 7208 15910 7236 16662
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7208 15366 7236 15846
rect 7484 15366 7512 15982
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7208 14550 7236 15302
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7300 13394 7328 13806
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7484 12646 7512 15302
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7668 13462 7696 13806
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7576 12374 7604 13330
rect 7668 12782 7696 13398
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7668 12442 7696 12718
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7208 11354 7236 12174
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7208 11082 7236 11290
rect 7484 11286 7512 11630
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7208 10606 7236 11018
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7484 10538 7512 11086
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7484 10130 7512 10474
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7668 9654 7696 12378
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7760 10470 7788 10542
rect 7748 10464 7800 10470
rect 7748 10406 7800 10412
rect 7760 10130 7788 10406
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7668 9518 7696 9590
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7024 8294 7052 8978
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7300 8430 7328 8910
rect 7668 8498 7696 8978
rect 7748 8968 7800 8974
rect 7852 8945 7880 18022
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8128 17338 8156 17614
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8772 16454 8800 17002
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8220 16250 8248 16390
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8312 15162 8340 15438
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8864 15026 8892 34342
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 9310 33416 9366 33425
rect 9310 33351 9366 33360
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9324 18426 9352 33351
rect 9508 19334 9536 34478
rect 9508 19306 9628 19334
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9324 17202 9352 18158
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8852 15020 8904 15026
rect 8852 14962 8904 14968
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8680 14618 8708 14826
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 13870 8064 14214
rect 8220 14006 8248 14350
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8024 13864 8076 13870
rect 7944 13812 8024 13814
rect 7944 13806 8076 13812
rect 7944 13786 8064 13806
rect 7944 13394 7972 13786
rect 8680 13734 8708 14418
rect 8864 14346 8892 14962
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 12102 7972 13330
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12782 8064 13126
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8024 12776 8076 12782
rect 8024 12718 8076 12724
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11830 7972 12038
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 10996 7972 11766
rect 8036 11694 8064 12718
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8312 12102 8340 12310
rect 8404 12306 8432 12786
rect 8680 12646 8708 13670
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 9324 12782 9352 13126
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8024 11008 8076 11014
rect 7944 10968 8024 10996
rect 8024 10950 8076 10956
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 7748 8910 7800 8916
rect 7838 8936 7894 8945
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6656 5098 6684 5714
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4826 6132 4966
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6196 4282 6224 4626
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6196 3602 6224 4218
rect 6380 4010 6408 4626
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6656 3602 6684 5034
rect 6748 4690 6776 5850
rect 7024 5370 7052 8230
rect 7300 7818 7328 8366
rect 7668 8090 7696 8434
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 7002 7144 7210
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7116 6458 7144 6938
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7300 5574 7328 7754
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7392 7206 7420 7414
rect 7668 7410 7696 7686
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 7002 7420 7142
rect 7760 7002 7788 8910
rect 7838 8871 7894 8880
rect 7944 8022 7972 10678
rect 8036 10606 8064 10950
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8036 10130 8064 10542
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8036 9518 8064 10066
rect 8128 9654 8156 11086
rect 8312 10470 8340 12038
rect 8404 11558 8432 12242
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8036 9178 8064 9454
rect 8128 9178 8156 9590
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7206 7972 7958
rect 8220 7410 8248 8298
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7760 6322 7788 6938
rect 7944 6934 7972 7142
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7852 6254 7880 6734
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7300 5166 7328 5510
rect 7852 5234 7880 6190
rect 7944 6186 7972 6870
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5574 7972 6122
rect 8128 5778 8156 6394
rect 8312 5914 8340 8230
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7024 3738 7052 4558
rect 7116 4146 7144 4762
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7300 3670 7328 3878
rect 7944 3670 7972 5510
rect 8128 5370 8156 5714
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8404 5098 8432 11494
rect 8588 10742 8616 11630
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8576 10532 8628 10538
rect 8680 10520 8708 11562
rect 8772 11150 8800 11698
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 11354 9168 11630
rect 9324 11558 9352 12718
rect 9416 12442 9444 13670
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9508 11898 9536 12310
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8852 11280 8904 11286
rect 9600 11257 9628 19306
rect 9784 18970 9812 39578
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18086 9720 18770
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17105 9720 17682
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9692 16998 9720 17031
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9784 13814 9812 14486
rect 9692 13786 9812 13814
rect 9692 13734 9720 13786
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9772 12164 9824 12170
rect 9772 12106 9824 12112
rect 8852 11222 8904 11228
rect 9586 11248 9642 11257
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8628 10492 8708 10520
rect 8576 10474 8628 10480
rect 8680 10266 8708 10492
rect 8864 10266 8892 11222
rect 9586 11183 9642 11192
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8680 9722 8708 10202
rect 9232 10198 9260 10542
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8668 9716 8720 9722
rect 9600 9674 9628 11183
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10674 9720 11086
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9784 10198 9812 12106
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 8668 9658 8720 9664
rect 8680 9450 8708 9658
rect 9508 9646 9628 9674
rect 9508 9518 9536 9646
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8680 9110 8708 9386
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8496 8498 8524 8842
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8680 7886 8708 8434
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8680 7274 8708 7822
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8680 6798 8708 7210
rect 9048 7002 9076 7346
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8668 6792 8720 6798
rect 9692 6780 9720 9318
rect 9784 9178 9812 10134
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9784 7546 9812 7958
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9772 6792 9824 6798
rect 9692 6752 9772 6780
rect 8668 6734 8720 6740
rect 9772 6734 9824 6740
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9784 6458 9812 6734
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9876 6338 9904 39646
rect 10782 39636 10838 40000
rect 12254 39658 12310 40000
rect 10782 39584 10784 39636
rect 10836 39584 10838 39636
rect 10782 39520 10838 39584
rect 11992 39630 12310 39658
rect 11518 38176 11574 38185
rect 11518 38111 11574 38120
rect 11336 27872 11388 27878
rect 11336 27814 11388 27820
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 9968 13802 9996 13942
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10060 13802 10088 13874
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 10048 13796 10100 13802
rect 10100 13756 10180 13784
rect 10048 13738 10100 13744
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 10060 12646 10088 13466
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12374 10088 12582
rect 10048 12368 10100 12374
rect 10048 12310 10100 12316
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9968 11694 9996 11834
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10060 11354 10088 12310
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10060 10538 10088 11290
rect 10152 10810 10180 13756
rect 10244 13394 10272 13874
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10336 11694 10364 11766
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 10152 10198 10180 10746
rect 10428 10198 10456 11018
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10152 9722 10180 10134
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9968 8634 9996 8774
rect 10336 8634 10364 8978
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 9968 8294 9996 8570
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 10336 8090 10364 8570
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10428 8022 10456 8298
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10416 7268 10468 7274
rect 10416 7210 10468 7216
rect 10428 6934 10456 7210
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 9784 6310 9904 6338
rect 9968 6322 9996 6870
rect 10428 6390 10456 6870
rect 10520 6390 10548 8842
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 9956 6316 10008 6322
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5846 9720 6054
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 9784 4826 9812 6310
rect 9956 6258 10008 6264
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9876 5914 9904 6122
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9876 5370 9904 5850
rect 10336 5778 10364 6258
rect 10612 6254 10640 16594
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12986 10732 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10796 12442 10824 12718
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11014 10824 12174
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 9586 10824 10950
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10336 5370 10364 5714
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6196 3058 6224 3538
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6196 2650 6224 2994
rect 6656 2922 6684 3538
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6840 3058 6868 3402
rect 7300 3194 7328 3606
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6840 2650 6868 2994
rect 7944 2990 7972 3606
rect 8036 3534 8064 3946
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 8128 2582 8156 4422
rect 8496 4282 8524 4626
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 3936 8444 3942
rect 8496 3924 8524 4218
rect 9968 4010 9996 4626
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 8444 3896 8524 3924
rect 8392 3878 8444 3884
rect 8680 3738 8708 3946
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8772 3670 8800 3946
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8680 3058 8708 3402
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8680 2582 8708 2994
rect 8772 2922 8800 3130
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8864 2650 8892 3878
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 9324 3058 9352 3946
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3194 9812 3538
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8864 2446 8892 2586
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 5814 54 6040 82
rect 6826 128 6882 480
rect 6826 76 6828 128
rect 6880 76 6882 128
rect 4710 0 4766 54
rect 5814 0 5870 54
rect 6826 0 6882 76
rect 7930 82 7986 480
rect 8036 82 8064 2314
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 7930 54 8064 82
rect 8864 82 8892 2246
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8942 82 8998 480
rect 8864 54 8998 82
rect 9968 82 9996 2790
rect 10060 2514 10088 4966
rect 10704 4282 10732 9454
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10704 4154 10732 4218
rect 10612 4146 10732 4154
rect 10600 4140 10732 4146
rect 10652 4126 10732 4140
rect 10600 4082 10652 4088
rect 10612 3194 10640 4082
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10612 2990 10640 3130
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10888 2514 10916 16934
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11256 14074 11284 14350
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11256 13814 11284 14010
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11164 13786 11284 13814
rect 11072 12850 11100 13738
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11164 12170 11192 13786
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 12374 11284 12582
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11256 11354 11284 12310
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11348 10130 11376 27814
rect 11426 19952 11482 19961
rect 11426 19887 11482 19896
rect 11440 17746 11468 19887
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 17338 11468 17682
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11532 13814 11560 38111
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11992 34746 12020 39630
rect 12254 39520 12310 39630
rect 13726 39704 13782 40000
rect 13726 39652 13728 39704
rect 13780 39652 13782 39704
rect 13726 39520 13782 39652
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 15198 39636 15254 40000
rect 15198 39584 15200 39636
rect 15252 39584 15254 39636
rect 11980 34740 12032 34746
rect 11980 34682 12032 34688
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 13634 30832 13690 30841
rect 13634 30767 13690 30776
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 13648 28762 13676 30767
rect 13636 28756 13688 28762
rect 13636 28698 13688 28704
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 13464 27878 13492 28562
rect 13452 27872 13504 27878
rect 13452 27814 13504 27820
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 13634 27432 13690 27441
rect 13634 27367 13690 27376
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 12070 23624 12126 23633
rect 12070 23559 12126 23568
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11440 13786 11560 13814
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9382 11376 10066
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11440 9178 11468 13786
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11716 12986 11744 13398
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11624 11898 11652 12310
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10810 11560 11086
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11808 10742 11836 11222
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11532 8294 11560 8978
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11072 7818 11100 8230
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11520 8016 11572 8022
rect 11520 7958 11572 7964
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11072 7410 11100 7754
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11532 7206 11560 7958
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7546 11836 7822
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11348 6866 11376 7142
rect 11532 7002 11560 7142
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11348 6458 11376 6802
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11992 4154 12020 17478
rect 12084 12782 12112 23559
rect 13648 14618 13676 27367
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12176 13462 12204 14282
rect 13464 13802 13492 14418
rect 13452 13796 13504 13802
rect 13452 13738 13504 13744
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12176 12646 12204 13262
rect 12268 12986 12296 13670
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13634 12744 13690 12753
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11082 12112 12106
rect 12176 11762 12204 12582
rect 13464 12306 13492 12718
rect 13634 12679 13690 12688
rect 13648 12442 13676 12679
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13464 11898 13492 12242
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12636 11626 12664 11834
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12452 11014 12480 11494
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10266 12480 10950
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 5817 12112 9318
rect 12898 8936 12954 8945
rect 12624 8900 12676 8906
rect 12898 8871 12954 8880
rect 12624 8842 12676 8848
rect 12636 8362 12664 8842
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12912 7342 12940 8871
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12070 5808 12126 5817
rect 12070 5743 12126 5752
rect 11992 4126 12112 4154
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10046 82 10102 480
rect 9968 54 10102 82
rect 7930 0 7986 54
rect 8942 0 8998 54
rect 10046 0 10102 54
rect 11150 128 11206 480
rect 12084 134 12112 4126
rect 11150 76 11152 128
rect 11204 76 11206 128
rect 11150 0 11206 76
rect 12072 128 12124 134
rect 12072 70 12124 76
rect 12162 82 12218 480
rect 12268 82 12296 6190
rect 13464 2990 13492 10406
rect 13634 9072 13690 9081
rect 13634 9007 13690 9016
rect 13648 8634 13676 9007
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13740 8430 13768 12786
rect 13832 9178 13860 39578
rect 15198 39520 15254 39584
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 15474 34504 15530 34513
rect 15474 34439 15530 34448
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 15488 33425 15516 34439
rect 15474 33416 15530 33425
rect 15474 33351 15530 33360
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14738 16280 14794 16289
rect 14738 16215 14794 16224
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14752 12850 14780 16215
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12162 54 12296 82
rect 12912 82 12940 2246
rect 13266 82 13322 480
rect 12912 54 13322 82
rect 13924 82 13952 2790
rect 14108 1873 14136 2790
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14094 1864 14150 1873
rect 14094 1799 14150 1808
rect 14278 82 14334 480
rect 13924 54 14334 82
rect 15212 82 15240 2314
rect 15382 82 15438 480
rect 15212 54 15438 82
rect 12162 0 12218 54
rect 13266 0 13322 54
rect 14278 0 14334 54
rect 15382 0 15438 54
<< via2 >>
rect 110 24928 166 24984
rect 110 21664 166 21720
rect 1582 34720 1638 34776
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 1582 17856 1638 17912
rect 4618 27784 4674 27840
rect 5354 31048 5410 31104
rect 1490 17040 1546 17096
rect 110 4936 166 4992
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 5078 14456 5134 14512
rect 4250 1944 4306 2000
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 8022 37712 8078 37768
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9310 33360 9366 33416
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 7838 8880 7894 8936
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 9678 17040 9734 17096
rect 9586 11192 9642 11248
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 11518 38120 11574 38176
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 11426 19896 11482 19952
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 13634 30776 13690 30832
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 13634 27376 13690 27432
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 12070 23568 12126 23624
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 13634 12688 13690 12744
rect 12898 8880 12954 8936
rect 12070 5752 12126 5808
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 13634 9016 13690 9072
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 15474 34448 15530 34504
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 15474 33360 15530 33416
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14738 16224 14794 16280
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 14094 1808 14150 1864
<< metal3 >>
rect 0 38224 480 38344
rect 62 37770 122 38224
rect 11513 38178 11579 38181
rect 15520 38178 16000 38208
rect 11513 38176 16000 38178
rect 11513 38120 11518 38176
rect 11574 38120 16000 38176
rect 11513 38118 16000 38120
rect 11513 38115 11579 38118
rect 15520 38088 16000 38118
rect 8017 37770 8083 37773
rect 62 37768 8083 37770
rect 62 37712 8022 37768
rect 8078 37712 8083 37768
rect 62 37710 8083 37712
rect 8017 37707 8083 37710
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 0 34960 480 35080
rect 62 34778 122 34960
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 1577 34778 1643 34781
rect 62 34776 1643 34778
rect 62 34720 1582 34776
rect 1638 34720 1643 34776
rect 62 34718 1643 34720
rect 1577 34715 1643 34718
rect 15520 34509 16000 34536
rect 15469 34506 16000 34509
rect 15388 34504 16000 34506
rect 15388 34448 15474 34504
rect 15530 34448 16000 34504
rect 15388 34446 16000 34448
rect 15469 34443 16000 34446
rect 15520 34416 16000 34443
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 9305 33418 9371 33421
rect 15469 33418 15535 33421
rect 9305 33416 15535 33418
rect 9305 33360 9310 33416
rect 9366 33360 15474 33416
rect 15530 33360 15535 33416
rect 9305 33358 15535 33360
rect 9305 33355 9371 33358
rect 15469 33355 15535 33358
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 0 31560 480 31680
rect 3610 31584 3930 31585
rect 62 31106 122 31560
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 5349 31106 5415 31109
rect 62 31104 5415 31106
rect 62 31048 5354 31104
rect 5410 31048 5415 31104
rect 62 31046 5415 31048
rect 5349 31043 5415 31046
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 13629 30834 13695 30837
rect 15520 30834 16000 30864
rect 13629 30832 16000 30834
rect 13629 30776 13634 30832
rect 13690 30776 16000 30832
rect 13629 30774 16000 30776
rect 13629 30771 13695 30774
rect 15520 30744 16000 30774
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 0 28296 480 28416
rect 3610 28320 3930 28321
rect 62 27842 122 28296
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 4613 27842 4679 27845
rect 62 27840 4679 27842
rect 62 27784 4618 27840
rect 4674 27784 4679 27840
rect 62 27782 4679 27784
rect 4613 27779 4679 27782
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 13629 27434 13695 27437
rect 13629 27432 15578 27434
rect 13629 27376 13634 27432
rect 13690 27376 15578 27432
rect 13629 27374 15578 27376
rect 13629 27371 13695 27374
rect 15518 27328 15578 27374
rect 15518 27238 16000 27328
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 15520 27208 16000 27238
rect 14277 27167 14597 27168
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 0 24984 480 25016
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 0 24928 110 24984
rect 166 24928 480 24984
rect 0 24896 480 24928
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 12065 23626 12131 23629
rect 15520 23626 16000 23656
rect 12065 23624 16000 23626
rect 12065 23568 12070 23624
rect 12126 23568 16000 23624
rect 12065 23566 16000 23568
rect 12065 23563 12131 23566
rect 15520 23536 16000 23566
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 3610 21792 3930 21793
rect 0 21720 480 21752
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 0 21664 110 21720
rect 166 21664 480 21720
rect 0 21632 480 21664
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 11421 19954 11487 19957
rect 15520 19954 16000 19984
rect 11421 19952 16000 19954
rect 11421 19896 11426 19952
rect 11482 19896 16000 19952
rect 11421 19894 16000 19896
rect 11421 19891 11487 19894
rect 15520 19864 16000 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 0 18232 480 18352
rect 62 17914 122 18232
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 1577 17914 1643 17917
rect 62 17912 1643 17914
rect 62 17856 1582 17912
rect 1638 17856 1643 17912
rect 62 17854 1643 17856
rect 1577 17851 1643 17854
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 1485 17098 1551 17101
rect 9673 17098 9739 17101
rect 1485 17096 9739 17098
rect 1485 17040 1490 17096
rect 1546 17040 9678 17096
rect 9734 17040 9739 17096
rect 1485 17038 9739 17040
rect 1485 17035 1551 17038
rect 9673 17035 9739 17038
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 14733 16282 14799 16285
rect 15520 16282 16000 16312
rect 14733 16280 16000 16282
rect 14733 16224 14738 16280
rect 14794 16224 16000 16280
rect 14733 16222 16000 16224
rect 14733 16219 14799 16222
rect 15520 16192 16000 16222
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 0 14968 480 15088
rect 62 14514 122 14968
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 5073 14514 5139 14517
rect 62 14512 5139 14514
rect 62 14456 5078 14512
rect 5134 14456 5139 14512
rect 62 14454 5139 14456
rect 5073 14451 5139 14454
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 13629 12746 13695 12749
rect 15520 12746 16000 12776
rect 13629 12744 16000 12746
rect 13629 12688 13634 12744
rect 13690 12688 16000 12744
rect 13629 12686 16000 12688
rect 13629 12683 13695 12686
rect 15520 12656 16000 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 0 11660 480 11688
rect 0 11596 60 11660
rect 124 11596 480 11660
rect 0 11568 480 11596
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 54 11188 60 11252
rect 124 11250 130 11252
rect 9581 11250 9647 11253
rect 124 11248 9647 11250
rect 124 11192 9586 11248
rect 9642 11192 9647 11248
rect 124 11190 9647 11192
rect 124 11188 130 11190
rect 9581 11187 9647 11190
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 13629 9074 13695 9077
rect 15520 9074 16000 9104
rect 13629 9072 16000 9074
rect 13629 9016 13634 9072
rect 13690 9016 16000 9072
rect 13629 9014 16000 9016
rect 13629 9011 13695 9014
rect 15520 8984 16000 9014
rect 7833 8938 7899 8941
rect 12893 8938 12959 8941
rect 62 8936 12959 8938
rect 62 8880 7838 8936
rect 7894 8880 12898 8936
rect 12954 8880 12959 8936
rect 62 8878 12959 8880
rect 62 8424 122 8878
rect 7833 8875 7899 8878
rect 12893 8875 12959 8878
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 0 8304 480 8424
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 12065 5810 12131 5813
rect 12065 5808 15578 5810
rect 12065 5752 12070 5808
rect 12126 5752 15578 5808
rect 12065 5750 15578 5752
rect 12065 5747 12131 5750
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 15518 5432 15578 5750
rect 15518 5342 16000 5432
rect 15520 5312 16000 5342
rect 0 4992 480 5024
rect 0 4936 110 4992
rect 166 4936 480 4992
rect 0 4904 480 4936
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 4245 2002 4311 2005
rect 62 2000 4311 2002
rect 62 1944 4250 2000
rect 4306 1944 4311 2000
rect 62 1942 4311 1944
rect 62 1760 122 1942
rect 4245 1939 4311 1942
rect 14089 1866 14155 1869
rect 15520 1866 16000 1896
rect 14089 1864 16000 1866
rect 14089 1808 14094 1864
rect 14150 1808 16000 1864
rect 14089 1806 16000 1808
rect 14089 1803 14155 1806
rect 15520 1776 16000 1806
rect 0 1640 480 1760
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 60 11596 124 11660
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 60 11188 124 11252
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 59 11660 125 11661
rect 59 11596 60 11660
rect 124 11596 125 11660
rect 59 11595 125 11596
rect 62 11253 122 11595
rect 59 11252 125 11253
rect 59 11188 60 11252
rect 124 11188 125 11252
rect 59 11187 125 11188
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_8  _33_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4140 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__33__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_1_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_42
timestamp 1586364061
transform 1 0 4968 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__C
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_46
timestamp 1586364061
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__B
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _82_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_8  _61_
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_58 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__82__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_81
timestamp 1586364061
transform 1 0 8556 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_73
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_77
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_90
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_102
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_114
timestamp 1586364061
transform 1 0 11592 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_122
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_138
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__91__A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__93__A
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _93_
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _91_
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_nor4_4  _64_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__63__C
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_8  _69_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 774 592
use scs8hd_conb_1  _75_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_137
timestamp 1586364061
transform 1 0 13708 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_or2_4  _62_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__D
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__B
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_121
timestamp 1586364061
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_143
timestamp 1586364061
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_nor4_4  _63_
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__62__B
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_8  _70_
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_82
timestamp 1586364061
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_96
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_120
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_144
timestamp 1586364061
transform 1 0 14352 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__32__A
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_43 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _60_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7176 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__31__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_79
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_40
timestamp 1586364061
transform 1 0 4784 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _32_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_49
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__34__A
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_8  _54_
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _31_
timestamp 1586364061
transform 1 0 5888 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__34__B
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__C
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_65
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__60__B
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__34__D
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _66_
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_73
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_103
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _68_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__B
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use scs8hd_or4_4  _34_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 866 592
use scs8hd_buf_1  _37_
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__46__C
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_8  _67_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _56_
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _45_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__D
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_36
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_40
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__B
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_72
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_76
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _47_
timestamp 1586364061
transform 1 0 4324 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use scs8hd_or4_4  _46_
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__55__B
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_38
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_42
timestamp 1586364061
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__D
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__B
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__B
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_59
timestamp 1586364061
transform 1 0 6532 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 774 592
use scs8hd_conb_1  _74_
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_130
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_142
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__55__C
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 130 592
use scs8hd_or4_4  _55_
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _59_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__58__B
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _72_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 406 592
use scs8hd_decap_6  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_buf_2  _84_
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__84__A
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use scs8hd_or4_4  _58_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__55__D
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__C
timestamp 1586364061
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_42
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _57_
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__42__D
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__42__B
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_75
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_79
timestamp 1586364061
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_8  _65_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_110
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_116
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_127
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_139
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__50__D
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__B
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_47
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_buf_1  _35_
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_51
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _41_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1602 592
use scs8hd_nor4_4  _42_
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__41__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__35__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__C
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__C
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_57
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__B
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__D
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__41__B
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_87
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_113
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_137
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__29__A
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 130 592
use scs8hd_inv_8  _39_
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__C
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_49
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _44_
timestamp 1586364061
transform 1 0 6900 0 1 10336
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__B
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__C
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_80
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_84
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_99
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_103
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__49__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_1  _29_
timestamp 1586364061
transform 1 0 4600 0 -1 11424
box -38 -48 314 592
use scs8hd_nor4_4  _50_
timestamp 1586364061
transform 1 0 5612 0 -1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_41
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_46
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__52__C
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_66
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__D
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_74
timestamp 1586364061
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_89
timestamp 1586364061
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__51__C
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__B
timestamp 1586364061
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__D
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_23
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_32
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _51_
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _52_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _43_
timestamp 1586364061
transform 1 0 9108 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_79
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_83
timestamp 1586364061
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__43__D
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__43__B
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_116
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_144
timestamp 1586364061
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_buf_1  _40_
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__30__A
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__D
timestamp 1586364061
transform 1 0 4968 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_38
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_51
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _49_
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 1602 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__43__C
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__D
timestamp 1586364061
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__C
timestamp 1586364061
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_72
timestamp 1586364061
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_76
timestamp 1586364061
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_104
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_133
timestamp 1586364061
transform 1 0 13340 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__53__C
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__D
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_8  _30_
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use scs8hd_nor4_4  _53_
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__53__B
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_38
timestamp 1586364061
transform 1 0 4600 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _38_
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 1602 592
use scs8hd_nor4_4  _48_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__38__B
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__C
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_57
timestamp 1586364061
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_78
timestamp 1586364061
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__D
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_86
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_82
timestamp 1586364061
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__B
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_102
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_109
timestamp 1586364061
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_142
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_133
timestamp 1586364061
transform 1 0 13340 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 406 592
use scs8hd_nor4_4  _36_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__C
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_83
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_87
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_120
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__89__A
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_131
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__36__B
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__36__D
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_91
timestamp 1586364061
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_114
timestamp 1586364061
transform 1 0 11592 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _89_
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_126
timestamp 1586364061
transform 1 0 12696 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_138
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_49
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_89
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_101
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_143
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_58
timestamp 1586364061
transform 1 0 6440 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_67
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 590 592
use scs8hd_conb_1  _71_
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_77
timestamp 1586364061
transform 1 0 8188 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_81
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_89
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_38
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_78
timestamp 1586364061
transform 1 0 8280 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_102
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_19
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_30
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_40
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_36
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_42
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5336 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7084 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_76
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_27_143
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_19
timestamp 1586364061
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_55
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _73_
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_91
timestamp 1586364061
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_96
timestamp 1586364061
transform 1 0 9936 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_116
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_28_140
timestamp 1586364061
transform 1 0 13984 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 314 592
use scs8hd_decap_6  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_79
timestamp 1586364061
transform 1 0 8372 0 1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__92__A
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_107
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_119
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_43
timestamp 1586364061
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_47
timestamp 1586364061
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use scs8hd_buf_2  _92_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_97
timestamp 1586364061
transform 1 0 10028 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_109
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_121
timestamp 1586364061
transform 1 0 12236 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_133
timestamp 1586364061
transform 1 0 13340 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_buf_2  _83_
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__83__A
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_47
timestamp 1586364061
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_55
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_58
timestamp 1586364061
transform 1 0 6440 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_119
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_143
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_59
timestamp 1586364061
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_76
timestamp 1586364061
transform 1 0 8096 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_19
timestamp 1586364061
transform 1 0 2852 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_55
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_7
timestamp 1586364061
transform 1 0 1748 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_19
timestamp 1586364061
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_105
timestamp 1586364061
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_117
timestamp 1586364061
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_129
timestamp 1586364061
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_1  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_43_35
timestamp 1586364061
transform 1 0 4324 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__88__A
timestamp 1586364061
transform 1 0 4416 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_38
timestamp 1586364061
transform 1 0 4600 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_50
timestamp 1586364061
transform 1 0 5704 0 1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_43_58
timestamp 1586364061
transform 1 0 6440 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_98
timestamp 1586364061
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_4  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 406 592
use scs8hd_buf_2  _88_
timestamp 1586364061
transform 1 0 4416 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_40
timestamp 1586364061
transform 1 0 4784 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_52
timestamp 1586364061
transform 1 0 5888 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_64
timestamp 1586364061
transform 1 0 6992 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_76
timestamp 1586364061
transform 1 0 8096 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_88
timestamp 1586364061
transform 1 0 9200 0 -1 26656
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_117
timestamp 1586364061
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_129
timestamp 1586364061
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_44_141
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_105
timestamp 1586364061
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_110
timestamp 1586364061
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__85__A
timestamp 1586364061
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_46_141
timestamp 1586364061
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_3  FILLER_47_131
timestamp 1586364061
transform 1 0 13156 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_47_136
timestamp 1586364061
transform 1 0 13616 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_144
timestamp 1586364061
transform 1 0 14352 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_105
timestamp 1586364061
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use scs8hd_buf_2  _85_
timestamp 1586364061
transform 1 0 13432 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_4  FILLER_48_129
timestamp 1586364061
transform 1 0 12972 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_133
timestamp 1586364061
transform 1 0 13340 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_138
timestamp 1586364061
transform 1 0 13800 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__87__A
timestamp 1586364061
transform 1 0 5152 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_43
timestamp 1586364061
transform 1 0 5060 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_46
timestamp 1586364061
transform 1 0 5336 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_decap_3  FILLER_49_58
timestamp 1586364061
transform 1 0 6440 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_98
timestamp 1586364061
transform 1 0 10120 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_110
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_buf_2  _87_
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_48
timestamp 1586364061
transform 1 0 5520 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_60
timestamp 1586364061
transform 1 0 6624 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_72
timestamp 1586364061
transform 1 0 7728 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_84
timestamp 1586364061
transform 1 0 8832 0 -1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_129
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_141
timestamp 1586364061
transform 1 0 14076 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_98
timestamp 1586364061
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_110
timestamp 1586364061
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_129
timestamp 1586364061
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_141
timestamp 1586364061
transform 1 0 14076 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_56_145
timestamp 1586364061
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_110
timestamp 1586364061
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_143
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_141
timestamp 1586364061
transform 1 0 14076 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_buf_2  _86_
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__86__A
timestamp 1586364061
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_7
timestamp 1586364061
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_11
timestamp 1586364061
transform 1 0 2116 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_23
timestamp 1586364061
transform 1 0 3220 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_35
timestamp 1586364061
transform 1 0 4324 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_47
timestamp 1586364061
transform 1 0 5428 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_79
timestamp 1586364061
transform 1 0 8372 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_83
timestamp 1586364061
transform 1 0 8740 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _90_
timestamp 1586364061
transform 1 0 10672 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_95
timestamp 1586364061
transform 1 0 9844 0 1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_59_103
timestamp 1586364061
transform 1 0 10580 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__90__A
timestamp 1586364061
transform 1 0 11224 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_108
timestamp 1586364061
transform 1 0 11040 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_59_112
timestamp 1586364061
transform 1 0 11408 0 1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_120
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_143
timestamp 1586364061
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 2594 0 2650 480 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 1640 480 1760 6 address[1]
port 1 nsew default input
rlabel metal2 s 662 39520 718 40000 6 address[2]
port 2 nsew default input
rlabel metal2 s 3606 0 3662 480 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 4904 480 5024 6 address[4]
port 4 nsew default input
rlabel metal2 s 4710 0 4766 480 6 address[5]
port 5 nsew default input
rlabel metal3 s 15520 1776 16000 1896 6 chany_bottom_in[0]
port 6 nsew default input
rlabel metal3 s 0 8304 480 8424 6 chany_bottom_in[1]
port 7 nsew default input
rlabel metal2 s 2042 39520 2098 40000 6 chany_bottom_in[2]
port 8 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chany_bottom_in[3]
port 9 nsew default input
rlabel metal3 s 0 14968 480 15088 6 chany_bottom_in[4]
port 10 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[5]
port 11 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_in[6]
port 12 nsew default input
rlabel metal2 s 3514 39520 3570 40000 6 chany_bottom_in[7]
port 13 nsew default input
rlabel metal3 s 15520 5312 16000 5432 6 chany_bottom_in[8]
port 14 nsew default input
rlabel metal3 s 15520 8984 16000 9104 6 chany_bottom_out[0]
port 15 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_bottom_out[1]
port 16 nsew default tristate
rlabel metal2 s 7930 0 7986 480 6 chany_bottom_out[2]
port 17 nsew default tristate
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_out[3]
port 18 nsew default tristate
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_out[4]
port 19 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_out[5]
port 20 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chany_bottom_out[6]
port 21 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chany_bottom_out[7]
port 22 nsew default tristate
rlabel metal3 s 15520 12656 16000 12776 6 chany_bottom_out[8]
port 23 nsew default tristate
rlabel metal3 s 15520 16192 16000 16312 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 6458 39520 6514 40000 6 chany_top_in[2]
port 26 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 7930 39520 7986 40000 6 chany_top_in[4]
port 28 nsew default input
rlabel metal3 s 15520 19864 16000 19984 6 chany_top_in[5]
port 29 nsew default input
rlabel metal2 s 9310 39520 9366 40000 6 chany_top_in[6]
port 30 nsew default input
rlabel metal3 s 0 24896 480 25016 6 chany_top_in[7]
port 31 nsew default input
rlabel metal3 s 15520 23536 16000 23656 6 chany_top_in[8]
port 32 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal2 s 10782 39520 10838 40000 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 12254 39520 12310 40000 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal3 s 15520 27208 16000 27328 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal3 s 0 28296 480 28416 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal3 s 0 31560 480 31680 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal3 s 0 34960 480 35080 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal3 s 15520 30744 16000 30864 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 data_in
port 42 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 43 nsew default input
rlabel metal3 s 15520 34416 16000 34536 6 left_grid_pin_1_
port 44 nsew default tristate
rlabel metal3 s 15520 38088 16000 38208 6 left_grid_pin_5_
port 45 nsew default tristate
rlabel metal2 s 13726 39520 13782 40000 6 left_grid_pin_9_
port 46 nsew default tristate
rlabel metal3 s 0 38224 480 38344 6 right_grid_pin_3_
port 47 nsew default tristate
rlabel metal2 s 15198 39520 15254 40000 6 right_grid_pin_7_
port 48 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 49 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 50 nsew default input
<< end >>
