magic
tech sky130A
magscale 1 2
timestamp 1609024634
<< locali >>
rect 8493 17663 8527 17833
rect 9505 14331 9539 14569
rect 12265 12631 12299 12733
rect 12173 3451 12207 3621
<< viali >>
rect 1961 20553 1995 20587
rect 6561 20553 6595 20587
rect 8217 20553 8251 20587
rect 2329 20485 2363 20519
rect 6101 20417 6135 20451
rect 6285 20417 6319 20451
rect 1777 20349 1811 20383
rect 2145 20349 2179 20383
rect 4997 20349 5031 20383
rect 5457 20281 5491 20315
rect 7389 20281 7423 20315
rect 5641 20213 5675 20247
rect 6009 20213 6043 20247
rect 7113 20213 7147 20247
rect 9597 20213 9631 20247
rect 1593 20009 1627 20043
rect 1961 20009 1995 20043
rect 4537 20009 4571 20043
rect 6837 20009 6871 20043
rect 6929 20009 6963 20043
rect 7297 20009 7331 20043
rect 7757 20009 7791 20043
rect 10057 20009 10091 20043
rect 10149 20009 10183 20043
rect 10609 20009 10643 20043
rect 12817 20009 12851 20043
rect 13277 20009 13311 20043
rect 13737 20009 13771 20043
rect 14749 20009 14783 20043
rect 16497 20009 16531 20043
rect 1409 19873 1443 19907
rect 1777 19873 1811 19907
rect 2237 19873 2271 19907
rect 3525 19873 3559 19907
rect 4445 19873 4479 19907
rect 5264 19873 5298 19907
rect 7665 19873 7699 19907
rect 8392 19873 8426 19907
rect 10977 19873 11011 19907
rect 11244 19873 11278 19907
rect 12633 19873 12667 19907
rect 13093 19873 13127 19907
rect 13553 19873 13587 19907
rect 13921 19873 13955 19907
rect 14565 19873 14599 19907
rect 16313 19873 16347 19907
rect 16681 19873 16715 19907
rect 17049 19873 17083 19907
rect 2421 19805 2455 19839
rect 3617 19805 3651 19839
rect 4721 19805 4755 19839
rect 4997 19805 5031 19839
rect 7113 19805 7147 19839
rect 7941 19805 7975 19839
rect 8125 19805 8159 19839
rect 10333 19805 10367 19839
rect 4077 19737 4111 19771
rect 6469 19737 6503 19771
rect 16865 19737 16899 19771
rect 6377 19669 6411 19703
rect 9505 19669 9539 19703
rect 9689 19669 9723 19703
rect 12357 19669 12391 19703
rect 12449 19669 12483 19703
rect 14381 19669 14415 19703
rect 14933 19669 14967 19703
rect 16129 19669 16163 19703
rect 18705 19669 18739 19703
rect 19073 19669 19107 19703
rect 1685 19465 1719 19499
rect 2421 19465 2455 19499
rect 4629 19465 4663 19499
rect 6101 19465 6135 19499
rect 12173 19465 12207 19499
rect 14657 19465 14691 19499
rect 14289 19397 14323 19431
rect 2053 19329 2087 19363
rect 2881 19329 2915 19363
rect 3065 19329 3099 19363
rect 7021 19329 7055 19363
rect 8677 19329 8711 19363
rect 12633 19329 12667 19363
rect 1501 19261 1535 19295
rect 1869 19261 1903 19295
rect 2789 19261 2823 19295
rect 3249 19261 3283 19295
rect 4721 19261 4755 19295
rect 4977 19261 5011 19295
rect 6193 19261 6227 19295
rect 7288 19261 7322 19295
rect 8493 19261 8527 19295
rect 9137 19261 9171 19295
rect 9404 19261 9438 19295
rect 10793 19261 10827 19295
rect 12449 19261 12483 19295
rect 13001 19261 13035 19295
rect 13277 19261 13311 19295
rect 13553 19261 13587 19295
rect 13921 19261 13955 19295
rect 14473 19261 14507 19295
rect 14841 19261 14875 19295
rect 15209 19261 15243 19295
rect 15669 19261 15703 19295
rect 16037 19261 16071 19295
rect 16589 19261 16623 19295
rect 17509 19261 17543 19295
rect 18061 19261 18095 19295
rect 18429 19261 18463 19295
rect 18797 19261 18831 19295
rect 19165 19261 19199 19295
rect 19533 19261 19567 19295
rect 3516 19193 3550 19227
rect 6469 19193 6503 19227
rect 11060 19193 11094 19227
rect 17233 19193 17267 19227
rect 8401 19125 8435 19159
rect 10517 19125 10551 19159
rect 13737 19125 13771 19159
rect 14105 19125 14139 19159
rect 15025 19125 15059 19159
rect 15393 19125 15427 19159
rect 15853 19125 15887 19159
rect 16221 19125 16255 19159
rect 17693 19125 17727 19159
rect 18245 19125 18279 19159
rect 18613 19125 18647 19159
rect 18981 19125 19015 19159
rect 19349 19125 19383 19159
rect 19717 19125 19751 19159
rect 1593 18921 1627 18955
rect 1961 18921 1995 18955
rect 8309 18921 8343 18955
rect 8769 18921 8803 18955
rect 9229 18921 9263 18955
rect 12265 18921 12299 18955
rect 18521 18921 18555 18955
rect 2513 18853 2547 18887
rect 5264 18853 5298 18887
rect 7196 18853 7230 18887
rect 12173 18853 12207 18887
rect 12633 18853 12667 18887
rect 14381 18853 14415 18887
rect 14933 18853 14967 18887
rect 16957 18853 16991 18887
rect 18981 18853 19015 18887
rect 1409 18785 1443 18819
rect 1777 18785 1811 18819
rect 2247 18785 2281 18819
rect 3617 18785 3651 18819
rect 4445 18785 4479 18819
rect 4997 18785 5031 18819
rect 6929 18785 6963 18819
rect 9137 18785 9171 18819
rect 9689 18785 9723 18819
rect 10241 18785 10275 18819
rect 11253 18785 11287 18819
rect 14105 18785 14139 18819
rect 14657 18785 14691 18819
rect 16681 18785 16715 18819
rect 18705 18785 18739 18819
rect 4537 18717 4571 18751
rect 4629 18717 4663 18751
rect 9321 18717 9355 18751
rect 10425 18717 10459 18751
rect 11345 18717 11379 18751
rect 11437 18717 11471 18751
rect 12357 18717 12391 18751
rect 17417 18717 17451 18751
rect 17601 18717 17635 18751
rect 4077 18649 4111 18683
rect 6377 18581 6411 18615
rect 10885 18581 10919 18615
rect 11805 18581 11839 18615
rect 12909 18581 12943 18615
rect 15393 18581 15427 18615
rect 15577 18581 15611 18615
rect 17969 18581 18003 18615
rect 2329 18377 2363 18411
rect 3985 18377 4019 18411
rect 4261 18377 4295 18411
rect 10885 18377 10919 18411
rect 13829 18377 13863 18411
rect 1961 18309 1995 18343
rect 5089 18309 5123 18343
rect 2605 18241 2639 18275
rect 4905 18241 4939 18275
rect 5549 18241 5583 18275
rect 5733 18241 5767 18275
rect 9505 18241 9539 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 1777 18173 1811 18207
rect 2145 18173 2179 18207
rect 2872 18173 2906 18207
rect 10701 18173 10735 18207
rect 11253 18173 11287 18207
rect 11345 18173 11379 18207
rect 12456 18173 12490 18207
rect 4721 18105 4755 18139
rect 5457 18105 5491 18139
rect 5917 18105 5951 18139
rect 12694 18105 12728 18139
rect 1409 18037 1443 18071
rect 4169 18037 4203 18071
rect 4629 18037 4663 18071
rect 8861 18037 8895 18071
rect 9229 18037 9263 18071
rect 9321 18037 9355 18071
rect 4537 17833 4571 17867
rect 4905 17833 4939 17867
rect 5181 17833 5215 17867
rect 8493 17833 8527 17867
rect 8585 17833 8619 17867
rect 8769 17833 8803 17867
rect 11069 17833 11103 17867
rect 13737 17833 13771 17867
rect 2237 17765 2271 17799
rect 2789 17765 2823 17799
rect 1593 17697 1627 17731
rect 1961 17697 1995 17731
rect 2513 17697 2547 17731
rect 4445 17697 4479 17731
rect 6929 17697 6963 17731
rect 11406 17765 11440 17799
rect 9137 17697 9171 17731
rect 9956 17697 9990 17731
rect 11161 17697 11195 17731
rect 13553 17697 13587 17731
rect 4721 17629 4755 17663
rect 6377 17629 6411 17663
rect 7021 17629 7055 17663
rect 7205 17629 7239 17663
rect 8493 17629 8527 17663
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 9689 17629 9723 17663
rect 1777 17561 1811 17595
rect 4077 17561 4111 17595
rect 3801 17493 3835 17527
rect 6561 17493 6595 17527
rect 12541 17493 12575 17527
rect 1777 17289 1811 17323
rect 4813 17289 4847 17323
rect 6285 17289 6319 17323
rect 9689 17289 9723 17323
rect 11161 17289 11195 17323
rect 2145 17153 2179 17187
rect 3065 17153 3099 17187
rect 3249 17153 3283 17187
rect 3433 17153 3467 17187
rect 6469 17153 6503 17187
rect 6837 17153 6871 17187
rect 8309 17153 8343 17187
rect 12081 17153 12115 17187
rect 13369 17153 13403 17187
rect 1593 17085 1627 17119
rect 1961 17085 1995 17119
rect 3700 17085 3734 17119
rect 4905 17085 4939 17119
rect 5161 17085 5195 17119
rect 7104 17085 7138 17119
rect 9781 17085 9815 17119
rect 10037 17085 10071 17119
rect 11897 17085 11931 17119
rect 12541 17085 12575 17119
rect 13093 17085 13127 17119
rect 8554 17017 8588 17051
rect 2605 16949 2639 16983
rect 2973 16949 3007 16983
rect 8217 16949 8251 16983
rect 11253 16949 11287 16983
rect 11529 16949 11563 16983
rect 11989 16949 12023 16983
rect 12725 16949 12759 16983
rect 1593 16745 1627 16779
rect 1961 16745 1995 16779
rect 3617 16745 3651 16779
rect 6561 16745 6595 16779
rect 7113 16745 7147 16779
rect 7205 16745 7239 16779
rect 7665 16745 7699 16779
rect 9137 16745 9171 16779
rect 9689 16745 9723 16779
rect 10057 16745 10091 16779
rect 10977 16745 11011 16779
rect 11345 16745 11379 16779
rect 12265 16745 12299 16779
rect 2421 16677 2455 16711
rect 3525 16677 3559 16711
rect 4537 16677 4571 16711
rect 12173 16677 12207 16711
rect 1409 16609 1443 16643
rect 1777 16609 1811 16643
rect 2145 16609 2179 16643
rect 4445 16609 4479 16643
rect 5437 16609 5471 16643
rect 8033 16609 8067 16643
rect 8125 16609 8159 16643
rect 8769 16609 8803 16643
rect 10885 16609 10919 16643
rect 4721 16541 4755 16575
rect 5181 16541 5215 16575
rect 7389 16541 7423 16575
rect 8217 16541 8251 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 10609 16541 10643 16575
rect 11437 16541 11471 16575
rect 11621 16541 11655 16575
rect 12357 16541 12391 16575
rect 6745 16473 6779 16507
rect 11805 16473 11839 16507
rect 4077 16405 4111 16439
rect 8585 16405 8619 16439
rect 10701 16405 10735 16439
rect 1961 16201 1995 16235
rect 5181 16201 5215 16235
rect 7941 16201 7975 16235
rect 6193 16133 6227 16167
rect 2329 16065 2363 16099
rect 3801 16065 3835 16099
rect 8401 16065 8435 16099
rect 8493 16065 8527 16099
rect 8769 16065 8803 16099
rect 10885 16065 10919 16099
rect 11713 16065 11747 16099
rect 1777 15997 1811 16031
rect 2145 15997 2179 16031
rect 6377 15997 6411 16031
rect 10701 15997 10735 16031
rect 13461 15997 13495 16031
rect 4068 15929 4102 15963
rect 11529 15929 11563 15963
rect 13728 15929 13762 15963
rect 8309 15861 8343 15895
rect 8953 15861 8987 15895
rect 10241 15861 10275 15895
rect 10609 15861 10643 15895
rect 11069 15861 11103 15895
rect 11437 15861 11471 15895
rect 14841 15861 14875 15895
rect 2789 15657 2823 15691
rect 4077 15657 4111 15691
rect 4537 15657 4571 15691
rect 8677 15657 8711 15691
rect 9413 15657 9447 15691
rect 9689 15657 9723 15691
rect 10793 15657 10827 15691
rect 12633 15657 12667 15691
rect 14105 15657 14139 15691
rect 9321 15589 9355 15623
rect 10057 15589 10091 15623
rect 10885 15589 10919 15623
rect 11498 15589 11532 15623
rect 14657 15589 14691 15623
rect 2053 15521 2087 15555
rect 2605 15521 2639 15555
rect 3893 15521 3927 15555
rect 4445 15521 4479 15555
rect 4905 15521 4939 15555
rect 5825 15521 5859 15555
rect 6092 15521 6126 15555
rect 7553 15521 7587 15555
rect 12725 15521 12759 15555
rect 12992 15521 13026 15555
rect 14565 15521 14599 15555
rect 2237 15453 2271 15487
rect 4629 15453 4663 15487
rect 7297 15453 7331 15487
rect 10149 15453 10183 15487
rect 10333 15453 10367 15487
rect 11253 15453 11287 15487
rect 14749 15453 14783 15487
rect 14197 15385 14231 15419
rect 7205 15317 7239 15351
rect 11069 15317 11103 15351
rect 5917 15113 5951 15147
rect 8677 15113 8711 15147
rect 8953 15113 8987 15147
rect 11345 15113 11379 15147
rect 13369 15113 13403 15147
rect 7941 15045 7975 15079
rect 9045 15045 9079 15079
rect 14197 15045 14231 15079
rect 2881 14977 2915 15011
rect 3801 14977 3835 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 9505 14977 9539 15011
rect 9689 14977 9723 15011
rect 11989 14977 12023 15011
rect 13093 14977 13127 15011
rect 13921 14977 13955 15011
rect 2053 14909 2087 14943
rect 2329 14909 2363 14943
rect 2605 14909 2639 14943
rect 8125 14909 8159 14943
rect 9413 14909 9447 14943
rect 9873 14909 9907 14943
rect 10140 14909 10174 14943
rect 12909 14909 12943 14943
rect 13829 14909 13863 14943
rect 14381 14909 14415 14943
rect 14648 14909 14682 14943
rect 6285 14841 6319 14875
rect 7205 14841 7239 14875
rect 7665 14841 7699 14875
rect 11713 14841 11747 14875
rect 13737 14841 13771 14875
rect 3157 14773 3191 14807
rect 3525 14773 3559 14807
rect 3617 14773 3651 14807
rect 6377 14773 6411 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 11253 14773 11287 14807
rect 11805 14773 11839 14807
rect 12541 14773 12575 14807
rect 13001 14773 13035 14807
rect 15761 14773 15795 14807
rect 1961 14569 1995 14603
rect 2329 14569 2363 14603
rect 3893 14569 3927 14603
rect 5457 14569 5491 14603
rect 7205 14569 7239 14603
rect 7665 14569 7699 14603
rect 8217 14569 8251 14603
rect 8677 14569 8711 14603
rect 9045 14569 9079 14603
rect 9413 14569 9447 14603
rect 9505 14569 9539 14603
rect 11529 14569 11563 14603
rect 12633 14569 12667 14603
rect 13093 14569 13127 14603
rect 14657 14569 14691 14603
rect 15393 14569 15427 14603
rect 4322 14501 4356 14535
rect 5816 14501 5850 14535
rect 1777 14433 1811 14467
rect 2145 14433 2179 14467
rect 2780 14433 2814 14467
rect 7573 14433 7607 14467
rect 8033 14433 8067 14467
rect 8585 14433 8619 14467
rect 9229 14433 9263 14467
rect 2513 14365 2547 14399
rect 4077 14365 4111 14399
rect 5549 14365 5583 14399
rect 7757 14365 7791 14399
rect 8769 14365 8803 14399
rect 11345 14501 11379 14535
rect 12725 14501 12759 14535
rect 13461 14501 13495 14535
rect 13921 14501 13955 14535
rect 14565 14501 14599 14535
rect 15025 14501 15059 14535
rect 9689 14433 9723 14467
rect 9965 14433 9999 14467
rect 10149 14433 10183 14467
rect 10425 14433 10459 14467
rect 10885 14433 10919 14467
rect 10977 14365 11011 14399
rect 11161 14365 11195 14399
rect 12817 14365 12851 14399
rect 13553 14365 13587 14399
rect 13737 14365 13771 14399
rect 14749 14365 14783 14399
rect 6929 14297 6963 14331
rect 9505 14297 9539 14331
rect 12265 14297 12299 14331
rect 7021 14229 7055 14263
rect 10241 14229 10275 14263
rect 10517 14229 10551 14263
rect 12081 14229 12115 14263
rect 14197 14229 14231 14263
rect 1869 14025 1903 14059
rect 2789 14025 2823 14059
rect 3341 14025 3375 14059
rect 4721 14025 4755 14059
rect 9321 14025 9355 14059
rect 10333 14025 10367 14059
rect 13553 14025 13587 14059
rect 14381 14025 14415 14059
rect 15577 14025 15611 14059
rect 14657 13957 14691 13991
rect 3893 13889 3927 13923
rect 5273 13889 5307 13923
rect 7665 13889 7699 13923
rect 10057 13889 10091 13923
rect 10793 13889 10827 13923
rect 10977 13889 11011 13923
rect 13369 13889 13403 13923
rect 14013 13889 14047 13923
rect 14197 13889 14231 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 1685 13821 1719 13855
rect 2053 13821 2087 13855
rect 2329 13821 2363 13855
rect 2605 13821 2639 13855
rect 5181 13821 5215 13855
rect 5733 13821 5767 13855
rect 5917 13821 5951 13855
rect 7573 13821 7607 13855
rect 7941 13821 7975 13855
rect 9873 13821 9907 13855
rect 12081 13821 12115 13855
rect 13093 13821 13127 13855
rect 15025 13821 15059 13855
rect 3709 13753 3743 13787
rect 4169 13753 4203 13787
rect 5089 13753 5123 13787
rect 7481 13753 7515 13787
rect 8208 13753 8242 13787
rect 9781 13753 9815 13787
rect 10701 13753 10735 13787
rect 12173 13753 12207 13787
rect 12633 13753 12667 13787
rect 13921 13753 13955 13787
rect 3249 13685 3283 13719
rect 3801 13685 3835 13719
rect 5549 13685 5583 13719
rect 7113 13685 7147 13719
rect 9413 13685 9447 13719
rect 11161 13685 11195 13719
rect 11897 13685 11931 13719
rect 12725 13685 12759 13719
rect 13185 13685 13219 13719
rect 1777 13481 1811 13515
rect 2421 13481 2455 13515
rect 2881 13481 2915 13515
rect 6009 13481 6043 13515
rect 6377 13481 6411 13515
rect 7757 13481 7791 13515
rect 8309 13481 8343 13515
rect 8677 13481 8711 13515
rect 9137 13481 9171 13515
rect 9505 13481 9539 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 10149 13481 10183 13515
rect 13001 13481 13035 13515
rect 14289 13481 14323 13515
rect 15761 13481 15795 13515
rect 17785 13481 17819 13515
rect 4804 13413 4838 13447
rect 7665 13413 7699 13447
rect 1593 13345 1627 13379
rect 2329 13345 2363 13379
rect 3249 13345 3283 13379
rect 4537 13345 4571 13379
rect 6929 13345 6963 13379
rect 11796 13345 11830 13379
rect 13369 13345 13403 13379
rect 14013 13345 14047 13379
rect 15669 13345 15703 13379
rect 16672 13345 16706 13379
rect 2605 13277 2639 13311
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 6469 13277 6503 13311
rect 6653 13277 6687 13311
rect 7849 13277 7883 13311
rect 8217 13277 8251 13311
rect 8769 13277 8803 13311
rect 8953 13277 8987 13311
rect 10241 13277 10275 13311
rect 10609 13277 10643 13311
rect 11529 13277 11563 13311
rect 13461 13277 13495 13311
rect 13645 13277 13679 13311
rect 15853 13277 15887 13311
rect 16405 13277 16439 13311
rect 5917 13209 5951 13243
rect 7113 13209 7147 13243
rect 13829 13209 13863 13243
rect 1961 13141 1995 13175
rect 7297 13141 7331 13175
rect 12909 13141 12943 13175
rect 15301 13141 15335 13175
rect 17969 13141 18003 13175
rect 3525 12937 3559 12971
rect 4629 12937 4663 12971
rect 13829 12937 13863 12971
rect 15669 12937 15703 12971
rect 16589 12937 16623 12971
rect 9689 12869 9723 12903
rect 10609 12869 10643 12903
rect 15577 12869 15611 12903
rect 3065 12801 3099 12835
rect 4077 12801 4111 12835
rect 10333 12801 10367 12835
rect 11161 12801 11195 12835
rect 11897 12801 11931 12835
rect 12081 12801 12115 12835
rect 16221 12801 16255 12835
rect 1409 12733 1443 12767
rect 2881 12733 2915 12767
rect 3985 12733 4019 12767
rect 4353 12733 4387 12767
rect 6837 12733 6871 12767
rect 7104 12733 7138 12767
rect 8309 12733 8343 12767
rect 10977 12733 11011 12767
rect 12265 12733 12299 12767
rect 12449 12733 12483 12767
rect 12716 12733 12750 12767
rect 14197 12733 14231 12767
rect 14464 12733 14498 12767
rect 16037 12733 16071 12767
rect 1676 12665 1710 12699
rect 3893 12665 3927 12699
rect 8554 12665 8588 12699
rect 11069 12665 11103 12699
rect 2789 12597 2823 12631
rect 8217 12597 8251 12631
rect 9781 12597 9815 12631
rect 10149 12597 10183 12631
rect 10241 12597 10275 12631
rect 11437 12597 11471 12631
rect 11805 12597 11839 12631
rect 12265 12597 12299 12631
rect 16129 12597 16163 12631
rect 3433 12393 3467 12427
rect 5549 12393 5583 12427
rect 7573 12393 7607 12427
rect 9045 12393 9079 12427
rect 9505 12393 9539 12427
rect 11069 12393 11103 12427
rect 12633 12393 12667 12427
rect 15301 12393 15335 12427
rect 15761 12393 15795 12427
rect 5908 12325 5942 12359
rect 9321 12325 9355 12359
rect 9956 12325 9990 12359
rect 14004 12325 14038 12359
rect 2053 12257 2087 12291
rect 2320 12257 2354 12291
rect 4169 12257 4203 12291
rect 4425 12257 4459 12291
rect 5641 12257 5675 12291
rect 7481 12257 7515 12291
rect 8585 12257 8619 12291
rect 9689 12257 9723 12291
rect 11161 12257 11195 12291
rect 11428 12257 11462 12291
rect 13001 12257 13035 12291
rect 13737 12257 13771 12291
rect 15669 12257 15703 12291
rect 7757 12189 7791 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 15853 12189 15887 12223
rect 15117 12121 15151 12155
rect 7021 12053 7055 12087
rect 7113 12053 7147 12087
rect 8769 12053 8803 12087
rect 12541 12053 12575 12087
rect 16221 12053 16255 12087
rect 1593 11849 1627 11883
rect 3617 11849 3651 11883
rect 4997 11849 5031 11883
rect 8033 11849 8067 11883
rect 8861 11849 8895 11883
rect 10149 11849 10183 11883
rect 11897 11849 11931 11883
rect 12449 11849 12483 11883
rect 10977 11781 11011 11815
rect 2237 11713 2271 11747
rect 3065 11713 3099 11747
rect 4169 11713 4203 11747
rect 4537 11713 4571 11747
rect 5641 11713 5675 11747
rect 8677 11713 8711 11747
rect 9321 11713 9355 11747
rect 9505 11713 9539 11747
rect 10609 11713 10643 11747
rect 10793 11713 10827 11747
rect 11437 11713 11471 11747
rect 11621 11713 11655 11747
rect 13001 11713 13035 11747
rect 14749 11713 14783 11747
rect 14933 11713 14967 11747
rect 2789 11645 2823 11679
rect 14013 11645 14047 11679
rect 15200 11645 15234 11679
rect 1501 11577 1535 11611
rect 2881 11577 2915 11611
rect 3525 11577 3559 11611
rect 3985 11577 4019 11611
rect 8493 11577 8527 11611
rect 9873 11577 9907 11611
rect 11345 11577 11379 11611
rect 14473 11577 14507 11611
rect 1961 11509 1995 11543
rect 2053 11509 2087 11543
rect 2421 11509 2455 11543
rect 4077 11509 4111 11543
rect 5365 11509 5399 11543
rect 5457 11509 5491 11543
rect 8401 11509 8435 11543
rect 9229 11509 9263 11543
rect 10057 11509 10091 11543
rect 10517 11509 10551 11543
rect 12817 11509 12851 11543
rect 12909 11509 12943 11543
rect 14105 11509 14139 11543
rect 14565 11509 14599 11543
rect 16313 11509 16347 11543
rect 2329 11305 2363 11339
rect 4721 11305 4755 11339
rect 9321 11305 9355 11339
rect 10977 11305 11011 11339
rect 11713 11305 11747 11339
rect 13277 11305 13311 11339
rect 14657 11305 14691 11339
rect 15301 11305 15335 11339
rect 1869 11237 1903 11271
rect 2789 11237 2823 11271
rect 9689 11237 9723 11271
rect 2145 11169 2179 11203
rect 2697 11169 2731 11203
rect 3157 11169 3191 11203
rect 5089 11169 5123 11203
rect 5549 11169 5583 11203
rect 6736 11169 6770 11203
rect 8208 11169 8242 11203
rect 12081 11169 12115 11203
rect 13645 11169 13679 11203
rect 2973 11101 3007 11135
rect 5181 11101 5215 11135
rect 5273 11101 5307 11135
rect 6469 11101 6503 11135
rect 7941 11101 7975 11135
rect 11621 11101 11655 11135
rect 12173 11101 12207 11135
rect 12265 11101 12299 11135
rect 13737 11101 13771 11135
rect 13921 11101 13955 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 4629 11033 4663 11067
rect 7849 11033 7883 11067
rect 9413 11033 9447 11067
rect 14289 11033 14323 11067
rect 5089 10761 5123 10795
rect 5917 10761 5951 10795
rect 10885 10761 10919 10795
rect 12725 10761 12759 10795
rect 15025 10761 15059 10795
rect 4721 10625 4755 10659
rect 4905 10625 4939 10659
rect 5641 10625 5675 10659
rect 6561 10625 6595 10659
rect 7481 10625 7515 10659
rect 9873 10625 9907 10659
rect 10701 10625 10735 10659
rect 11529 10625 11563 10659
rect 13277 10625 13311 10659
rect 15577 10625 15611 10659
rect 1777 10557 1811 10591
rect 2044 10557 2078 10591
rect 4169 10557 4203 10591
rect 5549 10557 5583 10591
rect 8309 10557 8343 10591
rect 10425 10557 10459 10591
rect 13185 10557 13219 10591
rect 13553 10557 13587 10591
rect 15485 10557 15519 10591
rect 3985 10489 4019 10523
rect 5457 10489 5491 10523
rect 6285 10489 6319 10523
rect 7205 10489 7239 10523
rect 7665 10489 7699 10523
rect 8576 10489 8610 10523
rect 11253 10489 11287 10523
rect 12081 10489 12115 10523
rect 13820 10489 13854 10523
rect 15393 10489 15427 10523
rect 3157 10421 3191 10455
rect 3801 10421 3835 10455
rect 4261 10421 4295 10455
rect 4629 10421 4663 10455
rect 6377 10421 6411 10455
rect 6837 10421 6871 10455
rect 7297 10421 7331 10455
rect 7941 10421 7975 10455
rect 9689 10421 9723 10455
rect 10057 10421 10091 10455
rect 10517 10421 10551 10455
rect 11345 10421 11379 10455
rect 11805 10421 11839 10455
rect 13093 10421 13127 10455
rect 14933 10421 14967 10455
rect 3709 10217 3743 10251
rect 5549 10217 5583 10251
rect 6377 10217 6411 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 10885 10217 10919 10251
rect 12909 10217 12943 10251
rect 14381 10217 14415 10251
rect 14657 10217 14691 10251
rect 14841 10217 14875 10251
rect 1961 10149 1995 10183
rect 4344 10149 4378 10183
rect 8493 10149 8527 10183
rect 9137 10149 9171 10183
rect 11796 10149 11830 10183
rect 13268 10149 13302 10183
rect 1685 10081 1719 10115
rect 2596 10081 2630 10115
rect 6745 10081 6779 10115
rect 7665 10081 7699 10115
rect 8677 10081 8711 10115
rect 10149 10081 10183 10115
rect 11437 10081 11471 10115
rect 13001 10081 13035 10115
rect 2329 10013 2363 10047
rect 4077 10013 4111 10047
rect 6101 10013 6135 10047
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 7757 10013 7791 10047
rect 7941 10013 7975 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 10333 10013 10367 10047
rect 10977 10013 11011 10047
rect 11069 10013 11103 10047
rect 11529 10013 11563 10047
rect 7297 9945 7331 9979
rect 8769 9945 8803 9979
rect 5457 9877 5491 9911
rect 6285 9877 6319 9911
rect 8217 9877 8251 9911
rect 10517 9877 10551 9911
rect 8217 9673 8251 9707
rect 13645 9673 13679 9707
rect 3985 9605 4019 9639
rect 10149 9605 10183 9639
rect 10241 9605 10275 9639
rect 11345 9605 11379 9639
rect 12449 9605 12483 9639
rect 2145 9537 2179 9571
rect 4537 9537 4571 9571
rect 5549 9537 5583 9571
rect 10793 9537 10827 9571
rect 11989 9537 12023 9571
rect 12081 9537 12115 9571
rect 13093 9537 13127 9571
rect 14289 9537 14323 9571
rect 1961 9469 1995 9503
rect 4353 9469 4387 9503
rect 4445 9469 4479 9503
rect 5917 9469 5951 9503
rect 6837 9469 6871 9503
rect 8769 9469 8803 9503
rect 9036 9469 9070 9503
rect 12909 9469 12943 9503
rect 7104 9401 7138 9435
rect 10701 9401 10735 9435
rect 12817 9401 12851 9435
rect 13369 9401 13403 9435
rect 14105 9401 14139 9435
rect 4905 9333 4939 9367
rect 5273 9333 5307 9367
rect 5365 9333 5399 9367
rect 5733 9333 5767 9367
rect 8309 9333 8343 9367
rect 8493 9333 8527 9367
rect 10609 9333 10643 9367
rect 11161 9333 11195 9367
rect 11529 9333 11563 9367
rect 11897 9333 11931 9367
rect 13461 9333 13495 9367
rect 14013 9333 14047 9367
rect 1869 9129 1903 9163
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 5733 9129 5767 9163
rect 7665 9129 7699 9163
rect 8125 9129 8159 9163
rect 8769 9129 8803 9163
rect 11161 9129 11195 9163
rect 11989 9129 12023 9163
rect 12265 9129 12299 9163
rect 13093 9129 13127 9163
rect 13737 9129 13771 9163
rect 2237 8993 2271 9027
rect 3157 8993 3191 9027
rect 4620 8993 4654 9027
rect 6081 8993 6115 9027
rect 8033 8993 8067 9027
rect 8677 8993 8711 9027
rect 9137 8993 9171 9027
rect 9956 8993 9990 9027
rect 11529 8993 11563 9027
rect 12449 8993 12483 9027
rect 13645 8993 13679 9027
rect 2513 8925 2547 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 4353 8925 4387 8959
rect 5825 8925 5859 8959
rect 8217 8925 8251 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 9689 8925 9723 8959
rect 11621 8925 11655 8959
rect 11805 8925 11839 8959
rect 13829 8925 13863 8959
rect 7205 8857 7239 8891
rect 12541 8857 12575 8891
rect 7297 8789 7331 8823
rect 8493 8789 8527 8823
rect 11069 8789 11103 8823
rect 13277 8789 13311 8823
rect 3525 8585 3559 8619
rect 4905 8585 4939 8619
rect 5733 8585 5767 8619
rect 9229 8585 9263 8619
rect 10333 8585 10367 8619
rect 7665 8517 7699 8551
rect 8401 8517 8435 8551
rect 10701 8517 10735 8551
rect 11529 8517 11563 8551
rect 1869 8449 1903 8483
rect 4077 8449 4111 8483
rect 4445 8449 4479 8483
rect 5549 8449 5583 8483
rect 6285 8449 6319 8483
rect 7389 8449 7423 8483
rect 8861 8449 8895 8483
rect 9045 8449 9079 8483
rect 9781 8449 9815 8483
rect 10057 8449 10091 8483
rect 11253 8449 11287 8483
rect 11805 8449 11839 8483
rect 12449 8449 12483 8483
rect 13369 8449 13403 8483
rect 13645 8449 13679 8483
rect 16221 8449 16255 8483
rect 2136 8381 2170 8415
rect 5365 8381 5399 8415
rect 6101 8381 6135 8415
rect 7297 8381 7331 8415
rect 7849 8381 7883 8415
rect 9597 8381 9631 8415
rect 10517 8381 10551 8415
rect 11161 8381 11195 8415
rect 14197 8381 14231 8415
rect 3985 8313 4019 8347
rect 4629 8313 4663 8347
rect 5273 8313 5307 8347
rect 6193 8313 6227 8347
rect 8125 8313 8159 8347
rect 9689 8313 9723 8347
rect 12633 8313 12667 8347
rect 13185 8313 13219 8347
rect 13277 8313 13311 8347
rect 14442 8313 14476 8347
rect 16037 8313 16071 8347
rect 3249 8245 3283 8279
rect 3341 8245 3375 8279
rect 3893 8245 3927 8279
rect 6653 8245 6687 8279
rect 6837 8245 6871 8279
rect 7205 8245 7239 8279
rect 8217 8245 8251 8279
rect 8769 8245 8803 8279
rect 11069 8245 11103 8279
rect 12817 8245 12851 8279
rect 15577 8245 15611 8279
rect 15669 8245 15703 8279
rect 16129 8245 16163 8279
rect 2789 8041 2823 8075
rect 3249 8041 3283 8075
rect 4169 8041 4203 8075
rect 5825 8041 5859 8075
rect 6009 8041 6043 8075
rect 7481 8041 7515 8075
rect 14565 8041 14599 8075
rect 15301 8041 15335 8075
rect 4712 7973 4746 8007
rect 10692 7973 10726 8007
rect 12900 7973 12934 8007
rect 15761 7973 15795 8007
rect 1409 7905 1443 7939
rect 1676 7905 1710 7939
rect 3341 7905 3375 7939
rect 6561 7905 6595 7939
rect 7389 7905 7423 7939
rect 8033 7905 8067 7939
rect 10425 7905 10459 7939
rect 12633 7905 12667 7939
rect 14473 7905 14507 7939
rect 15117 7905 15151 7939
rect 15669 7905 15703 7939
rect 3433 7837 3467 7871
rect 4445 7837 4479 7871
rect 6653 7837 6687 7871
rect 6837 7837 6871 7871
rect 7573 7837 7607 7871
rect 14657 7837 14691 7871
rect 15945 7837 15979 7871
rect 3801 7769 3835 7803
rect 14105 7769 14139 7803
rect 2881 7701 2915 7735
rect 4261 7701 4295 7735
rect 6193 7701 6227 7735
rect 7021 7701 7055 7735
rect 7849 7701 7883 7735
rect 8861 7701 8895 7735
rect 9137 7701 9171 7735
rect 11805 7701 11839 7735
rect 14013 7701 14047 7735
rect 3525 7497 3559 7531
rect 4353 7497 4387 7531
rect 5365 7497 5399 7531
rect 8861 7497 8895 7531
rect 12265 7497 12299 7531
rect 13277 7497 13311 7531
rect 15025 7497 15059 7531
rect 2237 7429 2271 7463
rect 9229 7429 9263 7463
rect 11345 7429 11379 7463
rect 12449 7429 12483 7463
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 4077 7361 4111 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 9873 7361 9907 7395
rect 10057 7361 10091 7395
rect 13001 7361 13035 7395
rect 13737 7361 13771 7395
rect 13921 7361 13955 7395
rect 5733 7293 5767 7327
rect 6285 7293 6319 7327
rect 7481 7293 7515 7327
rect 11529 7293 11563 7327
rect 12909 7293 12943 7327
rect 13645 7293 13679 7327
rect 15301 7293 15335 7327
rect 15568 7293 15602 7327
rect 2697 7225 2731 7259
rect 3157 7225 3191 7259
rect 3985 7225 4019 7259
rect 7748 7225 7782 7259
rect 12817 7225 12851 7259
rect 2329 7157 2363 7191
rect 3893 7157 3927 7191
rect 4537 7157 4571 7191
rect 4813 7157 4847 7191
rect 5549 7157 5583 7191
rect 5917 7157 5951 7191
rect 9413 7157 9447 7191
rect 9781 7157 9815 7191
rect 12081 7157 12115 7191
rect 16681 7157 16715 7191
rect 2421 6953 2455 6987
rect 3617 6953 3651 6987
rect 4077 6953 4111 6987
rect 4537 6953 4571 6987
rect 7849 6953 7883 6987
rect 8309 6953 8343 6987
rect 9229 6953 9263 6987
rect 10517 6953 10551 6987
rect 13829 6953 13863 6987
rect 14289 6953 14323 6987
rect 4445 6885 4479 6919
rect 6009 6885 6043 6919
rect 10057 6885 10091 6919
rect 11152 6885 11186 6919
rect 2513 6817 2547 6851
rect 3525 6817 3559 6851
rect 6736 6817 6770 6851
rect 13645 6817 13679 6851
rect 14381 6817 14415 6851
rect 2697 6749 2731 6783
rect 3065 6749 3099 6783
rect 3801 6749 3835 6783
rect 4721 6749 4755 6783
rect 6101 6749 6135 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 8401 6749 8435 6783
rect 8493 6749 8527 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 10885 6749 10919 6783
rect 14565 6749 14599 6783
rect 14749 6749 14783 6783
rect 2053 6681 2087 6715
rect 5273 6681 5307 6715
rect 9689 6681 9723 6715
rect 3157 6613 3191 6647
rect 5641 6613 5675 6647
rect 7941 6613 7975 6647
rect 9413 6613 9447 6647
rect 12265 6613 12299 6647
rect 13921 6613 13955 6647
rect 3249 6409 3283 6443
rect 7021 6409 7055 6443
rect 12449 6409 12483 6443
rect 6653 6341 6687 6375
rect 11989 6341 12023 6375
rect 15209 6341 15243 6375
rect 3985 6273 4019 6307
rect 4813 6273 4847 6307
rect 4997 6273 5031 6307
rect 7665 6273 7699 6307
rect 8953 6273 8987 6307
rect 9137 6273 9171 6307
rect 11345 6273 11379 6307
rect 13093 6273 13127 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 1869 6205 1903 6239
rect 4721 6205 4755 6239
rect 5273 6205 5307 6239
rect 5540 6205 5574 6239
rect 9321 6205 9355 6239
rect 11161 6205 11195 6239
rect 11253 6205 11287 6239
rect 12817 6205 12851 6239
rect 13829 6205 13863 6239
rect 14096 6205 14130 6239
rect 16405 6205 16439 6239
rect 2136 6137 2170 6171
rect 8861 6137 8895 6171
rect 9588 6137 9622 6171
rect 12909 6137 12943 6171
rect 15669 6137 15703 6171
rect 16672 6137 16706 6171
rect 3433 6069 3467 6103
rect 3801 6069 3835 6103
rect 3893 6069 3927 6103
rect 4353 6069 4387 6103
rect 7389 6069 7423 6103
rect 7481 6069 7515 6103
rect 7849 6069 7883 6103
rect 8493 6069 8527 6103
rect 10701 6069 10735 6103
rect 10793 6069 10827 6103
rect 12173 6069 12207 6103
rect 15301 6069 15335 6103
rect 17785 6069 17819 6103
rect 3157 5865 3191 5899
rect 3617 5865 3651 5899
rect 6101 5865 6135 5899
rect 7941 5865 7975 5899
rect 8309 5865 8343 5899
rect 9137 5865 9171 5899
rect 9229 5865 9263 5899
rect 11069 5865 11103 5899
rect 14105 5865 14139 5899
rect 14473 5865 14507 5899
rect 17417 5865 17451 5899
rect 17969 5865 18003 5899
rect 6736 5797 6770 5831
rect 9945 5797 9979 5831
rect 15761 5797 15795 5831
rect 17877 5797 17911 5831
rect 1777 5729 1811 5763
rect 2044 5729 2078 5763
rect 4721 5729 4755 5763
rect 4988 5729 5022 5763
rect 11529 5729 11563 5763
rect 12633 5729 12667 5763
rect 12900 5729 12934 5763
rect 14565 5729 14599 5763
rect 14933 5729 14967 5763
rect 16304 5729 16338 5763
rect 6469 5661 6503 5695
rect 8401 5661 8435 5695
rect 8493 5661 8527 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 11621 5661 11655 5695
rect 11805 5661 11839 5695
rect 14657 5661 14691 5695
rect 16037 5661 16071 5695
rect 18061 5661 18095 5695
rect 7849 5593 7883 5627
rect 11161 5593 11195 5627
rect 4169 5525 4203 5559
rect 8769 5525 8803 5559
rect 14013 5525 14047 5559
rect 17509 5525 17543 5559
rect 3709 5321 3743 5355
rect 4629 5321 4663 5355
rect 5917 5321 5951 5355
rect 8861 5321 8895 5355
rect 11161 5321 11195 5355
rect 16865 5321 16899 5355
rect 17785 5321 17819 5355
rect 8953 5253 8987 5287
rect 10333 5253 10367 5287
rect 4261 5185 4295 5219
rect 5273 5185 5307 5219
rect 6561 5185 6595 5219
rect 10977 5185 11011 5219
rect 11621 5185 11655 5219
rect 11805 5185 11839 5219
rect 15117 5185 15151 5219
rect 15485 5185 15519 5219
rect 17509 5185 17543 5219
rect 1869 5117 1903 5151
rect 2136 5117 2170 5151
rect 5825 5117 5859 5151
rect 7481 5117 7515 5151
rect 7748 5117 7782 5151
rect 13093 5117 13127 5151
rect 14933 5117 14967 5151
rect 19073 5117 19107 5151
rect 3525 5049 3559 5083
rect 4169 5049 4203 5083
rect 5641 5049 5675 5083
rect 9965 5049 9999 5083
rect 11529 5049 11563 5083
rect 13360 5049 13394 5083
rect 15025 5049 15059 5083
rect 15752 5049 15786 5083
rect 17325 5049 17359 5083
rect 19349 5049 19383 5083
rect 3249 4981 3283 5015
rect 3433 4981 3467 5015
rect 4077 4981 4111 5015
rect 4997 4981 5031 5015
rect 5089 4981 5123 5015
rect 6285 4981 6319 5015
rect 6377 4981 6411 5015
rect 10149 4981 10183 5015
rect 10701 4981 10735 5015
rect 10793 4981 10827 5015
rect 11989 4981 12023 5015
rect 12265 4981 12299 5015
rect 14473 4981 14507 5015
rect 14565 4981 14599 5015
rect 16957 4981 16991 5015
rect 17417 4981 17451 5015
rect 18061 4981 18095 5015
rect 2053 4777 2087 4811
rect 3433 4777 3467 4811
rect 6009 4777 6043 4811
rect 7297 4777 7331 4811
rect 8125 4777 8159 4811
rect 10333 4777 10367 4811
rect 11253 4777 11287 4811
rect 12449 4777 12483 4811
rect 12909 4777 12943 4811
rect 13737 4777 13771 4811
rect 15669 4777 15703 4811
rect 16129 4777 16163 4811
rect 16589 4777 16623 4811
rect 17325 4777 17359 4811
rect 1777 4709 1811 4743
rect 3341 4709 3375 4743
rect 15761 4709 15795 4743
rect 17417 4709 17451 4743
rect 1501 4641 1535 4675
rect 2421 4641 2455 4675
rect 2513 4641 2547 4675
rect 4629 4641 4663 4675
rect 4896 4641 4930 4675
rect 7665 4641 7699 4675
rect 8493 4641 8527 4675
rect 10241 4641 10275 4675
rect 11621 4641 11655 4675
rect 11713 4641 11747 4675
rect 13277 4641 13311 4675
rect 14105 4641 14139 4675
rect 16497 4641 16531 4675
rect 19993 4641 20027 4675
rect 2697 4573 2731 4607
rect 3617 4573 3651 4607
rect 7757 4573 7791 4607
rect 7941 4573 7975 4607
rect 8585 4573 8619 4607
rect 8769 4573 8803 4607
rect 10425 4573 10459 4607
rect 11805 4573 11839 4607
rect 12541 4573 12575 4607
rect 12725 4573 12759 4607
rect 13369 4573 13403 4607
rect 13553 4573 13587 4607
rect 14197 4573 14231 4607
rect 14381 4573 14415 4607
rect 15853 4573 15887 4607
rect 16773 4573 16807 4607
rect 17509 4573 17543 4607
rect 2973 4505 3007 4539
rect 9873 4505 9907 4539
rect 12081 4505 12115 4539
rect 6929 4437 6963 4471
rect 7113 4437 7147 4471
rect 10793 4437 10827 4471
rect 11069 4437 11103 4471
rect 14657 4437 14691 4471
rect 15301 4437 15335 4471
rect 16957 4437 16991 4471
rect 20177 4437 20211 4471
rect 3249 4233 3283 4267
rect 6837 4233 6871 4267
rect 7205 4233 7239 4267
rect 8401 4233 8435 4267
rect 10149 4233 10183 4267
rect 11161 4233 11195 4267
rect 11989 4233 12023 4267
rect 15025 4233 15059 4267
rect 12633 4165 12667 4199
rect 6101 4097 6135 4131
rect 8033 4097 8067 4131
rect 8217 4097 8251 4131
rect 9045 4097 9079 4131
rect 10609 4097 10643 4131
rect 10701 4097 10735 4131
rect 11713 4097 11747 4131
rect 12817 4097 12851 4131
rect 1869 4029 1903 4063
rect 3341 4029 3375 4063
rect 3597 4029 3631 4063
rect 5365 4029 5399 4063
rect 6009 4029 6043 4063
rect 7941 4029 7975 4063
rect 11069 4029 11103 4063
rect 11621 4029 11655 4063
rect 12173 4029 12207 4063
rect 13645 4029 13679 4063
rect 17141 4029 17175 4063
rect 2114 3961 2148 3995
rect 7021 3961 7055 3995
rect 8861 3961 8895 3995
rect 9229 3961 9263 3995
rect 11529 3961 11563 3995
rect 13912 3961 13946 3995
rect 17417 3961 17451 3995
rect 4721 3893 4755 3927
rect 5549 3893 5583 3927
rect 5917 3893 5951 3927
rect 6377 3893 6411 3927
rect 7389 3893 7423 3927
rect 7573 3893 7607 3927
rect 8769 3893 8803 3927
rect 9413 3893 9447 3927
rect 10517 3893 10551 3927
rect 3157 3689 3191 3723
rect 5917 3689 5951 3723
rect 6009 3689 6043 3723
rect 7205 3689 7239 3723
rect 7665 3689 7699 3723
rect 8953 3689 8987 3723
rect 9781 3689 9815 3723
rect 9873 3689 9907 3723
rect 10333 3689 10367 3723
rect 10701 3689 10735 3723
rect 11529 3689 11563 3723
rect 13921 3689 13955 3723
rect 1952 3621 1986 3655
rect 4782 3621 4816 3655
rect 8125 3621 8159 3655
rect 10241 3621 10275 3655
rect 12173 3621 12207 3655
rect 16037 3621 16071 3655
rect 1685 3553 1719 3587
rect 3525 3553 3559 3587
rect 3617 3553 3651 3587
rect 4537 3553 4571 3587
rect 6377 3553 6411 3587
rect 6469 3553 6503 3587
rect 8033 3553 8067 3587
rect 8861 3553 8895 3587
rect 9413 3553 9447 3587
rect 11069 3553 11103 3587
rect 3709 3485 3743 3519
rect 6561 3485 6595 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 8217 3485 8251 3519
rect 9045 3485 9079 3519
rect 10425 3485 10459 3519
rect 11161 3485 11195 3519
rect 11345 3485 11379 3519
rect 12532 3553 12566 3587
rect 14289 3553 14323 3587
rect 15485 3553 15519 3587
rect 18061 3553 18095 3587
rect 12265 3485 12299 3519
rect 14381 3485 14415 3519
rect 14473 3485 14507 3519
rect 15761 3485 15795 3519
rect 6837 3417 6871 3451
rect 8493 3417 8527 3451
rect 12173 3417 12207 3451
rect 13645 3417 13679 3451
rect 1501 3349 1535 3383
rect 3065 3349 3099 3383
rect 13829 3349 13863 3383
rect 18245 3349 18279 3383
rect 2789 3145 2823 3179
rect 3617 3145 3651 3179
rect 4721 3145 4755 3179
rect 8953 3145 8987 3179
rect 10425 3145 10459 3179
rect 11897 3145 11931 3179
rect 13829 3145 13863 3179
rect 18245 3145 18279 3179
rect 12449 3077 12483 3111
rect 16221 3077 16255 3111
rect 17417 3077 17451 3111
rect 18429 3077 18463 3111
rect 18797 3077 18831 3111
rect 19625 3077 19659 3111
rect 2421 3009 2455 3043
rect 2605 3009 2639 3043
rect 3341 3009 3375 3043
rect 4169 3009 4203 3043
rect 5365 3009 5399 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 6377 3009 6411 3043
rect 7573 3009 7607 3043
rect 9045 3009 9079 3043
rect 10517 3009 10551 3043
rect 13001 3009 13035 3043
rect 14289 3009 14323 3043
rect 19809 3009 19843 3043
rect 20177 3009 20211 3043
rect 2329 2941 2363 2975
rect 5089 2941 5123 2975
rect 5181 2941 5215 2975
rect 7021 2941 7055 2975
rect 7840 2941 7874 2975
rect 9301 2941 9335 2975
rect 13277 2941 13311 2975
rect 14013 2941 14047 2975
rect 14565 2941 14599 2975
rect 14933 2941 14967 2975
rect 15301 2941 15335 2975
rect 15669 2941 15703 2975
rect 16037 2941 16071 2975
rect 16405 2941 16439 2975
rect 16773 2941 16807 2975
rect 17233 2941 17267 2975
rect 17601 2941 17635 2975
rect 18061 2941 18095 2975
rect 18613 2941 18647 2975
rect 19073 2941 19107 2975
rect 19441 2941 19475 2975
rect 20361 2941 20395 2975
rect 1685 2873 1719 2907
rect 3985 2873 4019 2907
rect 4445 2873 4479 2907
rect 5917 2873 5951 2907
rect 6837 2873 6871 2907
rect 7297 2873 7331 2907
rect 10762 2873 10796 2907
rect 12909 2873 12943 2907
rect 13553 2873 13587 2907
rect 1593 2805 1627 2839
rect 1961 2805 1995 2839
rect 3157 2805 3191 2839
rect 3249 2805 3283 2839
rect 4077 2805 4111 2839
rect 5549 2805 5583 2839
rect 12817 2805 12851 2839
rect 14749 2805 14783 2839
rect 15117 2805 15151 2839
rect 15485 2805 15519 2839
rect 15853 2805 15887 2839
rect 16589 2805 16623 2839
rect 16957 2805 16991 2839
rect 17785 2805 17819 2839
rect 19257 2805 19291 2839
rect 20545 2805 20579 2839
rect 1409 2601 1443 2635
rect 1869 2601 1903 2635
rect 2237 2601 2271 2635
rect 2605 2601 2639 2635
rect 3709 2601 3743 2635
rect 4721 2601 4755 2635
rect 5549 2601 5583 2635
rect 6377 2601 6411 2635
rect 8033 2601 8067 2635
rect 10333 2601 10367 2635
rect 10793 2601 10827 2635
rect 10977 2601 11011 2635
rect 11437 2601 11471 2635
rect 11897 2601 11931 2635
rect 14381 2601 14415 2635
rect 15209 2601 15243 2635
rect 15945 2601 15979 2635
rect 16129 2601 16163 2635
rect 16681 2601 16715 2635
rect 17141 2601 17175 2635
rect 17417 2601 17451 2635
rect 17969 2601 18003 2635
rect 18981 2601 19015 2635
rect 1777 2533 1811 2567
rect 7941 2533 7975 2567
rect 8493 2533 8527 2567
rect 11345 2533 11379 2567
rect 4997 2465 5031 2499
rect 5917 2465 5951 2499
rect 7665 2465 7699 2499
rect 8401 2465 8435 2499
rect 10425 2465 10459 2499
rect 12633 2465 12667 2499
rect 12909 2465 12943 2499
rect 13185 2465 13219 2499
rect 13553 2465 13587 2499
rect 13921 2465 13955 2499
rect 15577 2465 15611 2499
rect 2053 2397 2087 2431
rect 2697 2397 2731 2431
rect 2789 2397 2823 2431
rect 6009 2397 6043 2431
rect 6193 2397 6227 2431
rect 8585 2397 8619 2431
rect 10609 2397 10643 2431
rect 11529 2397 11563 2431
rect 3249 2329 3283 2363
rect 9965 2329 9999 2363
rect 3065 2261 3099 2295
rect 5181 2261 5215 2295
rect 5365 2261 5399 2295
rect 13369 2261 13403 2295
rect 13737 2261 13771 2295
rect 14105 2261 14139 2295
rect 15761 2261 15795 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2774 20584 2780 20596
rect 1995 20556 2780 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 6549 20587 6607 20593
rect 6549 20553 6561 20587
rect 6595 20584 6607 20587
rect 7098 20584 7104 20596
rect 6595 20556 7104 20584
rect 6595 20553 6607 20556
rect 6549 20547 6607 20553
rect 2317 20519 2375 20525
rect 2317 20485 2329 20519
rect 2363 20516 2375 20519
rect 2866 20516 2872 20528
rect 2363 20488 2872 20516
rect 2363 20485 2375 20488
rect 2317 20479 2375 20485
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 6564 20516 6592 20547
rect 7098 20544 7104 20556
rect 7156 20544 7162 20596
rect 7742 20544 7748 20596
rect 7800 20584 7806 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7800 20556 8217 20584
rect 7800 20544 7806 20556
rect 8205 20553 8217 20556
rect 8251 20584 8263 20587
rect 10778 20584 10784 20596
rect 8251 20556 10784 20584
rect 8251 20553 8263 20556
rect 8205 20547 8263 20553
rect 10778 20544 10784 20556
rect 10836 20544 10842 20596
rect 6104 20488 6592 20516
rect 6104 20457 6132 20488
rect 6089 20451 6147 20457
rect 6089 20417 6101 20451
rect 6135 20417 6147 20451
rect 6270 20448 6276 20460
rect 6231 20420 6276 20448
rect 6089 20411 6147 20417
rect 6270 20408 6276 20420
rect 6328 20408 6334 20460
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 2130 20380 2136 20392
rect 2091 20352 2136 20380
rect 2130 20340 2136 20352
rect 2188 20340 2194 20392
rect 4522 20340 4528 20392
rect 4580 20380 4586 20392
rect 4985 20383 5043 20389
rect 4985 20380 4997 20383
rect 4580 20352 4997 20380
rect 4580 20340 4586 20352
rect 4985 20349 4997 20352
rect 5031 20380 5043 20383
rect 8938 20380 8944 20392
rect 5031 20352 8944 20380
rect 5031 20349 5043 20352
rect 4985 20343 5043 20349
rect 8938 20340 8944 20352
rect 8996 20340 9002 20392
rect 5445 20315 5503 20321
rect 5445 20281 5457 20315
rect 5491 20312 5503 20315
rect 5491 20284 6040 20312
rect 5491 20281 5503 20284
rect 5445 20275 5503 20281
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 6012 20253 6040 20284
rect 6822 20272 6828 20324
rect 6880 20312 6886 20324
rect 7377 20315 7435 20321
rect 7377 20312 7389 20315
rect 6880 20284 7389 20312
rect 6880 20272 6886 20284
rect 7377 20281 7389 20284
rect 7423 20281 7435 20315
rect 7377 20275 7435 20281
rect 13262 20272 13268 20324
rect 13320 20312 13326 20324
rect 21818 20312 21824 20324
rect 13320 20284 21824 20312
rect 13320 20272 13326 20284
rect 21818 20272 21824 20284
rect 21876 20272 21882 20324
rect 5629 20247 5687 20253
rect 5629 20244 5641 20247
rect 5592 20216 5641 20244
rect 5592 20204 5598 20216
rect 5629 20213 5641 20216
rect 5675 20213 5687 20247
rect 5629 20207 5687 20213
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6546 20244 6552 20256
rect 6043 20216 6552 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 7064 20216 7113 20244
rect 7064 20204 7070 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 9582 20244 9588 20256
rect 9543 20216 9588 20244
rect 7101 20207 7159 20213
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 13722 20204 13728 20256
rect 13780 20244 13786 20256
rect 19518 20244 19524 20256
rect 13780 20216 19524 20244
rect 13780 20204 13786 20216
rect 19518 20204 19524 20216
rect 19576 20204 19582 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 4522 20040 4528 20052
rect 4483 20012 4528 20040
rect 4522 20000 4528 20012
rect 4580 20000 4586 20052
rect 6822 20040 6828 20052
rect 6783 20012 6828 20040
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 6917 20043 6975 20049
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 6963 20012 7297 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 7742 20040 7748 20052
rect 7703 20012 7748 20040
rect 7285 20003 7343 20009
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 8294 20000 8300 20052
rect 8352 20040 8358 20052
rect 9582 20040 9588 20052
rect 8352 20012 9588 20040
rect 8352 20000 8358 20012
rect 9582 20000 9588 20012
rect 9640 20040 9646 20052
rect 10045 20043 10103 20049
rect 10045 20040 10057 20043
rect 9640 20012 10057 20040
rect 9640 20000 9646 20012
rect 10045 20009 10057 20012
rect 10091 20009 10103 20043
rect 10045 20003 10103 20009
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 10597 20043 10655 20049
rect 10597 20040 10609 20043
rect 10183 20012 10609 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 10597 20009 10609 20012
rect 10643 20040 10655 20043
rect 12618 20040 12624 20052
rect 10643 20012 12624 20040
rect 10643 20009 10655 20012
rect 10597 20003 10655 20009
rect 12618 20000 12624 20012
rect 12676 20000 12682 20052
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13078 20040 13084 20052
rect 12851 20012 13084 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 13262 20040 13268 20052
rect 13223 20012 13268 20040
rect 13262 20000 13268 20012
rect 13320 20000 13326 20052
rect 13722 20040 13728 20052
rect 13683 20012 13728 20040
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20009 14795 20043
rect 14737 20003 14795 20009
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 17218 20040 17224 20052
rect 16531 20012 17224 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 8662 19972 8668 19984
rect 1780 19944 8668 19972
rect 1780 19913 1808 19944
rect 8662 19932 8668 19944
rect 8720 19932 8726 19984
rect 11974 19932 11980 19984
rect 12032 19972 12038 19984
rect 14752 19972 14780 20003
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 21358 19972 21364 19984
rect 12032 19944 13584 19972
rect 14752 19944 21364 19972
rect 12032 19932 12038 19944
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19873 1455 19907
rect 1397 19867 1455 19873
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 2222 19904 2228 19916
rect 2183 19876 2228 19904
rect 1765 19867 1823 19873
rect 1412 19836 1440 19867
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 3513 19907 3571 19913
rect 3513 19873 3525 19907
rect 3559 19904 3571 19907
rect 4154 19904 4160 19916
rect 3559 19876 4160 19904
rect 3559 19873 3571 19876
rect 3513 19867 3571 19873
rect 4154 19864 4160 19876
rect 4212 19904 4218 19916
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 4212 19876 4445 19904
rect 4212 19864 4218 19876
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 5252 19907 5310 19913
rect 5252 19873 5264 19907
rect 5298 19904 5310 19907
rect 6270 19904 6276 19916
rect 5298 19876 6276 19904
rect 5298 19873 5310 19876
rect 5252 19867 5310 19873
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 7006 19864 7012 19916
rect 7064 19904 7070 19916
rect 7653 19907 7711 19913
rect 7653 19904 7665 19907
rect 7064 19876 7665 19904
rect 7064 19864 7070 19876
rect 7653 19873 7665 19876
rect 7699 19873 7711 19907
rect 7653 19867 7711 19873
rect 8380 19907 8438 19913
rect 8380 19873 8392 19907
rect 8426 19904 8438 19907
rect 9306 19904 9312 19916
rect 8426 19876 9312 19904
rect 8426 19873 8438 19876
rect 8380 19867 8438 19873
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19904 11023 19907
rect 11054 19904 11060 19916
rect 11011 19876 11060 19904
rect 11011 19873 11023 19876
rect 10965 19867 11023 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11232 19907 11290 19913
rect 11232 19873 11244 19907
rect 11278 19904 11290 19907
rect 12158 19904 12164 19916
rect 11278 19876 12164 19904
rect 11278 19873 11290 19876
rect 11232 19867 11290 19873
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13556 19913 13584 19944
rect 21358 19932 21364 19944
rect 21416 19932 21422 19984
rect 13081 19907 13139 19913
rect 13081 19873 13093 19907
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 13541 19907 13599 19913
rect 13541 19873 13553 19907
rect 13587 19904 13599 19907
rect 13909 19907 13967 19913
rect 13909 19904 13921 19907
rect 13587 19876 13921 19904
rect 13587 19873 13599 19876
rect 13541 19867 13599 19873
rect 13909 19873 13921 19876
rect 13955 19873 13967 19907
rect 14553 19907 14611 19913
rect 14553 19904 14565 19907
rect 13909 19867 13967 19873
rect 14200 19876 14565 19904
rect 2409 19839 2467 19845
rect 2409 19836 2421 19839
rect 1412 19808 2421 19836
rect 2409 19805 2421 19808
rect 2455 19805 2467 19839
rect 2409 19799 2467 19805
rect 2774 19796 2780 19848
rect 2832 19836 2838 19848
rect 3605 19839 3663 19845
rect 3605 19836 3617 19839
rect 2832 19808 3617 19836
rect 2832 19796 2838 19808
rect 3605 19805 3617 19808
rect 3651 19805 3663 19839
rect 3605 19799 3663 19805
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 4798 19836 4804 19848
rect 4755 19808 4804 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 4890 19796 4896 19848
rect 4948 19836 4954 19848
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 4948 19808 4997 19836
rect 4948 19796 4954 19808
rect 4985 19805 4997 19808
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19836 7159 19839
rect 7374 19836 7380 19848
rect 7147 19808 7380 19836
rect 7147 19805 7159 19808
rect 7101 19799 7159 19805
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 7929 19839 7987 19845
rect 7929 19805 7941 19839
rect 7975 19805 7987 19839
rect 8110 19836 8116 19848
rect 8071 19808 8116 19836
rect 7929 19799 7987 19805
rect 2866 19728 2872 19780
rect 2924 19768 2930 19780
rect 4065 19771 4123 19777
rect 4065 19768 4077 19771
rect 2924 19740 4077 19768
rect 2924 19728 2930 19740
rect 4065 19737 4077 19740
rect 4111 19737 4123 19771
rect 4065 19731 4123 19737
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 6457 19771 6515 19777
rect 6457 19768 6469 19771
rect 6236 19740 6469 19768
rect 6236 19728 6242 19740
rect 6457 19737 6469 19740
rect 6503 19737 6515 19771
rect 6457 19731 6515 19737
rect 6362 19700 6368 19712
rect 6323 19672 6368 19700
rect 6362 19660 6368 19672
rect 6420 19660 6426 19712
rect 7282 19660 7288 19712
rect 7340 19700 7346 19712
rect 7944 19700 7972 19799
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 10321 19839 10379 19845
rect 10321 19805 10333 19839
rect 10367 19805 10379 19839
rect 13096 19836 13124 19867
rect 10321 19799 10379 19805
rect 12452 19808 13124 19836
rect 10336 19712 10364 19799
rect 12452 19712 12480 19808
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 7340 19672 9505 19700
rect 7340 19660 7346 19672
rect 9493 19669 9505 19672
rect 9539 19669 9551 19703
rect 9674 19700 9680 19712
rect 9635 19672 9680 19700
rect 9493 19663 9551 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 10318 19700 10324 19712
rect 10231 19672 10324 19700
rect 10318 19660 10324 19672
rect 10376 19700 10382 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 10376 19672 12357 19700
rect 10376 19660 10382 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 12345 19663 12403 19669
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 12492 19672 12537 19700
rect 12492 19660 12498 19672
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 14200 19700 14228 19876
rect 14553 19873 14565 19876
rect 14599 19873 14611 19907
rect 16301 19907 16359 19913
rect 16301 19904 16313 19907
rect 14553 19867 14611 19873
rect 16132 19876 16313 19904
rect 14369 19703 14427 19709
rect 14369 19700 14381 19703
rect 12952 19672 14381 19700
rect 12952 19660 12958 19672
rect 14369 19669 14381 19672
rect 14415 19669 14427 19703
rect 14369 19663 14427 19669
rect 14550 19660 14556 19712
rect 14608 19700 14614 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 14608 19672 14933 19700
rect 14608 19660 14614 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16132 19709 16160 19876
rect 16301 19873 16313 19876
rect 16347 19873 16359 19907
rect 16301 19867 16359 19873
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 16632 19876 16681 19904
rect 16632 19864 16638 19876
rect 16669 19873 16681 19876
rect 16715 19904 16727 19907
rect 17037 19907 17095 19913
rect 17037 19904 17049 19907
rect 16715 19876 17049 19904
rect 16715 19873 16727 19876
rect 16669 19867 16727 19873
rect 17037 19873 17049 19876
rect 17083 19873 17095 19907
rect 17037 19867 17095 19873
rect 16853 19771 16911 19777
rect 16853 19737 16865 19771
rect 16899 19768 16911 19771
rect 20898 19768 20904 19780
rect 16899 19740 20904 19768
rect 16899 19737 16911 19740
rect 16853 19731 16911 19737
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 16080 19672 16129 19700
rect 16080 19660 16086 19672
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 16117 19663 16175 19669
rect 18693 19703 18751 19709
rect 18693 19669 18705 19703
rect 18739 19700 18751 19703
rect 18782 19700 18788 19712
rect 18739 19672 18788 19700
rect 18739 19669 18751 19672
rect 18693 19663 18751 19669
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 19061 19703 19119 19709
rect 19061 19669 19073 19703
rect 19107 19700 19119 19703
rect 19150 19700 19156 19712
rect 19107 19672 19156 19700
rect 19107 19669 19119 19672
rect 19061 19663 19119 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1670 19496 1676 19508
rect 1631 19468 1676 19496
rect 1670 19456 1676 19468
rect 1728 19456 1734 19508
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 2409 19499 2467 19505
rect 2409 19496 2421 19499
rect 2280 19468 2421 19496
rect 2280 19456 2286 19468
rect 2409 19465 2421 19468
rect 2455 19465 2467 19499
rect 4617 19499 4675 19505
rect 4617 19496 4629 19499
rect 2409 19459 2467 19465
rect 3068 19468 4629 19496
rect 1762 19320 1768 19372
rect 1820 19360 1826 19372
rect 2041 19363 2099 19369
rect 2041 19360 2053 19363
rect 1820 19332 2053 19360
rect 1820 19320 1826 19332
rect 2041 19329 2053 19332
rect 2087 19329 2099 19363
rect 2866 19360 2872 19372
rect 2827 19332 2872 19360
rect 2041 19323 2099 19329
rect 2866 19320 2872 19332
rect 2924 19320 2930 19372
rect 3068 19369 3096 19468
rect 4617 19465 4629 19468
rect 4663 19465 4675 19499
rect 4890 19496 4896 19508
rect 4617 19459 4675 19465
rect 4724 19468 4896 19496
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 4632 19360 4660 19459
rect 4724 19440 4752 19468
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 6089 19499 6147 19505
rect 6089 19465 6101 19499
rect 6135 19496 6147 19499
rect 6270 19496 6276 19508
rect 6135 19468 6276 19496
rect 6135 19465 6147 19468
rect 6089 19459 6147 19465
rect 6270 19456 6276 19468
rect 6328 19456 6334 19508
rect 8110 19496 8116 19508
rect 7024 19468 8116 19496
rect 4706 19388 4712 19440
rect 4764 19388 4770 19440
rect 4632 19332 4844 19360
rect 3053 19323 3111 19329
rect 1489 19295 1547 19301
rect 1489 19261 1501 19295
rect 1535 19261 1547 19295
rect 1489 19255 1547 19261
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 2498 19292 2504 19304
rect 1903 19264 2504 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 1504 19224 1532 19255
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 2774 19252 2780 19304
rect 2832 19292 2838 19304
rect 3237 19295 3295 19301
rect 2832 19264 2877 19292
rect 2832 19252 2838 19264
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 4706 19292 4712 19304
rect 3283 19264 4712 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 1504 19196 2084 19224
rect 2056 19156 2084 19196
rect 2590 19184 2596 19236
rect 2648 19224 2654 19236
rect 3252 19224 3280 19255
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 4816 19292 4844 19332
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 7024 19369 7052 19468
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 11054 19496 11060 19508
rect 10796 19468 11060 19496
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6972 19332 7021 19360
rect 6972 19320 6978 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 8662 19360 8668 19372
rect 8623 19332 8668 19360
rect 7009 19323 7067 19329
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 4965 19295 5023 19301
rect 4965 19292 4977 19295
rect 4816 19264 4977 19292
rect 4965 19261 4977 19264
rect 5011 19261 5023 19295
rect 6178 19292 6184 19304
rect 6139 19264 6184 19292
rect 4965 19255 5023 19261
rect 6178 19252 6184 19264
rect 6236 19252 6242 19304
rect 7282 19301 7288 19304
rect 7276 19292 7288 19301
rect 6380 19264 7144 19292
rect 7243 19264 7288 19292
rect 2648 19196 3280 19224
rect 3504 19227 3562 19233
rect 2648 19184 2654 19196
rect 3504 19193 3516 19227
rect 3550 19224 3562 19227
rect 4798 19224 4804 19236
rect 3550 19196 4804 19224
rect 3550 19193 3562 19196
rect 3504 19187 3562 19193
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 5074 19184 5080 19236
rect 5132 19224 5138 19236
rect 6380 19224 6408 19264
rect 5132 19196 6408 19224
rect 6457 19227 6515 19233
rect 5132 19184 5138 19196
rect 6457 19193 6469 19227
rect 6503 19193 6515 19227
rect 7116 19224 7144 19264
rect 7276 19255 7288 19264
rect 7282 19252 7288 19255
rect 7340 19252 7346 19304
rect 8478 19292 8484 19304
rect 8439 19264 8484 19292
rect 8478 19252 8484 19264
rect 8536 19252 8542 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 9392 19295 9450 19301
rect 9392 19261 9404 19295
rect 9438 19292 9450 19295
rect 10318 19292 10324 19304
rect 9438 19264 10324 19292
rect 9438 19261 9450 19264
rect 9392 19255 9450 19261
rect 9030 19224 9036 19236
rect 7116 19196 9036 19224
rect 6457 19187 6515 19193
rect 6472 19156 6500 19187
rect 9030 19184 9036 19196
rect 9088 19184 9094 19236
rect 9140 19224 9168 19255
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 10796 19301 10824 19468
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 12158 19496 12164 19508
rect 12119 19468 12164 19496
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 14645 19499 14703 19505
rect 14645 19465 14657 19499
rect 14691 19496 14703 19499
rect 15378 19496 15384 19508
rect 14691 19468 15384 19496
rect 14691 19465 14703 19468
rect 14645 19459 14703 19465
rect 15378 19456 15384 19468
rect 15436 19456 15442 19508
rect 14277 19431 14335 19437
rect 14277 19428 14289 19431
rect 14200 19400 14289 19428
rect 12618 19360 12624 19372
rect 12579 19332 12624 19360
rect 12618 19320 12624 19332
rect 12676 19320 12682 19372
rect 10781 19295 10839 19301
rect 10781 19292 10793 19295
rect 10691 19264 10793 19292
rect 10781 19261 10793 19264
rect 10827 19261 10839 19295
rect 10781 19255 10839 19261
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12710 19292 12716 19304
rect 12483 19264 12716 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 10796 19224 10824 19255
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 12986 19292 12992 19304
rect 12947 19264 12992 19292
rect 12986 19252 12992 19264
rect 13044 19252 13050 19304
rect 13265 19295 13323 19301
rect 13265 19261 13277 19295
rect 13311 19292 13323 19295
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 13311 19264 13553 19292
rect 13311 19261 13323 19264
rect 13265 19255 13323 19261
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 13909 19295 13967 19301
rect 13909 19261 13921 19295
rect 13955 19292 13967 19295
rect 14200 19292 14228 19400
rect 14277 19397 14289 19400
rect 14323 19397 14335 19431
rect 14277 19391 14335 19397
rect 13955 19264 14228 19292
rect 13955 19261 13967 19264
rect 13909 19255 13967 19261
rect 9140 19196 10824 19224
rect 11048 19227 11106 19233
rect 11048 19193 11060 19227
rect 11094 19224 11106 19227
rect 11422 19224 11428 19236
rect 11094 19196 11428 19224
rect 11094 19193 11106 19196
rect 11048 19187 11106 19193
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 13446 19184 13452 19236
rect 13504 19224 13510 19236
rect 13924 19224 13952 19255
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14332 19264 14473 19292
rect 14332 19252 14338 19264
rect 14461 19261 14473 19264
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14792 19264 14841 19292
rect 14792 19252 14798 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15197 19295 15255 19301
rect 15197 19261 15209 19295
rect 15243 19292 15255 19295
rect 15378 19292 15384 19304
rect 15243 19264 15384 19292
rect 15243 19261 15255 19264
rect 15197 19255 15255 19261
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 15654 19292 15660 19304
rect 15615 19264 15660 19292
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 15930 19252 15936 19304
rect 15988 19292 15994 19304
rect 16025 19295 16083 19301
rect 16025 19292 16037 19295
rect 15988 19264 16037 19292
rect 15988 19252 15994 19264
rect 16025 19261 16037 19264
rect 16071 19261 16083 19295
rect 16025 19255 16083 19261
rect 16577 19295 16635 19301
rect 16577 19261 16589 19295
rect 16623 19292 16635 19295
rect 16850 19292 16856 19304
rect 16623 19264 16856 19292
rect 16623 19261 16635 19264
rect 16577 19255 16635 19261
rect 16850 19252 16856 19264
rect 16908 19252 16914 19304
rect 17494 19292 17500 19304
rect 17455 19264 17500 19292
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18782 19292 18788 19304
rect 18743 19264 18788 19292
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 19150 19292 19156 19304
rect 19111 19264 19156 19292
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19518 19292 19524 19304
rect 19479 19264 19524 19292
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 14366 19224 14372 19236
rect 13504 19196 13952 19224
rect 14108 19196 14372 19224
rect 13504 19184 13510 19196
rect 2056 19128 6500 19156
rect 7374 19116 7380 19168
rect 7432 19156 7438 19168
rect 8389 19159 8447 19165
rect 8389 19156 8401 19159
rect 7432 19128 8401 19156
rect 7432 19116 7438 19128
rect 8389 19125 8401 19128
rect 8435 19125 8447 19159
rect 8389 19119 8447 19125
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 10505 19159 10563 19165
rect 10505 19156 10517 19159
rect 9364 19128 10517 19156
rect 9364 19116 9370 19128
rect 10505 19125 10517 19128
rect 10551 19125 10563 19159
rect 10505 19119 10563 19125
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 14108 19165 14136 19196
rect 14366 19184 14372 19196
rect 14424 19184 14430 19236
rect 14918 19184 14924 19236
rect 14976 19224 14982 19236
rect 16298 19224 16304 19236
rect 14976 19196 15056 19224
rect 14976 19184 14982 19196
rect 15028 19165 15056 19196
rect 15856 19196 16304 19224
rect 13725 19159 13783 19165
rect 13725 19156 13737 19159
rect 13596 19128 13737 19156
rect 13596 19116 13602 19128
rect 13725 19125 13737 19128
rect 13771 19125 13783 19159
rect 13725 19119 13783 19125
rect 14093 19159 14151 19165
rect 14093 19125 14105 19159
rect 14139 19125 14151 19159
rect 14093 19119 14151 19125
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19125 15071 19159
rect 15013 19119 15071 19125
rect 15381 19159 15439 19165
rect 15381 19125 15393 19159
rect 15427 19156 15439 19159
rect 15746 19156 15752 19168
rect 15427 19128 15752 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 15856 19165 15884 19196
rect 16298 19184 16304 19196
rect 16356 19184 16362 19236
rect 17218 19224 17224 19236
rect 17179 19196 17224 19224
rect 17218 19184 17224 19196
rect 17276 19184 17282 19236
rect 19978 19224 19984 19236
rect 19352 19196 19984 19224
rect 15841 19159 15899 19165
rect 15841 19125 15853 19159
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 16209 19159 16267 19165
rect 16209 19125 16221 19159
rect 16255 19156 16267 19159
rect 16758 19156 16764 19168
rect 16255 19128 16764 19156
rect 16255 19125 16267 19128
rect 16209 19119 16267 19125
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 17678 19156 17684 19168
rect 17639 19128 17684 19156
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 18196 19128 18245 19156
rect 18196 19116 18202 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18598 19156 18604 19168
rect 18559 19128 18604 19156
rect 18233 19119 18291 19125
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 18969 19159 19027 19165
rect 18969 19125 18981 19159
rect 19015 19156 19027 19159
rect 19058 19156 19064 19168
rect 19015 19128 19064 19156
rect 19015 19125 19027 19128
rect 18969 19119 19027 19125
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 19352 19165 19380 19196
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 19337 19159 19395 19165
rect 19337 19125 19349 19159
rect 19383 19125 19395 19159
rect 19337 19119 19395 19125
rect 19705 19159 19763 19165
rect 19705 19125 19717 19159
rect 19751 19156 19763 19159
rect 20438 19156 20444 19168
rect 19751 19128 20444 19156
rect 19751 19125 19763 19128
rect 19705 19119 19763 19125
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 4614 18952 4620 18964
rect 2056 18924 4620 18952
rect 1118 18844 1124 18896
rect 1176 18884 1182 18896
rect 2056 18884 2084 18924
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 4798 18912 4804 18964
rect 4856 18952 4862 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 4856 18924 8309 18952
rect 4856 18912 4862 18924
rect 8297 18921 8309 18924
rect 8343 18921 8355 18955
rect 8297 18915 8355 18921
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 8757 18955 8815 18961
rect 8757 18952 8769 18955
rect 8536 18924 8769 18952
rect 8536 18912 8542 18924
rect 8757 18921 8769 18924
rect 8803 18921 8815 18955
rect 8757 18915 8815 18921
rect 9217 18955 9275 18961
rect 9217 18921 9229 18955
rect 9263 18952 9275 18955
rect 9674 18952 9680 18964
rect 9263 18924 9680 18952
rect 9263 18921 9275 18924
rect 9217 18915 9275 18921
rect 9674 18912 9680 18924
rect 9732 18912 9738 18964
rect 12250 18952 12256 18964
rect 12163 18924 12256 18952
rect 12250 18912 12256 18924
rect 12308 18952 12314 18964
rect 12802 18952 12808 18964
rect 12308 18924 12808 18952
rect 12308 18912 12314 18924
rect 12802 18912 12808 18924
rect 12860 18912 12866 18964
rect 15930 18952 15936 18964
rect 14384 18924 15936 18952
rect 1176 18856 2084 18884
rect 1176 18844 1182 18856
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 2501 18887 2559 18893
rect 2501 18884 2513 18887
rect 2188 18856 2513 18884
rect 2188 18844 2194 18856
rect 2501 18853 2513 18856
rect 2547 18853 2559 18887
rect 2501 18847 2559 18853
rect 5252 18887 5310 18893
rect 5252 18853 5264 18887
rect 5298 18884 5310 18887
rect 5718 18884 5724 18896
rect 5298 18856 5724 18884
rect 5298 18853 5310 18856
rect 5252 18847 5310 18853
rect 5718 18844 5724 18856
rect 5776 18884 5782 18896
rect 6362 18884 6368 18896
rect 5776 18856 6368 18884
rect 5776 18844 5782 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 7184 18887 7242 18893
rect 7184 18853 7196 18887
rect 7230 18884 7242 18887
rect 7374 18884 7380 18896
rect 7230 18856 7380 18884
rect 7230 18853 7242 18856
rect 7184 18847 7242 18853
rect 7374 18844 7380 18856
rect 7432 18844 7438 18896
rect 12161 18887 12219 18893
rect 8864 18856 11836 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2235 18819 2293 18825
rect 2235 18785 2247 18819
rect 2281 18785 2293 18819
rect 2235 18779 2293 18785
rect 3605 18819 3663 18825
rect 3605 18785 3617 18819
rect 3651 18816 3663 18819
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3651 18788 4445 18816
rect 3651 18785 3663 18788
rect 3605 18779 3663 18785
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 2240 18680 2268 18779
rect 4706 18776 4712 18828
rect 4764 18816 4770 18828
rect 4985 18819 5043 18825
rect 4985 18816 4997 18819
rect 4764 18788 4997 18816
rect 4764 18776 4770 18788
rect 4985 18785 4997 18788
rect 5031 18816 5043 18819
rect 6914 18816 6920 18828
rect 5031 18788 6920 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 6914 18776 6920 18788
rect 6972 18776 6978 18828
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 8864 18816 8892 18856
rect 8812 18788 8892 18816
rect 9125 18819 9183 18825
rect 8812 18776 8818 18788
rect 9125 18785 9137 18819
rect 9171 18816 9183 18819
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9171 18788 9689 18816
rect 9171 18785 9183 18788
rect 9125 18779 9183 18785
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 10229 18819 10287 18825
rect 10229 18785 10241 18819
rect 10275 18816 10287 18819
rect 10870 18816 10876 18828
rect 10275 18788 10876 18816
rect 10275 18785 10287 18788
rect 10229 18779 10287 18785
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18816 11299 18819
rect 11698 18816 11704 18828
rect 11287 18788 11704 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11808 18816 11836 18856
rect 12161 18853 12173 18887
rect 12207 18884 12219 18887
rect 12434 18884 12440 18896
rect 12207 18856 12440 18884
rect 12207 18853 12219 18856
rect 12161 18847 12219 18853
rect 12434 18844 12440 18856
rect 12492 18884 12498 18896
rect 14384 18893 14412 18924
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 16500 18924 18521 18952
rect 12621 18887 12679 18893
rect 12621 18884 12633 18887
rect 12492 18856 12633 18884
rect 12492 18844 12498 18856
rect 12621 18853 12633 18856
rect 12667 18853 12679 18887
rect 12621 18847 12679 18853
rect 14369 18887 14427 18893
rect 14369 18853 14381 18887
rect 14415 18853 14427 18887
rect 14369 18847 14427 18853
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 14921 18887 14979 18893
rect 14921 18884 14933 18887
rect 14792 18856 14933 18884
rect 14792 18844 14798 18856
rect 14921 18853 14933 18856
rect 14967 18853 14979 18887
rect 14921 18847 14979 18853
rect 11808 18788 13860 18816
rect 4246 18708 4252 18760
rect 4304 18748 4310 18760
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4304 18720 4537 18748
rect 4304 18708 4310 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18717 4675 18751
rect 9306 18748 9312 18760
rect 9267 18720 9312 18748
rect 4617 18711 4675 18717
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 2240 18652 4077 18680
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4065 18643 4123 18649
rect 658 18572 664 18624
rect 716 18612 722 18624
rect 2682 18612 2688 18624
rect 716 18584 2688 18612
rect 716 18572 722 18584
rect 2682 18572 2688 18584
rect 2740 18572 2746 18624
rect 3970 18572 3976 18624
rect 4028 18612 4034 18624
rect 4632 18612 4660 18711
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 10410 18748 10416 18760
rect 10371 18720 10416 18748
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10686 18708 10692 18760
rect 10744 18748 10750 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 10744 18720 11345 18748
rect 10744 18708 10750 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 11422 18708 11428 18760
rect 11480 18748 11486 18760
rect 12342 18748 12348 18760
rect 11480 18720 12348 18748
rect 11480 18708 11486 18720
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 13832 18748 13860 18788
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 13964 18788 14105 18816
rect 13964 18776 13970 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 14645 18819 14703 18825
rect 14645 18785 14657 18819
rect 14691 18816 14703 18819
rect 15194 18816 15200 18828
rect 14691 18788 15200 18816
rect 14691 18785 14703 18788
rect 14645 18779 14703 18785
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 16500 18748 16528 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 16945 18887 17003 18893
rect 16945 18853 16957 18887
rect 16991 18884 17003 18887
rect 18414 18884 18420 18896
rect 16991 18856 18420 18884
rect 16991 18853 17003 18856
rect 16945 18847 17003 18853
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 16669 18819 16727 18825
rect 16669 18785 16681 18819
rect 16715 18785 16727 18819
rect 16669 18779 16727 18785
rect 13832 18720 16528 18748
rect 5994 18640 6000 18692
rect 6052 18680 6058 18692
rect 6052 18652 6960 18680
rect 6052 18640 6058 18652
rect 4028 18584 4660 18612
rect 4028 18572 4034 18584
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 6365 18615 6423 18621
rect 6365 18612 6377 18615
rect 4948 18584 6377 18612
rect 4948 18572 4954 18584
rect 6365 18581 6377 18584
rect 6411 18581 6423 18615
rect 6932 18612 6960 18652
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 16684 18680 16712 18779
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 18524 18816 18552 18915
rect 18969 18887 19027 18893
rect 18969 18853 18981 18887
rect 19015 18884 19027 18887
rect 19518 18884 19524 18896
rect 19015 18856 19524 18884
rect 19015 18853 19027 18856
rect 18969 18847 19027 18853
rect 19518 18844 19524 18856
rect 19576 18844 19582 18896
rect 18693 18819 18751 18825
rect 18693 18816 18705 18819
rect 16908 18788 17632 18816
rect 18524 18788 18705 18816
rect 16908 18776 16914 18788
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17494 18748 17500 18760
rect 17451 18720 17500 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17604 18757 17632 18788
rect 18693 18785 18705 18788
rect 18739 18785 18751 18819
rect 18693 18779 18751 18785
rect 17589 18751 17647 18757
rect 17589 18717 17601 18751
rect 17635 18748 17647 18751
rect 22278 18748 22284 18760
rect 17635 18720 22284 18748
rect 17635 18717 17647 18720
rect 17589 18711 17647 18717
rect 22278 18708 22284 18720
rect 22336 18708 22342 18760
rect 12492 18652 16712 18680
rect 12492 18640 12498 18652
rect 8938 18612 8944 18624
rect 6932 18584 8944 18612
rect 6365 18575 6423 18581
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 10873 18615 10931 18621
rect 10873 18581 10885 18615
rect 10919 18612 10931 18615
rect 11238 18612 11244 18624
rect 10919 18584 11244 18612
rect 10919 18581 10931 18584
rect 10873 18575 10931 18581
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 11790 18612 11796 18624
rect 11751 18584 11796 18612
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 12897 18615 12955 18621
rect 12897 18612 12909 18615
rect 12860 18584 12909 18612
rect 12860 18572 12866 18584
rect 12897 18581 12909 18584
rect 12943 18612 12955 18615
rect 14090 18612 14096 18624
rect 12943 18584 14096 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 14090 18572 14096 18584
rect 14148 18572 14154 18624
rect 15378 18612 15384 18624
rect 15339 18584 15384 18612
rect 15378 18572 15384 18584
rect 15436 18572 15442 18624
rect 15565 18615 15623 18621
rect 15565 18581 15577 18615
rect 15611 18612 15623 18615
rect 15654 18612 15660 18624
rect 15611 18584 15660 18612
rect 15611 18581 15623 18584
rect 15565 18575 15623 18581
rect 15654 18572 15660 18584
rect 15712 18612 15718 18624
rect 16298 18612 16304 18624
rect 15712 18584 16304 18612
rect 15712 18572 15718 18584
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 17957 18615 18015 18621
rect 17957 18581 17969 18615
rect 18003 18612 18015 18615
rect 18046 18612 18052 18624
rect 18003 18584 18052 18612
rect 18003 18581 18015 18584
rect 17957 18575 18015 18581
rect 18046 18572 18052 18584
rect 18104 18572 18110 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1578 18368 1584 18420
rect 1636 18408 1642 18420
rect 2317 18411 2375 18417
rect 2317 18408 2329 18411
rect 1636 18380 2329 18408
rect 1636 18368 1642 18380
rect 2317 18377 2329 18380
rect 2363 18377 2375 18411
rect 2317 18371 2375 18377
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 2556 18380 3547 18408
rect 2556 18368 2562 18380
rect 1946 18340 1952 18352
rect 1907 18312 1952 18340
rect 1946 18300 1952 18312
rect 2004 18300 2010 18352
rect 3519 18340 3547 18380
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 4246 18408 4252 18420
rect 4028 18380 4073 18408
rect 4207 18380 4252 18408
rect 4028 18368 4034 18380
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 4347 18380 4752 18408
rect 4347 18340 4375 18380
rect 3519 18312 4375 18340
rect 4724 18340 4752 18380
rect 4798 18368 4804 18420
rect 4856 18408 4862 18420
rect 10134 18408 10140 18420
rect 4856 18380 10140 18408
rect 4856 18368 4862 18380
rect 10134 18368 10140 18380
rect 10192 18368 10198 18420
rect 10870 18408 10876 18420
rect 10831 18380 10876 18408
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 10980 18380 12296 18408
rect 5077 18343 5135 18349
rect 5077 18340 5089 18343
rect 4724 18312 5089 18340
rect 5077 18309 5089 18312
rect 5123 18309 5135 18343
rect 5077 18303 5135 18309
rect 7742 18300 7748 18352
rect 7800 18340 7806 18352
rect 10980 18340 11008 18380
rect 12158 18340 12164 18352
rect 7800 18312 11008 18340
rect 11532 18312 12164 18340
rect 7800 18300 7806 18312
rect 2590 18272 2596 18284
rect 2551 18244 2596 18272
rect 2590 18232 2596 18244
rect 2648 18232 2654 18284
rect 4890 18272 4896 18284
rect 3804 18244 4896 18272
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 2860 18207 2918 18213
rect 2860 18173 2872 18207
rect 2906 18204 2918 18207
rect 3804 18204 3832 18244
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 5534 18272 5540 18284
rect 5495 18244 5540 18272
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5718 18272 5724 18284
rect 5679 18244 5724 18272
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 9950 18272 9956 18284
rect 9539 18244 9956 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 11532 18281 11560 18312
rect 12158 18300 12164 18312
rect 12216 18300 12222 18352
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18241 11575 18275
rect 11698 18272 11704 18284
rect 11659 18244 11704 18272
rect 11517 18235 11575 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 12268 18272 12296 18380
rect 12342 18368 12348 18420
rect 12400 18408 12406 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 12400 18380 13829 18408
rect 12400 18368 12406 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 14090 18368 14096 18420
rect 14148 18408 14154 18420
rect 17770 18408 17776 18420
rect 14148 18380 17776 18408
rect 14148 18368 14154 18380
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 12434 18300 12440 18352
rect 12492 18300 12498 18352
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 19150 18340 19156 18352
rect 14516 18312 19156 18340
rect 14516 18300 14522 18312
rect 19150 18300 19156 18312
rect 19208 18300 19214 18352
rect 12452 18272 12480 18300
rect 12268 18244 12480 18272
rect 2906 18176 3832 18204
rect 2906 18173 2918 18176
rect 2860 18167 2918 18173
rect 2148 18136 2176 18167
rect 5074 18164 5080 18216
rect 5132 18204 5138 18216
rect 10686 18204 10692 18216
rect 5132 18176 10692 18204
rect 5132 18164 5138 18176
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 11238 18204 11244 18216
rect 11199 18176 11244 18204
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 11333 18207 11391 18213
rect 11333 18173 11345 18207
rect 11379 18204 11391 18207
rect 11790 18204 11796 18216
rect 11379 18176 11796 18204
rect 11379 18173 11391 18176
rect 11333 18167 11391 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 12434 18164 12440 18216
rect 12492 18213 12498 18216
rect 12492 18204 12502 18213
rect 12492 18176 12537 18204
rect 12492 18167 12502 18176
rect 12492 18164 12498 18167
rect 2774 18136 2780 18148
rect 2148 18108 2780 18136
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 4709 18139 4767 18145
rect 4709 18105 4721 18139
rect 4755 18136 4767 18139
rect 5258 18136 5264 18148
rect 4755 18108 5264 18136
rect 4755 18105 4767 18108
rect 4709 18099 4767 18105
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 5445 18139 5503 18145
rect 5445 18105 5457 18139
rect 5491 18136 5503 18139
rect 5905 18139 5963 18145
rect 5905 18136 5917 18139
rect 5491 18108 5917 18136
rect 5491 18105 5503 18108
rect 5445 18099 5503 18105
rect 5905 18105 5917 18108
rect 5951 18105 5963 18139
rect 5905 18099 5963 18105
rect 6270 18096 6276 18148
rect 6328 18136 6334 18148
rect 10778 18136 10784 18148
rect 6328 18108 10784 18136
rect 6328 18096 6334 18108
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 12682 18139 12740 18145
rect 12682 18136 12694 18139
rect 12584 18108 12694 18136
rect 12584 18096 12590 18108
rect 12682 18105 12694 18108
rect 12728 18105 12740 18139
rect 12682 18099 12740 18105
rect 1394 18068 1400 18080
rect 1355 18040 1400 18068
rect 1394 18028 1400 18040
rect 1452 18028 1458 18080
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18068 4215 18071
rect 4430 18068 4436 18080
rect 4203 18040 4436 18068
rect 4203 18037 4215 18040
rect 4157 18031 4215 18037
rect 4430 18028 4436 18040
rect 4488 18068 4494 18080
rect 4617 18071 4675 18077
rect 4617 18068 4629 18071
rect 4488 18040 4629 18068
rect 4488 18028 4494 18040
rect 4617 18037 4629 18040
rect 4663 18068 4675 18071
rect 5350 18068 5356 18080
rect 4663 18040 5356 18068
rect 4663 18037 4675 18040
rect 4617 18031 4675 18037
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 8846 18068 8852 18080
rect 8807 18040 8852 18068
rect 8846 18028 8852 18040
rect 8904 18028 8910 18080
rect 9214 18068 9220 18080
rect 9175 18040 9220 18068
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 9309 18071 9367 18077
rect 9309 18037 9321 18071
rect 9355 18068 9367 18071
rect 9674 18068 9680 18080
rect 9355 18040 9680 18068
rect 9355 18037 9367 18040
rect 9309 18031 9367 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4396 17836 4537 17864
rect 4396 17824 4402 17836
rect 4525 17833 4537 17836
rect 4571 17864 4583 17867
rect 4893 17867 4951 17873
rect 4893 17864 4905 17867
rect 4571 17836 4905 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4893 17833 4905 17836
rect 4939 17833 4951 17867
rect 4893 17827 4951 17833
rect 5169 17867 5227 17873
rect 5169 17833 5181 17867
rect 5215 17864 5227 17867
rect 5258 17864 5264 17876
rect 5215 17836 5264 17864
rect 5215 17833 5227 17836
rect 5169 17827 5227 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5350 17824 5356 17876
rect 5408 17864 5414 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 5408 17836 8493 17864
rect 5408 17824 5414 17836
rect 8481 17833 8493 17836
rect 8527 17864 8539 17867
rect 8573 17867 8631 17873
rect 8573 17864 8585 17867
rect 8527 17836 8585 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 8573 17833 8585 17836
rect 8619 17833 8631 17867
rect 8573 17827 8631 17833
rect 8757 17867 8815 17873
rect 8757 17833 8769 17867
rect 8803 17864 8815 17867
rect 9214 17864 9220 17876
rect 8803 17836 9220 17864
rect 8803 17833 8815 17836
rect 8757 17827 8815 17833
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 11057 17867 11115 17873
rect 11057 17833 11069 17867
rect 11103 17833 11115 17867
rect 11057 17827 11115 17833
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 13998 17864 14004 17876
rect 13771 17836 14004 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2225 17799 2283 17805
rect 2225 17796 2237 17799
rect 1820 17768 2237 17796
rect 1820 17756 1826 17768
rect 2225 17765 2237 17768
rect 2271 17765 2283 17799
rect 2225 17759 2283 17765
rect 2774 17756 2780 17808
rect 2832 17796 2838 17808
rect 8846 17796 8852 17808
rect 2832 17768 2877 17796
rect 2976 17768 8852 17796
rect 2832 17756 2838 17768
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 1854 17728 1860 17740
rect 1627 17700 1860 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17697 2007 17731
rect 1949 17691 2007 17697
rect 1964 17660 1992 17691
rect 2498 17688 2504 17740
rect 2556 17728 2562 17740
rect 2556 17700 2601 17728
rect 2556 17688 2562 17700
rect 2976 17660 3004 17768
rect 8846 17756 8852 17768
rect 8904 17756 8910 17808
rect 10686 17796 10692 17808
rect 9324 17768 10692 17796
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 1964 17632 3004 17660
rect 4417 17697 4445 17728
rect 4479 17697 4491 17731
rect 4417 17691 4491 17697
rect 1765 17595 1823 17601
rect 1765 17561 1777 17595
rect 1811 17592 1823 17595
rect 2958 17592 2964 17604
rect 1811 17564 2964 17592
rect 1811 17561 1823 17564
rect 1765 17555 1823 17561
rect 2958 17552 2964 17564
rect 3016 17552 3022 17604
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 4065 17595 4123 17601
rect 4065 17592 4077 17595
rect 3108 17564 4077 17592
rect 3108 17552 3114 17564
rect 4065 17561 4077 17564
rect 4111 17561 4123 17595
rect 4065 17555 4123 17561
rect 4417 17592 4445 17691
rect 6454 17688 6460 17740
rect 6512 17728 6518 17740
rect 6917 17731 6975 17737
rect 6917 17728 6929 17731
rect 6512 17700 6929 17728
rect 6512 17688 6518 17700
rect 6917 17697 6929 17700
rect 6963 17697 6975 17731
rect 9122 17728 9128 17740
rect 9083 17700 9128 17728
rect 6917 17691 6975 17697
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 4798 17660 4804 17672
rect 4755 17632 4804 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4798 17620 4804 17632
rect 4856 17620 4862 17672
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17660 6423 17663
rect 6546 17660 6552 17672
rect 6411 17632 6552 17660
rect 6411 17629 6423 17632
rect 6365 17623 6423 17629
rect 6546 17620 6552 17632
rect 6604 17660 6610 17672
rect 7009 17663 7067 17669
rect 7009 17660 7021 17663
rect 6604 17632 7021 17660
rect 6604 17620 6610 17632
rect 7009 17629 7021 17632
rect 7055 17629 7067 17663
rect 7009 17623 7067 17629
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17660 7251 17663
rect 7374 17660 7380 17672
rect 7239 17632 7380 17660
rect 7239 17629 7251 17632
rect 7193 17623 7251 17629
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 8481 17663 8539 17669
rect 8481 17629 8493 17663
rect 8527 17660 8539 17663
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 8527 17632 9229 17660
rect 8527 17629 8539 17632
rect 8481 17623 8539 17629
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9324 17592 9352 17768
rect 10686 17756 10692 17768
rect 10744 17756 10750 17808
rect 11072 17796 11100 17827
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 11394 17799 11452 17805
rect 11394 17796 11406 17799
rect 11072 17768 11406 17796
rect 11394 17765 11406 17768
rect 11440 17796 11452 17799
rect 12066 17796 12072 17808
rect 11440 17768 12072 17796
rect 11440 17765 11452 17768
rect 11394 17759 11452 17765
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 9766 17728 9772 17740
rect 9416 17700 9772 17728
rect 9416 17669 9444 17700
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 9950 17737 9956 17740
rect 9944 17728 9956 17737
rect 9911 17700 9956 17728
rect 9944 17691 9956 17700
rect 9950 17688 9956 17691
rect 10008 17688 10014 17740
rect 11054 17688 11060 17740
rect 11112 17728 11118 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 11112 17700 11161 17728
rect 11112 17688 11118 17700
rect 11149 17697 11161 17700
rect 11195 17728 11207 17731
rect 11238 17728 11244 17740
rect 11195 17700 11244 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 4417 17564 9352 17592
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3200 17496 3801 17524
rect 3200 17484 3206 17496
rect 3789 17493 3801 17496
rect 3835 17524 3847 17527
rect 4417 17524 4445 17564
rect 3835 17496 4445 17524
rect 6549 17527 6607 17533
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 6549 17493 6561 17527
rect 6595 17524 6607 17527
rect 7098 17524 7104 17536
rect 6595 17496 7104 17524
rect 6595 17493 6607 17496
rect 6549 17487 6607 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 9692 17524 9720 17623
rect 11164 17524 11192 17691
rect 11238 17688 11244 17700
rect 11296 17728 11302 17740
rect 12434 17728 12440 17740
rect 11296 17700 12440 17728
rect 11296 17688 11302 17700
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 13412 17700 13553 17728
rect 13412 17688 13418 17700
rect 13541 17697 13553 17700
rect 13587 17697 13599 17731
rect 13541 17691 13599 17697
rect 12526 17524 12532 17536
rect 9640 17496 11192 17524
rect 12487 17496 12532 17524
rect 9640 17484 9646 17496
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1670 17280 1676 17332
rect 1728 17320 1734 17332
rect 1765 17323 1823 17329
rect 1765 17320 1777 17323
rect 1728 17292 1777 17320
rect 1728 17280 1734 17292
rect 1765 17289 1777 17292
rect 1811 17289 1823 17323
rect 4062 17320 4068 17332
rect 1765 17283 1823 17289
rect 3436 17292 4068 17320
rect 2133 17187 2191 17193
rect 2133 17184 2145 17187
rect 1596 17156 2145 17184
rect 1596 17125 1624 17156
rect 2133 17153 2145 17156
rect 2179 17153 2191 17187
rect 3050 17184 3056 17196
rect 2133 17147 2191 17153
rect 2608 17156 2912 17184
rect 3011 17156 3056 17184
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17085 1639 17119
rect 1581 17079 1639 17085
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 2608 17116 2636 17156
rect 1995 17088 2636 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2884 17048 2912 17156
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 3234 17184 3240 17196
rect 3195 17156 3240 17184
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 3436 17193 3464 17292
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4798 17320 4804 17332
rect 4759 17292 4804 17320
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 4890 17280 4896 17332
rect 4948 17320 4954 17332
rect 6273 17323 6331 17329
rect 6273 17320 6285 17323
rect 4948 17292 6285 17320
rect 4948 17280 4954 17292
rect 6273 17289 6285 17292
rect 6319 17320 6331 17323
rect 9677 17323 9735 17329
rect 6319 17292 9352 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 4816 17184 4844 17280
rect 6454 17184 6460 17196
rect 4816 17156 5028 17184
rect 6415 17156 6460 17184
rect 3421 17147 3479 17153
rect 3688 17119 3746 17125
rect 3688 17085 3700 17119
rect 3734 17116 3746 17119
rect 3970 17116 3976 17128
rect 3734 17088 3976 17116
rect 3734 17085 3746 17088
rect 3688 17079 3746 17085
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4798 17116 4804 17128
rect 4120 17088 4804 17116
rect 4120 17076 4126 17088
rect 4798 17076 4804 17088
rect 4856 17116 4862 17128
rect 4893 17119 4951 17125
rect 4893 17116 4905 17119
rect 4856 17088 4905 17116
rect 4856 17076 4862 17088
rect 4893 17085 4905 17088
rect 4939 17085 4951 17119
rect 5000 17116 5028 17156
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 6822 17184 6828 17196
rect 6783 17156 6828 17184
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 8110 17144 8116 17196
rect 8168 17184 8174 17196
rect 8297 17187 8355 17193
rect 8297 17184 8309 17187
rect 8168 17156 8309 17184
rect 8168 17144 8174 17156
rect 8297 17153 8309 17156
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 5149 17119 5207 17125
rect 5149 17116 5161 17119
rect 5000 17088 5161 17116
rect 4893 17079 4951 17085
rect 5149 17085 5161 17088
rect 5195 17085 5207 17119
rect 5149 17079 5207 17085
rect 6730 17048 6736 17060
rect 2884 17020 6736 17048
rect 6730 17008 6736 17020
rect 6788 17008 6794 17060
rect 6840 17048 6868 17144
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7092 17119 7150 17125
rect 7092 17116 7104 17119
rect 6972 17088 7104 17116
rect 6972 17076 6978 17088
rect 7092 17085 7104 17088
rect 7138 17116 7150 17119
rect 7374 17116 7380 17128
rect 7138 17088 7380 17116
rect 7138 17085 7150 17088
rect 7092 17079 7150 17085
rect 7374 17076 7380 17088
rect 7432 17116 7438 17128
rect 8202 17116 8208 17128
rect 7432 17088 8208 17116
rect 7432 17076 7438 17088
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 7190 17048 7196 17060
rect 6840 17020 7196 17048
rect 7190 17008 7196 17020
rect 7248 17048 7254 17060
rect 8110 17048 8116 17060
rect 7248 17020 8116 17048
rect 7248 17008 7254 17020
rect 8110 17008 8116 17020
rect 8168 17008 8174 17060
rect 8542 17051 8600 17057
rect 8542 17048 8554 17051
rect 8220 17020 8554 17048
rect 2130 16940 2136 16992
rect 2188 16980 2194 16992
rect 2593 16983 2651 16989
rect 2593 16980 2605 16983
rect 2188 16952 2605 16980
rect 2188 16940 2194 16952
rect 2593 16949 2605 16952
rect 2639 16949 2651 16983
rect 2958 16980 2964 16992
rect 2919 16952 2964 16980
rect 2593 16943 2651 16949
rect 2958 16940 2964 16952
rect 3016 16940 3022 16992
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 6638 16980 6644 16992
rect 3476 16952 6644 16980
rect 3476 16940 3482 16952
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 8220 16989 8248 17020
rect 8542 17017 8554 17020
rect 8588 17017 8600 17051
rect 9324 17048 9352 17292
rect 9677 17289 9689 17323
rect 9723 17320 9735 17323
rect 9766 17320 9772 17332
rect 9723 17292 9772 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 11149 17323 11207 17329
rect 11149 17320 11161 17323
rect 10008 17292 11161 17320
rect 10008 17280 10014 17292
rect 11149 17289 11161 17292
rect 11195 17289 11207 17323
rect 11149 17283 11207 17289
rect 9784 17184 9812 17280
rect 12066 17184 12072 17196
rect 9784 17156 9904 17184
rect 12027 17156 12072 17184
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 9640 17088 9781 17116
rect 9640 17076 9646 17088
rect 9769 17085 9781 17088
rect 9815 17085 9827 17119
rect 9876 17116 9904 17156
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 13354 17184 13360 17196
rect 13315 17156 13360 17184
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 10025 17119 10083 17125
rect 10025 17116 10037 17119
rect 9876 17088 10037 17116
rect 9769 17079 9827 17085
rect 10025 17085 10037 17088
rect 10071 17116 10083 17119
rect 10318 17116 10324 17128
rect 10071 17088 10324 17116
rect 10071 17085 10083 17088
rect 10025 17079 10083 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 11885 17119 11943 17125
rect 11885 17085 11897 17119
rect 11931 17116 11943 17119
rect 12529 17119 12587 17125
rect 12529 17116 12541 17119
rect 11931 17088 12541 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 12529 17085 12541 17088
rect 12575 17116 12587 17119
rect 12894 17116 12900 17128
rect 12575 17088 12900 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13081 17119 13139 17125
rect 13081 17085 13093 17119
rect 13127 17116 13139 17119
rect 14182 17116 14188 17128
rect 13127 17088 14188 17116
rect 13127 17085 13139 17088
rect 13081 17079 13139 17085
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 17954 17048 17960 17060
rect 9324 17020 17960 17048
rect 8542 17011 8600 17017
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 8205 16983 8263 16989
rect 8205 16980 8217 16983
rect 7432 16952 8217 16980
rect 7432 16940 7438 16952
rect 8205 16949 8217 16952
rect 8251 16949 8263 16983
rect 8205 16943 8263 16949
rect 11241 16983 11299 16989
rect 11241 16949 11253 16983
rect 11287 16980 11299 16983
rect 11330 16980 11336 16992
rect 11287 16952 11336 16980
rect 11287 16949 11299 16952
rect 11241 16943 11299 16949
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 11514 16980 11520 16992
rect 11475 16952 11520 16980
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 11977 16983 12035 16989
rect 11977 16980 11989 16983
rect 11940 16952 11989 16980
rect 11940 16940 11946 16952
rect 11977 16949 11989 16952
rect 12023 16980 12035 16983
rect 12713 16983 12771 16989
rect 12713 16980 12725 16983
rect 12023 16952 12725 16980
rect 12023 16949 12035 16952
rect 11977 16943 12035 16949
rect 12713 16949 12725 16952
rect 12759 16980 12771 16983
rect 15470 16980 15476 16992
rect 12759 16952 15476 16980
rect 12759 16949 12771 16952
rect 12713 16943 12771 16949
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3605 16779 3663 16785
rect 3605 16776 3617 16779
rect 3016 16748 3617 16776
rect 3016 16736 3022 16748
rect 3605 16745 3617 16748
rect 3651 16745 3663 16779
rect 4890 16776 4896 16788
rect 3605 16739 3663 16745
rect 4448 16748 4896 16776
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 2409 16711 2467 16717
rect 2409 16708 2421 16711
rect 1912 16680 2421 16708
rect 1912 16668 1918 16680
rect 2409 16677 2421 16680
rect 2455 16677 2467 16711
rect 2409 16671 2467 16677
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 3513 16711 3571 16717
rect 3513 16708 3525 16711
rect 3292 16680 3525 16708
rect 3292 16668 3298 16680
rect 3513 16677 3525 16680
rect 3559 16708 3571 16711
rect 4448 16708 4476 16748
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 6549 16779 6607 16785
rect 6549 16745 6561 16779
rect 6595 16776 6607 16779
rect 6914 16776 6920 16788
rect 6595 16748 6920 16776
rect 6595 16745 6607 16748
rect 6549 16739 6607 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7098 16776 7104 16788
rect 7059 16748 7104 16776
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7193 16779 7251 16785
rect 7193 16745 7205 16779
rect 7239 16776 7251 16779
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7239 16748 7665 16776
rect 7239 16745 7251 16748
rect 7193 16739 7251 16745
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 9122 16776 9128 16788
rect 9083 16748 9128 16776
rect 7653 16739 7711 16745
rect 9122 16736 9128 16748
rect 9180 16736 9186 16788
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10045 16779 10103 16785
rect 10045 16745 10057 16779
rect 10091 16776 10103 16779
rect 10594 16776 10600 16788
rect 10091 16748 10600 16776
rect 10091 16745 10103 16748
rect 10045 16739 10103 16745
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 10965 16779 11023 16785
rect 10965 16745 10977 16779
rect 11011 16776 11023 16779
rect 11330 16776 11336 16788
rect 11011 16748 11192 16776
rect 11291 16748 11336 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 3559 16680 4476 16708
rect 4525 16711 4583 16717
rect 3559 16677 3571 16680
rect 3513 16671 3571 16677
rect 4525 16677 4537 16711
rect 4571 16708 4583 16711
rect 6822 16708 6828 16720
rect 4571 16680 6828 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 7282 16668 7288 16720
rect 7340 16708 7346 16720
rect 11164 16708 11192 16748
rect 11330 16736 11336 16748
rect 11388 16736 11394 16788
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 12253 16779 12311 16785
rect 12253 16776 12265 16779
rect 11572 16748 12265 16776
rect 11572 16736 11578 16748
rect 12253 16745 12265 16748
rect 12299 16745 12311 16779
rect 12253 16739 12311 16745
rect 12161 16711 12219 16717
rect 12161 16708 12173 16711
rect 7340 16680 11008 16708
rect 11164 16680 12173 16708
rect 7340 16668 7346 16680
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2130 16640 2136 16652
rect 2091 16612 2136 16640
rect 2130 16600 2136 16612
rect 2188 16600 2194 16652
rect 4246 16600 4252 16652
rect 4304 16640 4310 16652
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4304 16612 4445 16640
rect 4304 16600 4310 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 5258 16640 5264 16652
rect 4433 16603 4491 16609
rect 4724 16612 5264 16640
rect 4724 16581 4752 16612
rect 5258 16600 5264 16612
rect 5316 16640 5322 16652
rect 5425 16643 5483 16649
rect 5425 16640 5437 16643
rect 5316 16612 5437 16640
rect 5316 16600 5322 16612
rect 5425 16609 5437 16612
rect 5471 16609 5483 16643
rect 5425 16603 5483 16609
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16640 8171 16643
rect 8757 16643 8815 16649
rect 8757 16640 8769 16643
rect 8159 16612 8769 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 8757 16609 8769 16612
rect 8803 16640 8815 16643
rect 10042 16640 10048 16652
rect 8803 16612 10048 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16541 4767 16575
rect 4709 16535 4767 16541
rect 4798 16532 4804 16584
rect 4856 16572 4862 16584
rect 5169 16575 5227 16581
rect 5169 16572 5181 16575
rect 4856 16544 5181 16572
rect 4856 16532 4862 16544
rect 5169 16541 5181 16544
rect 5215 16541 5227 16575
rect 7374 16572 7380 16584
rect 7335 16544 7380 16572
rect 5169 16535 5227 16541
rect 4890 16464 4896 16516
rect 4948 16504 4954 16516
rect 5074 16504 5080 16516
rect 4948 16476 5080 16504
rect 4948 16464 4954 16476
rect 5074 16464 5080 16476
rect 5132 16464 5138 16516
rect 3510 16396 3516 16448
rect 3568 16436 3574 16448
rect 4065 16439 4123 16445
rect 4065 16436 4077 16439
rect 3568 16408 4077 16436
rect 3568 16396 3574 16408
rect 4065 16405 4077 16408
rect 4111 16405 4123 16439
rect 5184 16436 5212 16535
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 6730 16504 6736 16516
rect 6691 16476 6736 16504
rect 6730 16464 6736 16476
rect 6788 16464 6794 16516
rect 7190 16436 7196 16448
rect 5184 16408 7196 16436
rect 4065 16399 4123 16405
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 8036 16436 8064 16603
rect 10042 16600 10048 16612
rect 10100 16600 10106 16652
rect 10226 16600 10232 16652
rect 10284 16640 10290 16652
rect 10873 16643 10931 16649
rect 10873 16640 10885 16643
rect 10284 16612 10885 16640
rect 10284 16600 10290 16612
rect 10873 16609 10885 16612
rect 10919 16609 10931 16643
rect 10980 16640 11008 16680
rect 12161 16677 12173 16680
rect 12207 16677 12219 16711
rect 12161 16671 12219 16677
rect 10980 16612 11560 16640
rect 10873 16603 10931 16609
rect 8202 16572 8208 16584
rect 8163 16544 8208 16572
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 10137 16575 10195 16581
rect 10137 16541 10149 16575
rect 10183 16541 10195 16575
rect 10318 16572 10324 16584
rect 10279 16544 10324 16572
rect 10137 16535 10195 16541
rect 10152 16504 10180 16535
rect 10318 16532 10324 16544
rect 10376 16532 10382 16584
rect 10594 16572 10600 16584
rect 10555 16544 10600 16572
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10686 16532 10692 16584
rect 10744 16572 10750 16584
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10744 16544 11437 16572
rect 10744 16532 10750 16544
rect 11425 16541 11437 16544
rect 11471 16541 11483 16575
rect 11425 16535 11483 16541
rect 11146 16504 11152 16516
rect 10152 16476 11152 16504
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 11532 16504 11560 16612
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 12066 16572 12072 16584
rect 11655 16544 12072 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 12526 16572 12532 16584
rect 12391 16544 12532 16572
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 11793 16507 11851 16513
rect 11793 16504 11805 16507
rect 11532 16476 11805 16504
rect 11793 16473 11805 16476
rect 11839 16473 11851 16507
rect 11793 16467 11851 16473
rect 8573 16439 8631 16445
rect 8573 16436 8585 16439
rect 8036 16408 8585 16436
rect 8573 16405 8585 16408
rect 8619 16436 8631 16439
rect 10502 16436 10508 16448
rect 8619 16408 10508 16436
rect 8619 16405 8631 16408
rect 8573 16399 8631 16405
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 10689 16439 10747 16445
rect 10689 16405 10701 16439
rect 10735 16436 10747 16439
rect 10870 16436 10876 16448
rect 10735 16408 10876 16436
rect 10735 16405 10747 16408
rect 10689 16399 10747 16405
rect 10870 16396 10876 16408
rect 10928 16436 10934 16448
rect 11238 16436 11244 16448
rect 10928 16408 11244 16436
rect 10928 16396 10934 16408
rect 11238 16396 11244 16408
rect 11296 16436 11302 16448
rect 12526 16436 12532 16448
rect 11296 16408 12532 16436
rect 11296 16396 11302 16408
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 4062 16232 4068 16244
rect 3804 16204 4068 16232
rect 1394 16056 1400 16108
rect 1452 16096 1458 16108
rect 3804 16105 3832 16204
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 5258 16232 5264 16244
rect 5215 16204 5264 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6822 16192 6828 16244
rect 6880 16232 6886 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 6880 16204 7941 16232
rect 6880 16192 6886 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 8846 16232 8852 16244
rect 7929 16195 7987 16201
rect 8312 16204 8852 16232
rect 6181 16167 6239 16173
rect 6181 16133 6193 16167
rect 6227 16164 6239 16167
rect 7190 16164 7196 16176
rect 6227 16136 7196 16164
rect 6227 16133 6239 16136
rect 6181 16127 6239 16133
rect 7190 16124 7196 16136
rect 7248 16124 7254 16176
rect 2317 16099 2375 16105
rect 2317 16096 2329 16099
rect 1452 16068 2329 16096
rect 1452 16056 1458 16068
rect 2317 16065 2329 16068
rect 2363 16065 2375 16099
rect 2317 16059 2375 16065
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16065 3847 16099
rect 8312 16096 8340 16204
rect 8846 16192 8852 16204
rect 8904 16232 8910 16244
rect 9858 16232 9864 16244
rect 8904 16204 9864 16232
rect 8904 16192 8910 16204
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 11790 16232 11796 16244
rect 10336 16204 11796 16232
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 8312 16068 8401 16096
rect 3789 16059 3847 16065
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16096 8815 16099
rect 10336 16096 10364 16204
rect 11790 16192 11796 16204
rect 11848 16232 11854 16244
rect 11974 16232 11980 16244
rect 11848 16204 11980 16232
rect 11848 16192 11854 16204
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 8803 16068 10364 16096
rect 10873 16099 10931 16105
rect 8803 16065 8815 16068
rect 8757 16059 8815 16065
rect 10873 16065 10885 16099
rect 10919 16096 10931 16099
rect 11422 16096 11428 16108
rect 10919 16068 11428 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 3510 16028 3516 16040
rect 2179 16000 3516 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 1780 15892 1808 15991
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 5718 15988 5724 16040
rect 5776 16028 5782 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 5776 16000 6377 16028
rect 5776 15988 5782 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 2866 15960 2872 15972
rect 2516 15932 2872 15960
rect 2516 15892 2544 15932
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 4056 15963 4114 15969
rect 4056 15929 4068 15963
rect 4102 15960 4114 15963
rect 4614 15960 4620 15972
rect 4102 15932 4620 15960
rect 4102 15929 4114 15932
rect 4056 15923 4114 15929
rect 4614 15920 4620 15932
rect 4672 15960 4678 15972
rect 8496 15960 8524 16059
rect 8662 15960 8668 15972
rect 4672 15932 8668 15960
rect 4672 15920 4678 15932
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 1780 15864 2544 15892
rect 2682 15852 2688 15904
rect 2740 15892 2746 15904
rect 8202 15892 8208 15904
rect 2740 15864 8208 15892
rect 2740 15852 2746 15864
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8297 15895 8355 15901
rect 8297 15861 8309 15895
rect 8343 15892 8355 15895
rect 8772 15892 8800 16059
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16096 11759 16099
rect 12618 16096 12624 16108
rect 11747 16068 12624 16096
rect 11747 16065 11759 16068
rect 11701 16059 11759 16065
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 11238 16028 11244 16040
rect 10735 16000 11244 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 13449 16031 13507 16037
rect 13449 16028 13461 16031
rect 12584 16000 13461 16028
rect 12584 15988 12590 16000
rect 13449 15997 13461 16000
rect 13495 15997 13507 16031
rect 13449 15991 13507 15997
rect 11517 15963 11575 15969
rect 11517 15960 11529 15963
rect 10244 15932 11529 15960
rect 8343 15864 8800 15892
rect 8343 15861 8355 15864
rect 8297 15855 8355 15861
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 10244 15901 10272 15932
rect 11517 15929 11529 15932
rect 11563 15929 11575 15963
rect 11517 15923 11575 15929
rect 13716 15963 13774 15969
rect 13716 15929 13728 15963
rect 13762 15960 13774 15963
rect 14090 15960 14096 15972
rect 13762 15932 14096 15960
rect 13762 15929 13774 15932
rect 13716 15923 13774 15929
rect 14090 15920 14096 15932
rect 14148 15920 14154 15972
rect 8941 15895 8999 15901
rect 8941 15892 8953 15895
rect 8904 15864 8953 15892
rect 8904 15852 8910 15864
rect 8941 15861 8953 15864
rect 8987 15861 8999 15895
rect 8941 15855 8999 15861
rect 10229 15895 10287 15901
rect 10229 15861 10241 15895
rect 10275 15861 10287 15895
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10229 15855 10287 15861
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 11054 15892 11060 15904
rect 11015 15864 11060 15892
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11425 15895 11483 15901
rect 11425 15892 11437 15895
rect 11204 15864 11437 15892
rect 11204 15852 11210 15864
rect 11425 15861 11437 15864
rect 11471 15861 11483 15895
rect 11425 15855 11483 15861
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 14829 15895 14887 15901
rect 14829 15892 14841 15895
rect 14700 15864 14841 15892
rect 14700 15852 14706 15864
rect 14829 15861 14841 15864
rect 14875 15861 14887 15895
rect 14829 15855 14887 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 4065 15691 4123 15697
rect 2832 15660 2877 15688
rect 2832 15648 2838 15660
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4246 15688 4252 15700
rect 4111 15660 4252 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 4525 15691 4583 15697
rect 4525 15688 4537 15691
rect 4396 15660 4537 15688
rect 4396 15648 4402 15660
rect 4525 15657 4537 15660
rect 4571 15657 4583 15691
rect 8662 15688 8668 15700
rect 8623 15660 8668 15688
rect 4525 15651 4583 15657
rect 8662 15648 8668 15660
rect 8720 15648 8726 15700
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9401 15691 9459 15697
rect 9401 15688 9413 15691
rect 9088 15660 9413 15688
rect 9088 15648 9094 15660
rect 9401 15657 9413 15660
rect 9447 15657 9459 15691
rect 9401 15651 9459 15657
rect 9677 15691 9735 15697
rect 9677 15657 9689 15691
rect 9723 15688 9735 15691
rect 10594 15688 10600 15700
rect 9723 15660 10600 15688
rect 9723 15657 9735 15660
rect 9677 15651 9735 15657
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 10962 15688 10968 15700
rect 10827 15660 10968 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 12618 15688 12624 15700
rect 11112 15660 12480 15688
rect 12531 15660 12624 15688
rect 11112 15648 11118 15660
rect 5534 15620 5540 15632
rect 2056 15592 5540 15620
rect 2056 15561 2084 15592
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 7282 15620 7288 15632
rect 5828 15592 7288 15620
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 2314 15512 2320 15564
rect 2372 15552 2378 15564
rect 2593 15555 2651 15561
rect 2593 15552 2605 15555
rect 2372 15524 2605 15552
rect 2372 15512 2378 15524
rect 2593 15521 2605 15524
rect 2639 15521 2651 15555
rect 2593 15515 2651 15521
rect 3418 15512 3424 15564
rect 3476 15552 3482 15564
rect 3881 15555 3939 15561
rect 3881 15552 3893 15555
rect 3476 15524 3893 15552
rect 3476 15512 3482 15524
rect 3881 15521 3893 15524
rect 3927 15552 3939 15555
rect 4154 15552 4160 15564
rect 3927 15524 4160 15552
rect 3927 15521 3939 15524
rect 3881 15515 3939 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 5828 15561 5856 15592
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 7374 15580 7380 15632
rect 7432 15620 7438 15632
rect 7742 15620 7748 15632
rect 7432 15592 7748 15620
rect 7432 15580 7438 15592
rect 7742 15580 7748 15592
rect 7800 15580 7806 15632
rect 8202 15580 8208 15632
rect 8260 15580 8266 15632
rect 9309 15623 9367 15629
rect 9309 15589 9321 15623
rect 9355 15620 9367 15623
rect 9950 15620 9956 15632
rect 9355 15592 9956 15620
rect 9355 15589 9367 15592
rect 9309 15583 9367 15589
rect 9950 15580 9956 15592
rect 10008 15620 10014 15632
rect 10045 15623 10103 15629
rect 10045 15620 10057 15623
rect 10008 15592 10057 15620
rect 10008 15580 10014 15592
rect 10045 15589 10057 15592
rect 10091 15620 10103 15623
rect 10134 15620 10140 15632
rect 10091 15592 10140 15620
rect 10091 15589 10103 15592
rect 10045 15583 10103 15589
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 10873 15623 10931 15629
rect 10873 15620 10885 15623
rect 10744 15592 10885 15620
rect 10744 15580 10750 15592
rect 10873 15589 10885 15592
rect 10919 15589 10931 15623
rect 10873 15583 10931 15589
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4893 15555 4951 15561
rect 4893 15552 4905 15555
rect 4479 15524 4905 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4893 15521 4905 15524
rect 4939 15521 4951 15555
rect 4893 15515 4951 15521
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 6080 15555 6138 15561
rect 6080 15521 6092 15555
rect 6126 15552 6138 15555
rect 6914 15552 6920 15564
rect 6126 15524 6920 15552
rect 6126 15521 6138 15524
rect 6080 15515 6138 15521
rect 6914 15512 6920 15524
rect 6972 15512 6978 15564
rect 7190 15512 7196 15564
rect 7248 15552 7254 15564
rect 7541 15555 7599 15561
rect 7541 15552 7553 15555
rect 7248 15524 7553 15552
rect 7248 15512 7254 15524
rect 7541 15521 7553 15524
rect 7587 15521 7599 15555
rect 8220 15552 8248 15580
rect 8220 15524 10272 15552
rect 7541 15515 7599 15521
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2225 15487 2283 15493
rect 2225 15484 2237 15487
rect 1820 15456 2237 15484
rect 1820 15444 1826 15456
rect 2225 15453 2237 15456
rect 2271 15453 2283 15487
rect 4614 15484 4620 15496
rect 4575 15456 4620 15484
rect 2225 15447 2283 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 7282 15484 7288 15496
rect 7243 15456 7288 15484
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 9030 15484 9036 15496
rect 8720 15456 9036 15484
rect 8720 15444 8726 15456
rect 9030 15444 9036 15456
rect 9088 15484 9094 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 9088 15456 10149 15484
rect 9088 15444 9094 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 7190 15348 7196 15360
rect 7151 15320 7196 15348
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 10244 15348 10272 15524
rect 10321 15487 10379 15493
rect 10321 15453 10333 15487
rect 10367 15484 10379 15487
rect 10410 15484 10416 15496
rect 10367 15456 10416 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 10980 15416 11008 15648
rect 11422 15580 11428 15632
rect 11480 15629 11486 15632
rect 11480 15623 11544 15629
rect 11480 15589 11498 15623
rect 11532 15620 11544 15623
rect 11698 15620 11704 15632
rect 11532 15592 11704 15620
rect 11532 15589 11544 15592
rect 11480 15583 11544 15589
rect 11480 15580 11486 15583
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 12452 15620 12480 15660
rect 12618 15648 12624 15660
rect 12676 15688 12682 15700
rect 13262 15688 13268 15700
rect 12676 15660 13268 15688
rect 12676 15648 12682 15660
rect 13262 15648 13268 15660
rect 13320 15648 13326 15700
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 14090 15648 14096 15660
rect 14148 15688 14154 15700
rect 14148 15660 14780 15688
rect 14148 15648 14154 15660
rect 14645 15623 14703 15629
rect 14645 15620 14657 15623
rect 12452 15592 14657 15620
rect 14645 15589 14657 15592
rect 14691 15589 14703 15623
rect 14645 15583 14703 15589
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 12584 15524 12725 15552
rect 12584 15512 12590 15524
rect 12713 15521 12725 15524
rect 12759 15521 12771 15555
rect 12713 15515 12771 15521
rect 12980 15555 13038 15561
rect 12980 15521 12992 15555
rect 13026 15552 13038 15555
rect 13262 15552 13268 15564
rect 13026 15524 13268 15552
rect 13026 15521 13038 15524
rect 12980 15515 13038 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 14550 15552 14556 15564
rect 14511 15524 14556 15552
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 14752 15493 14780 15660
rect 11241 15487 11299 15493
rect 11241 15484 11253 15487
rect 11112 15456 11253 15484
rect 11112 15444 11118 15456
rect 11241 15453 11253 15456
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14182 15416 14188 15428
rect 10980 15388 11192 15416
rect 14143 15388 14188 15416
rect 10962 15348 10968 15360
rect 10244 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15348 11026 15360
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 11020 15320 11069 15348
rect 11020 15308 11026 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11164 15348 11192 15388
rect 14182 15376 14188 15388
rect 14240 15376 14246 15428
rect 13998 15348 14004 15360
rect 11164 15320 14004 15348
rect 11057 15311 11115 15317
rect 13998 15308 14004 15320
rect 14056 15308 14062 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5905 15147 5963 15153
rect 5905 15144 5917 15147
rect 5592 15116 5917 15144
rect 5592 15104 5598 15116
rect 5905 15113 5917 15116
rect 5951 15113 5963 15147
rect 5905 15107 5963 15113
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 8665 15147 8723 15153
rect 8665 15144 8677 15147
rect 6696 15116 8677 15144
rect 6696 15104 6702 15116
rect 8665 15113 8677 15116
rect 8711 15113 8723 15147
rect 8938 15144 8944 15156
rect 8899 15116 8944 15144
rect 8665 15107 8723 15113
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 7929 15079 7987 15085
rect 7929 15076 7941 15079
rect 5776 15048 7941 15076
rect 5776 15036 5782 15048
rect 7929 15045 7941 15048
rect 7975 15045 7987 15079
rect 7929 15039 7987 15045
rect 2866 15008 2872 15020
rect 2056 14980 2728 15008
rect 2827 14980 2872 15008
rect 2056 14949 2084 14980
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14909 2099 14943
rect 2314 14940 2320 14952
rect 2275 14912 2320 14940
rect 2041 14903 2099 14909
rect 2314 14900 2320 14912
rect 2372 14900 2378 14952
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 2700 14940 2728 14980
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 15008 3847 15011
rect 3878 15008 3884 15020
rect 3835 14980 3884 15008
rect 3835 14977 3847 14980
rect 3789 14971 3847 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 7190 15008 7196 15020
rect 6595 14980 7196 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 8680 15008 8708 15107
rect 8938 15104 8944 15116
rect 8996 15144 9002 15156
rect 8996 15116 9536 15144
rect 8996 15104 9002 15116
rect 9033 15079 9091 15085
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 9214 15076 9220 15088
rect 9079 15048 9220 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 9214 15036 9220 15048
rect 9272 15036 9278 15088
rect 9508 15020 9536 15116
rect 9858 15104 9864 15156
rect 9916 15144 9922 15156
rect 11054 15144 11060 15156
rect 9916 15116 11060 15144
rect 9916 15104 9922 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11333 15147 11391 15153
rect 11333 15144 11345 15147
rect 11296 15116 11345 15144
rect 11296 15104 11302 15116
rect 11333 15113 11345 15116
rect 11379 15113 11391 15147
rect 13170 15144 13176 15156
rect 11333 15107 11391 15113
rect 11808 15116 13176 15144
rect 9122 15008 9128 15020
rect 8680 14980 9128 15008
rect 7377 14971 7435 14977
rect 2700 14912 3832 14940
rect 2593 14903 2651 14909
rect 2608 14804 2636 14903
rect 3804 14884 3832 14912
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7392 14940 7420 14971
rect 9122 14968 9128 14980
rect 9180 15008 9186 15020
rect 9180 14980 9444 15008
rect 9180 14968 9186 14980
rect 6972 14912 7420 14940
rect 8113 14943 8171 14949
rect 6972 14900 6978 14912
rect 8113 14909 8125 14943
rect 8159 14940 8171 14943
rect 9030 14940 9036 14952
rect 8159 14912 9036 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9416 14949 9444 14980
rect 9490 14968 9496 15020
rect 9548 15008 9554 15020
rect 9677 15011 9735 15017
rect 9548 14980 9641 15008
rect 9548 14968 9554 14980
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 9723 14980 9996 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14909 9459 14943
rect 9858 14940 9864 14952
rect 9819 14912 9864 14940
rect 9401 14903 9459 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 9968 14940 9996 14980
rect 10870 14968 10876 15020
rect 10928 15008 10934 15020
rect 11808 15008 11836 15116
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 14550 15144 14556 15156
rect 13403 15116 14556 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 14182 15076 14188 15088
rect 12360 15048 14188 15076
rect 11974 15008 11980 15020
rect 10928 14980 11836 15008
rect 11935 14980 11980 15008
rect 10928 14968 10934 14980
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 10128 14943 10186 14949
rect 10128 14940 10140 14943
rect 9968 14912 10140 14940
rect 10128 14909 10140 14912
rect 10174 14940 10186 14943
rect 10410 14940 10416 14952
rect 10174 14912 10416 14940
rect 10174 14909 10186 14912
rect 10128 14903 10186 14909
rect 10410 14900 10416 14912
rect 10468 14940 10474 14952
rect 11992 14940 12020 14968
rect 10468 14912 12020 14940
rect 10468 14900 10474 14912
rect 3786 14832 3792 14884
rect 3844 14832 3850 14884
rect 6273 14875 6331 14881
rect 6273 14841 6285 14875
rect 6319 14872 6331 14875
rect 7193 14875 7251 14881
rect 6319 14844 6868 14872
rect 6319 14841 6331 14844
rect 6273 14835 6331 14841
rect 3145 14807 3203 14813
rect 3145 14804 3157 14807
rect 2608 14776 3157 14804
rect 3145 14773 3157 14776
rect 3191 14773 3203 14807
rect 3145 14767 3203 14773
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 3513 14807 3571 14813
rect 3513 14804 3525 14807
rect 3384 14776 3525 14804
rect 3384 14764 3390 14776
rect 3513 14773 3525 14776
rect 3559 14773 3571 14807
rect 3513 14767 3571 14773
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 6362 14804 6368 14816
rect 3660 14776 3705 14804
rect 6323 14776 6368 14804
rect 3660 14764 3666 14776
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6840 14813 6868 14844
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 7239 14844 7665 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7653 14841 7665 14844
rect 7699 14841 7711 14875
rect 7653 14835 7711 14841
rect 9214 14832 9220 14884
rect 9272 14872 9278 14884
rect 10686 14872 10692 14884
rect 9272 14844 10692 14872
rect 9272 14832 9278 14844
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 10962 14832 10968 14884
rect 11020 14872 11026 14884
rect 11701 14875 11759 14881
rect 11701 14872 11713 14875
rect 11020 14844 11713 14872
rect 11020 14832 11026 14844
rect 11701 14841 11713 14844
rect 11747 14872 11759 14875
rect 11882 14872 11888 14884
rect 11747 14844 11888 14872
rect 11747 14841 11759 14844
rect 11701 14835 11759 14841
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7064 14776 7297 14804
rect 7064 14764 7070 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 7285 14767 7343 14773
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 10778 14804 10784 14816
rect 8536 14776 10784 14804
rect 8536 14764 8542 14776
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11238 14804 11244 14816
rect 11112 14776 11244 14804
rect 11112 14764 11118 14776
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11793 14807 11851 14813
rect 11793 14804 11805 14807
rect 11388 14776 11805 14804
rect 11388 14764 11394 14776
rect 11793 14773 11805 14776
rect 11839 14804 11851 14807
rect 12360 14804 12388 15048
rect 14182 15036 14188 15048
rect 14240 15036 14246 15088
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12584 14980 13093 15008
rect 12584 14968 12590 14980
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13320 14980 13921 15008
rect 13320 14968 13326 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14940 12955 14943
rect 13538 14940 13544 14952
rect 12943 14912 13544 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 13538 14900 13544 14912
rect 13596 14900 13602 14952
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 13872 14912 13917 14940
rect 13872 14900 13878 14912
rect 14090 14900 14096 14952
rect 14148 14940 14154 14952
rect 14642 14949 14648 14952
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 14148 14912 14381 14940
rect 14148 14900 14154 14912
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 14636 14940 14648 14949
rect 14603 14912 14648 14940
rect 14369 14903 14427 14909
rect 14636 14903 14648 14912
rect 14642 14900 14648 14903
rect 14700 14900 14706 14952
rect 13446 14872 13452 14884
rect 12544 14844 13452 14872
rect 12544 14813 12572 14844
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 13722 14832 13728 14884
rect 13780 14872 13786 14884
rect 18782 14872 18788 14884
rect 13780 14844 13825 14872
rect 15212 14844 18788 14872
rect 13780 14832 13786 14844
rect 11839 14776 12388 14804
rect 12529 14807 12587 14813
rect 11839 14773 11851 14776
rect 11793 14767 11851 14773
rect 12529 14773 12541 14807
rect 12575 14773 12587 14807
rect 12529 14767 12587 14773
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13078 14804 13084 14816
rect 13035 14776 13084 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13170 14764 13176 14816
rect 13228 14804 13234 14816
rect 15212 14804 15240 14844
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 13228 14776 15240 14804
rect 13228 14764 13234 14776
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 15749 14807 15807 14813
rect 15749 14804 15761 14807
rect 15344 14776 15761 14804
rect 15344 14764 15350 14776
rect 15749 14773 15761 14776
rect 15795 14773 15807 14807
rect 15749 14767 15807 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2317 14603 2375 14609
rect 2317 14569 2329 14603
rect 2363 14600 2375 14603
rect 2774 14600 2780 14612
rect 2363 14572 2780 14600
rect 2363 14569 2375 14572
rect 2317 14563 2375 14569
rect 2774 14560 2780 14572
rect 2832 14560 2838 14612
rect 3878 14600 3884 14612
rect 3839 14572 3884 14600
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 3896 14532 3924 14560
rect 4310 14535 4368 14541
rect 4310 14532 4322 14535
rect 3896 14504 4322 14532
rect 4310 14501 4322 14504
rect 4356 14501 4368 14535
rect 5460 14532 5488 14563
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 6420 14572 7205 14600
rect 6420 14560 6426 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7699 14572 8217 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 8665 14603 8723 14609
rect 8665 14569 8677 14603
rect 8711 14600 8723 14603
rect 9030 14600 9036 14612
rect 8711 14572 8892 14600
rect 8991 14572 9036 14600
rect 8711 14569 8723 14572
rect 8665 14563 8723 14569
rect 5804 14535 5862 14541
rect 5804 14532 5816 14535
rect 5460 14504 5816 14532
rect 4310 14495 4368 14501
rect 5804 14501 5816 14504
rect 5850 14532 5862 14535
rect 5850 14504 8800 14532
rect 5850 14501 5862 14504
rect 5804 14495 5862 14501
rect 1765 14467 1823 14473
rect 1765 14433 1777 14467
rect 1811 14433 1823 14467
rect 2130 14464 2136 14476
rect 2091 14436 2136 14464
rect 1765 14427 1823 14433
rect 1780 14396 1808 14427
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 2768 14467 2826 14473
rect 2768 14433 2780 14467
rect 2814 14464 2826 14467
rect 3878 14464 3884 14476
rect 2814 14436 3884 14464
rect 2814 14433 2826 14436
rect 2768 14427 2826 14433
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 7650 14464 7656 14476
rect 7607 14436 7656 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 7650 14424 7656 14436
rect 7708 14464 7714 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 7708 14436 8033 14464
rect 7708 14424 7714 14436
rect 8021 14433 8033 14436
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14433 8631 14467
rect 8573 14427 8631 14433
rect 2314 14396 2320 14408
rect 1780 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14365 2559 14399
rect 2501 14359 2559 14365
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 5534 14396 5540 14408
rect 5495 14368 5540 14396
rect 4065 14359 4123 14365
rect 2038 14288 2044 14340
rect 2096 14328 2102 14340
rect 2516 14328 2544 14359
rect 2096 14300 2544 14328
rect 2096 14288 2102 14300
rect 2516 14260 2544 14300
rect 4080 14272 4108 14359
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 7745 14399 7803 14405
rect 7745 14365 7757 14399
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 6914 14328 6920 14340
rect 6875 14300 6920 14328
rect 6914 14288 6920 14300
rect 6972 14328 6978 14340
rect 7760 14328 7788 14359
rect 6972 14300 7788 14328
rect 8588 14328 8616 14427
rect 8772 14405 8800 14504
rect 8757 14399 8815 14405
rect 8757 14365 8769 14399
rect 8803 14365 8815 14399
rect 8864 14396 8892 14572
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 9401 14603 9459 14609
rect 9401 14569 9413 14603
rect 9447 14600 9459 14603
rect 9493 14603 9551 14609
rect 9493 14600 9505 14603
rect 9447 14572 9505 14600
rect 9447 14569 9459 14572
rect 9401 14563 9459 14569
rect 9493 14569 9505 14572
rect 9539 14600 9551 14603
rect 9674 14600 9680 14612
rect 9539 14572 9680 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9674 14560 9680 14572
rect 9732 14600 9738 14612
rect 10870 14600 10876 14612
rect 9732 14572 10876 14600
rect 9732 14560 9738 14572
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 11020 14572 11529 14600
rect 11020 14560 11026 14572
rect 11517 14569 11529 14572
rect 11563 14569 11575 14603
rect 11517 14563 11575 14569
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 13078 14600 13084 14612
rect 12667 14572 12940 14600
rect 13039 14572 13084 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 9048 14532 9076 14560
rect 9048 14504 10456 14532
rect 9214 14464 9220 14476
rect 9175 14436 9220 14464
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9398 14424 9404 14476
rect 9456 14464 9462 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9456 14436 9689 14464
rect 9456 14424 9462 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9416 14396 9444 14424
rect 8864 14368 9444 14396
rect 8757 14359 8815 14365
rect 9493 14331 9551 14337
rect 9493 14328 9505 14331
rect 8588 14300 9505 14328
rect 6972 14288 6978 14300
rect 9493 14297 9505 14300
rect 9539 14297 9551 14331
rect 9692 14328 9720 14427
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 9953 14467 10011 14473
rect 9953 14464 9965 14467
rect 9916 14436 9965 14464
rect 9916 14424 9922 14436
rect 9953 14433 9965 14436
rect 9999 14464 10011 14467
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 9999 14436 10149 14464
rect 9999 14433 10011 14436
rect 9953 14427 10011 14433
rect 10137 14433 10149 14436
rect 10183 14464 10195 14467
rect 10318 14464 10324 14476
rect 10183 14436 10324 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 10428 14473 10456 14504
rect 10778 14492 10784 14544
rect 10836 14532 10842 14544
rect 11330 14532 11336 14544
rect 10836 14504 11336 14532
rect 10836 14492 10842 14504
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 12713 14535 12771 14541
rect 12713 14501 12725 14535
rect 12759 14532 12771 14535
rect 12802 14532 12808 14544
rect 12759 14504 12808 14532
rect 12759 14501 12771 14504
rect 12713 14495 12771 14501
rect 12802 14492 12808 14504
rect 12860 14492 12866 14544
rect 12912 14532 12940 14572
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 13722 14600 13728 14612
rect 13228 14572 13728 14600
rect 13228 14560 13234 14572
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 14240 14572 14657 14600
rect 14240 14560 14246 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 14645 14563 14703 14569
rect 15381 14603 15439 14609
rect 15381 14569 15393 14603
rect 15427 14600 15439 14603
rect 15562 14600 15568 14612
rect 15427 14572 15568 14600
rect 15427 14569 15439 14572
rect 15381 14563 15439 14569
rect 15562 14560 15568 14572
rect 15620 14600 15626 14612
rect 22738 14600 22744 14612
rect 15620 14572 22744 14600
rect 15620 14560 15626 14572
rect 22738 14560 22744 14572
rect 22796 14560 22802 14612
rect 13446 14532 13452 14544
rect 12912 14504 13216 14532
rect 13407 14504 13452 14532
rect 10413 14467 10471 14473
rect 10413 14433 10425 14467
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 10870 14464 10876 14476
rect 10652 14436 10876 14464
rect 10652 14424 10658 14436
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12526 14464 12532 14476
rect 11756 14436 12532 14464
rect 11756 14424 11762 14436
rect 12526 14424 12532 14436
rect 12584 14464 12590 14476
rect 12584 14436 12848 14464
rect 12584 14424 12590 14436
rect 10336 14396 10364 14424
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10336 14368 10977 14396
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11974 14396 11980 14408
rect 11195 14368 11980 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 12820 14405 12848 14436
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14365 12863 14399
rect 13188 14396 13216 14504
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 13909 14535 13967 14541
rect 13909 14532 13921 14535
rect 13556 14504 13921 14532
rect 13556 14464 13584 14504
rect 13909 14501 13921 14504
rect 13955 14501 13967 14535
rect 14550 14532 14556 14544
rect 14511 14504 14556 14532
rect 13909 14495 13967 14501
rect 14550 14492 14556 14504
rect 14608 14532 14614 14544
rect 15013 14535 15071 14541
rect 15013 14532 15025 14535
rect 14608 14504 15025 14532
rect 14608 14492 14614 14504
rect 15013 14501 15025 14504
rect 15059 14501 15071 14535
rect 15013 14495 15071 14501
rect 14366 14464 14372 14476
rect 13464 14436 13584 14464
rect 13648 14436 14372 14464
rect 13464 14396 13492 14436
rect 13188 14368 13492 14396
rect 13541 14399 13599 14405
rect 12805 14359 12863 14365
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13648 14396 13676 14436
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 13587 14368 13676 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 11238 14328 11244 14340
rect 9692 14300 11244 14328
rect 9493 14291 9551 14297
rect 11238 14288 11244 14300
rect 11296 14288 11302 14340
rect 12253 14331 12311 14337
rect 12253 14297 12265 14331
rect 12299 14328 12311 14331
rect 13170 14328 13176 14340
rect 12299 14300 13176 14328
rect 12299 14297 12311 14300
rect 12253 14291 12311 14297
rect 13170 14288 13176 14300
rect 13228 14288 13234 14340
rect 4062 14260 4068 14272
rect 2516 14232 4068 14260
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 7006 14260 7012 14272
rect 6967 14232 7012 14260
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 10226 14260 10232 14272
rect 10187 14232 10232 14260
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 10505 14263 10563 14269
rect 10505 14229 10517 14263
rect 10551 14260 10563 14263
rect 10778 14260 10784 14272
rect 10551 14232 10784 14260
rect 10551 14229 10563 14232
rect 10505 14223 10563 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 12069 14263 12127 14269
rect 12069 14260 12081 14263
rect 12032 14232 12081 14260
rect 12032 14220 12038 14232
rect 12069 14229 12081 14232
rect 12115 14260 12127 14263
rect 12618 14260 12624 14272
rect 12115 14232 12624 14260
rect 12115 14229 12127 14232
rect 12069 14223 12127 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 13556 14260 13584 14359
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 13780 14368 13825 14396
rect 13780 14356 13786 14368
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 14792 14368 14837 14396
rect 14792 14356 14798 14368
rect 13136 14232 13584 14260
rect 14185 14263 14243 14269
rect 13136 14220 13142 14232
rect 14185 14229 14197 14263
rect 14231 14260 14243 14263
rect 15102 14260 15108 14272
rect 14231 14232 15108 14260
rect 14231 14229 14243 14232
rect 14185 14223 14243 14229
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3326 14056 3332 14068
rect 2832 14028 2877 14056
rect 3287 14028 3332 14056
rect 2832 14016 2838 14028
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 3660 14028 4721 14056
rect 3660 14016 3666 14028
rect 4709 14025 4721 14028
rect 4755 14025 4767 14059
rect 9306 14056 9312 14068
rect 4709 14019 4767 14025
rect 7668 14028 9312 14056
rect 3878 13920 3884 13932
rect 2056 13892 3740 13920
rect 3839 13892 3884 13920
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2056 13861 2084 13892
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2314 13852 2320 13864
rect 2275 13824 2320 13852
rect 2041 13815 2099 13821
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 2498 13812 2504 13864
rect 2556 13852 2562 13864
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2556 13824 2605 13852
rect 2556 13812 2562 13824
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 3712 13852 3740 13892
rect 3878 13880 3884 13892
rect 3936 13920 3942 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 3936 13892 5273 13920
rect 3936 13880 3942 13892
rect 5261 13889 5273 13892
rect 5307 13920 5319 13923
rect 5810 13920 5816 13932
rect 5307 13892 5816 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7668 13929 7696 14028
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 10321 14059 10379 14065
rect 10321 14025 10333 14059
rect 10367 14056 10379 14059
rect 11146 14056 11152 14068
rect 10367 14028 11152 14056
rect 10367 14025 10379 14028
rect 10321 14019 10379 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13170 14056 13176 14068
rect 12952 14028 13176 14056
rect 12952 14016 12958 14028
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 13538 14056 13544 14068
rect 13499 14028 13544 14056
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 14369 14059 14427 14065
rect 14369 14056 14381 14059
rect 14016 14028 14381 14056
rect 10060 13960 13400 13988
rect 7653 13923 7711 13929
rect 7653 13920 7665 13923
rect 7248 13892 7665 13920
rect 7248 13880 7254 13892
rect 7653 13889 7665 13892
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 10060 13929 10088 13960
rect 10045 13923 10103 13929
rect 10045 13920 10057 13923
rect 8996 13892 10057 13920
rect 8996 13880 9002 13892
rect 10045 13889 10057 13892
rect 10091 13889 10103 13923
rect 10778 13920 10784 13932
rect 10739 13892 10784 13920
rect 10045 13883 10103 13889
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11054 13920 11060 13932
rect 11011 13892 11060 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 13372 13929 13400 13960
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 4798 13852 4804 13864
rect 3712 13824 4804 13852
rect 2593 13815 2651 13821
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 5169 13855 5227 13861
rect 5169 13821 5181 13855
rect 5215 13852 5227 13855
rect 5626 13852 5632 13864
rect 5215 13824 5632 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 5718 13812 5724 13864
rect 5776 13852 5782 13864
rect 5905 13855 5963 13861
rect 5776 13824 5821 13852
rect 5776 13812 5782 13824
rect 5905 13821 5917 13855
rect 5951 13852 5963 13855
rect 6086 13852 6092 13864
rect 5951 13824 6092 13852
rect 5951 13821 5963 13824
rect 5905 13815 5963 13821
rect 3697 13787 3755 13793
rect 3697 13753 3709 13787
rect 3743 13784 3755 13787
rect 4157 13787 4215 13793
rect 4157 13784 4169 13787
rect 3743 13756 4169 13784
rect 3743 13753 3755 13756
rect 3697 13747 3755 13753
rect 4157 13753 4169 13756
rect 4203 13753 4215 13787
rect 4157 13747 4215 13753
rect 5077 13787 5135 13793
rect 5077 13753 5089 13787
rect 5123 13784 5135 13787
rect 5920 13784 5948 13815
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13852 7619 13855
rect 7834 13852 7840 13864
rect 7607 13824 7840 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13852 7987 13855
rect 8018 13852 8024 13864
rect 7975 13824 8024 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 8956 13852 8984 13880
rect 9858 13852 9864 13864
rect 8312 13824 8984 13852
rect 9819 13824 9864 13852
rect 5123 13756 5948 13784
rect 7469 13787 7527 13793
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 7469 13753 7481 13787
rect 7515 13784 7527 13787
rect 8196 13787 8254 13793
rect 7515 13756 7880 13784
rect 7515 13753 7527 13756
rect 7469 13747 7527 13753
rect 2958 13676 2964 13728
rect 3016 13716 3022 13728
rect 3237 13719 3295 13725
rect 3237 13716 3249 13719
rect 3016 13688 3249 13716
rect 3016 13676 3022 13688
rect 3237 13685 3249 13688
rect 3283 13716 3295 13719
rect 3789 13719 3847 13725
rect 3789 13716 3801 13719
rect 3283 13688 3801 13716
rect 3283 13685 3295 13688
rect 3237 13679 3295 13685
rect 3789 13685 3801 13688
rect 3835 13716 3847 13719
rect 3878 13716 3884 13728
rect 3835 13688 3884 13716
rect 3835 13685 3847 13688
rect 3789 13679 3847 13685
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 5534 13716 5540 13728
rect 4120 13688 5540 13716
rect 4120 13676 4126 13688
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 7098 13716 7104 13728
rect 7059 13688 7104 13716
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 7852 13716 7880 13756
rect 8196 13753 8208 13787
rect 8242 13784 8254 13787
rect 8312 13784 8340 13824
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 10284 13824 12081 13852
rect 10284 13812 10290 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12069 13815 12127 13821
rect 12176 13824 13093 13852
rect 8242 13756 8340 13784
rect 8242 13753 8254 13756
rect 8196 13747 8254 13753
rect 9490 13744 9496 13796
rect 9548 13784 9554 13796
rect 9769 13787 9827 13793
rect 9769 13784 9781 13787
rect 9548 13756 9781 13784
rect 9548 13744 9554 13756
rect 9769 13753 9781 13756
rect 9815 13753 9827 13787
rect 10686 13784 10692 13796
rect 10647 13756 10692 13784
rect 9769 13747 9827 13753
rect 9401 13719 9459 13725
rect 9401 13716 9413 13719
rect 7852 13688 9413 13716
rect 9401 13685 9413 13688
rect 9447 13685 9459 13719
rect 9784 13716 9812 13747
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 12176 13793 12204 13824
rect 13081 13821 13093 13824
rect 13127 13852 13139 13855
rect 13262 13852 13268 13864
rect 13127 13824 13268 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13372 13852 13400 13883
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14016 13929 14044 14028
rect 14369 14025 14381 14028
rect 14415 14056 14427 14059
rect 14458 14056 14464 14068
rect 14415 14028 14464 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 15562 14056 15568 14068
rect 15523 14028 15568 14056
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 14645 13991 14703 13997
rect 14645 13957 14657 13991
rect 14691 13988 14703 13991
rect 15746 13988 15752 14000
rect 14691 13960 15752 13988
rect 14691 13957 14703 13960
rect 14645 13951 14703 13957
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13504 13892 14013 13920
rect 13504 13880 13510 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 14185 13883 14243 13889
rect 13538 13852 13544 13864
rect 13372 13824 13544 13852
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14200 13852 14228 13883
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15286 13920 15292 13932
rect 15247 13892 15292 13920
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 13688 13824 14228 13852
rect 13688 13812 13694 13824
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 15013 13855 15071 13861
rect 15013 13852 15025 13855
rect 14424 13824 15025 13852
rect 14424 13812 14430 13824
rect 15013 13821 15025 13824
rect 15059 13852 15071 13855
rect 15562 13852 15568 13864
rect 15059 13824 15568 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 12161 13787 12219 13793
rect 12161 13784 12173 13787
rect 10836 13756 12173 13784
rect 10836 13744 10842 13756
rect 12161 13753 12173 13756
rect 12207 13753 12219 13787
rect 12161 13747 12219 13753
rect 12621 13787 12679 13793
rect 12621 13753 12633 13787
rect 12667 13784 12679 13787
rect 12802 13784 12808 13796
rect 12667 13756 12808 13784
rect 12667 13753 12679 13756
rect 12621 13747 12679 13753
rect 12802 13744 12808 13756
rect 12860 13784 12866 13796
rect 13909 13787 13967 13793
rect 13909 13784 13921 13787
rect 12860 13756 13921 13784
rect 12860 13744 12866 13756
rect 13909 13753 13921 13756
rect 13955 13753 13967 13787
rect 18046 13784 18052 13796
rect 13909 13747 13967 13753
rect 14007 13756 18052 13784
rect 11149 13719 11207 13725
rect 11149 13716 11161 13719
rect 9784 13688 11161 13716
rect 9401 13679 9459 13685
rect 11149 13685 11161 13688
rect 11195 13685 11207 13719
rect 11149 13679 11207 13685
rect 11514 13676 11520 13728
rect 11572 13716 11578 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11572 13688 11897 13716
rect 11572 13676 11578 13688
rect 11885 13685 11897 13688
rect 11931 13685 11943 13719
rect 12710 13716 12716 13728
rect 12671 13688 12716 13716
rect 11885 13679 11943 13685
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13173 13719 13231 13725
rect 13173 13716 13185 13719
rect 13136 13688 13185 13716
rect 13136 13676 13142 13688
rect 13173 13685 13185 13688
rect 13219 13685 13231 13719
rect 13173 13679 13231 13685
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 14007 13716 14035 13756
rect 18046 13744 18052 13756
rect 18104 13744 18110 13796
rect 13320 13688 14035 13716
rect 13320 13676 13326 13688
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 1762 13512 1768 13524
rect 1723 13484 1768 13512
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2455 13484 2881 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 5684 13484 6009 13512
rect 5684 13472 5690 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 5997 13475 6055 13481
rect 6365 13515 6423 13521
rect 6365 13481 6377 13515
rect 6411 13512 6423 13515
rect 6411 13484 6960 13512
rect 6411 13481 6423 13484
rect 6365 13475 6423 13481
rect 4792 13447 4850 13453
rect 4792 13413 4804 13447
rect 4838 13444 4850 13447
rect 5534 13444 5540 13456
rect 4838 13416 5540 13444
rect 4838 13413 4850 13416
rect 4792 13407 4850 13413
rect 5534 13404 5540 13416
rect 5592 13444 5598 13456
rect 5592 13416 6684 13444
rect 5592 13404 5598 13416
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13345 1639 13379
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 1581 13339 1639 13345
rect 1596 13308 1624 13339
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 3234 13376 3240 13388
rect 3195 13348 3240 13376
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4120 13348 4537 13376
rect 4120 13336 4126 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 2406 13308 2412 13320
rect 1596 13280 2412 13308
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 2590 13308 2596 13320
rect 2551 13280 2596 13308
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 3326 13308 3332 13320
rect 3287 13280 3332 13308
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3510 13308 3516 13320
rect 3471 13280 3516 13308
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 6656 13317 6684 13416
rect 6932 13385 6960 13484
rect 7098 13472 7104 13524
rect 7156 13512 7162 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 7156 13484 7757 13512
rect 7156 13472 7162 13484
rect 7745 13481 7757 13484
rect 7791 13481 7803 13515
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 7745 13475 7803 13481
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8662 13512 8668 13524
rect 8623 13484 8668 13512
rect 8662 13472 8668 13484
rect 8720 13512 8726 13524
rect 9125 13515 9183 13521
rect 9125 13512 9137 13515
rect 8720 13484 9137 13512
rect 8720 13472 8726 13484
rect 9125 13481 9137 13484
rect 9171 13481 9183 13515
rect 9125 13475 9183 13481
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 9456 13484 9505 13512
rect 9456 13472 9462 13484
rect 9493 13481 9505 13484
rect 9539 13512 9551 13515
rect 9582 13512 9588 13524
rect 9539 13484 9588 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 7653 13447 7711 13453
rect 7653 13413 7665 13447
rect 7699 13444 7711 13447
rect 9692 13444 9720 13475
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 9916 13484 10057 13512
rect 9916 13472 9922 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 12710 13512 12716 13524
rect 10183 13484 12716 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12952 13484 13001 13512
rect 12952 13472 12958 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 14277 13515 14335 13521
rect 13596 13484 14228 13512
rect 13596 13472 13602 13484
rect 7699 13416 9720 13444
rect 7699 13413 7711 13416
rect 7653 13407 7711 13413
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 14090 13444 14096 13456
rect 9824 13416 14096 13444
rect 9824 13404 9830 13416
rect 14090 13404 14096 13416
rect 14148 13404 14154 13456
rect 14200 13444 14228 13484
rect 14277 13481 14289 13515
rect 14323 13512 14335 13515
rect 14366 13512 14372 13524
rect 14323 13484 14372 13512
rect 14323 13481 14335 13484
rect 14277 13475 14335 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15746 13512 15752 13524
rect 15707 13484 15752 13512
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 17773 13515 17831 13521
rect 17773 13481 17785 13515
rect 17819 13481 17831 13515
rect 17773 13475 17831 13481
rect 17788 13444 17816 13475
rect 14200 13416 17816 13444
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 9122 13376 9128 13388
rect 6963 13348 9128 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 9122 13336 9128 13348
rect 9180 13376 9186 13388
rect 11606 13376 11612 13388
rect 9180 13348 11612 13376
rect 9180 13336 9186 13348
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 11784 13379 11842 13385
rect 11784 13345 11796 13379
rect 11830 13376 11842 13379
rect 12066 13376 12072 13388
rect 11830 13348 12072 13376
rect 11830 13345 11842 13348
rect 11784 13339 11842 13345
rect 12066 13336 12072 13348
rect 12124 13336 12130 13388
rect 12710 13336 12716 13388
rect 12768 13376 12774 13388
rect 12894 13376 12900 13388
rect 12768 13348 12900 13376
rect 12768 13336 12774 13348
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 13354 13376 13360 13388
rect 13267 13348 13360 13376
rect 13354 13336 13360 13348
rect 13412 13376 13418 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13412 13348 14013 13376
rect 13412 13336 13418 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 14001 13339 14059 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16660 13379 16718 13385
rect 16660 13345 16672 13379
rect 16706 13376 16718 13379
rect 16706 13348 18000 13376
rect 16706 13345 16718 13348
rect 16660 13339 16718 13345
rect 6457 13311 6515 13317
rect 6457 13277 6469 13311
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 7834 13308 7840 13320
rect 7795 13280 7840 13308
rect 6641 13271 6699 13277
rect 5810 13200 5816 13252
rect 5868 13240 5874 13252
rect 5905 13243 5963 13249
rect 5905 13240 5917 13243
rect 5868 13212 5917 13240
rect 5868 13200 5874 13212
rect 5905 13209 5917 13212
rect 5951 13209 5963 13243
rect 6472 13240 6500 13271
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8478 13308 8484 13320
rect 8251 13280 8484 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8478 13268 8484 13280
rect 8536 13308 8542 13320
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 8536 13280 8769 13308
rect 8536 13268 8542 13280
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8938 13308 8944 13320
rect 8899 13280 8944 13308
rect 8757 13271 8815 13277
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9364 13280 10241 13308
rect 9364 13268 9370 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 10962 13308 10968 13320
rect 10643 13280 10968 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11514 13308 11520 13320
rect 11204 13280 11520 13308
rect 11204 13268 11210 13280
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 13449 13311 13507 13317
rect 13449 13308 13461 13311
rect 12676 13280 13461 13308
rect 12676 13268 12682 13280
rect 13449 13277 13461 13280
rect 13495 13277 13507 13311
rect 13630 13308 13636 13320
rect 13591 13280 13636 13308
rect 13449 13271 13507 13277
rect 6730 13240 6736 13252
rect 6472 13212 6736 13240
rect 5905 13203 5963 13209
rect 6730 13200 6736 13212
rect 6788 13240 6794 13252
rect 7101 13243 7159 13249
rect 7101 13240 7113 13243
rect 6788 13212 7113 13240
rect 6788 13200 6794 13212
rect 7101 13209 7113 13212
rect 7147 13240 7159 13243
rect 8386 13240 8392 13252
rect 7147 13212 8392 13240
rect 7147 13209 7159 13212
rect 7101 13203 7159 13209
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 13354 13240 13360 13252
rect 12636 13212 13360 13240
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13172 2007 13175
rect 2866 13172 2872 13184
rect 1995 13144 2872 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 7282 13172 7288 13184
rect 7243 13144 7288 13172
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 12636 13172 12664 13212
rect 13354 13200 13360 13212
rect 13412 13200 13418 13252
rect 13464 13240 13492 13271
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 13817 13243 13875 13249
rect 13817 13240 13829 13243
rect 13464 13212 13829 13240
rect 13817 13209 13829 13212
rect 13863 13209 13875 13243
rect 13817 13203 13875 13209
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 16408 13240 16436 13271
rect 14240 13212 16436 13240
rect 14240 13200 14246 13212
rect 9640 13144 12664 13172
rect 9640 13132 9646 13144
rect 12710 13132 12716 13184
rect 12768 13172 12774 13184
rect 12897 13175 12955 13181
rect 12897 13172 12909 13175
rect 12768 13144 12909 13172
rect 12768 13132 12774 13144
rect 12897 13141 12909 13144
rect 12943 13141 12955 13175
rect 12897 13135 12955 13141
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15746 13172 15752 13184
rect 15335 13144 15752 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 17972 13181 18000 13348
rect 17957 13175 18015 13181
rect 17957 13141 17969 13175
rect 18003 13172 18015 13175
rect 18598 13172 18604 13184
rect 18003 13144 18604 13172
rect 18003 13141 18015 13144
rect 17957 13135 18015 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 3513 12931 3571 12937
rect 3804 12940 4629 12968
rect 2406 12792 2412 12844
rect 2464 12832 2470 12844
rect 3053 12835 3111 12841
rect 3053 12832 3065 12835
rect 2464 12804 3065 12832
rect 2464 12792 2470 12804
rect 3053 12801 3065 12804
rect 3099 12801 3111 12835
rect 3053 12795 3111 12801
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2038 12764 2044 12776
rect 1443 12736 2044 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 2866 12764 2872 12776
rect 2827 12736 2872 12764
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 1664 12699 1722 12705
rect 1664 12665 1676 12699
rect 1710 12696 1722 12699
rect 2222 12696 2228 12708
rect 1710 12668 2228 12696
rect 1710 12665 1722 12668
rect 1664 12659 1722 12665
rect 2222 12656 2228 12668
rect 2280 12696 2286 12708
rect 3510 12696 3516 12708
rect 2280 12668 3516 12696
rect 2280 12656 2286 12668
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 3804 12696 3832 12940
rect 4617 12937 4629 12940
rect 4663 12968 4675 12971
rect 4982 12968 4988 12980
rect 4663 12940 4988 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 9766 12968 9772 12980
rect 5092 12940 9772 12968
rect 3878 12860 3884 12912
rect 3936 12900 3942 12912
rect 5092 12900 5120 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 13630 12928 13636 12980
rect 13688 12968 13694 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 13688 12940 13829 12968
rect 13688 12928 13694 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 15654 12968 15660 12980
rect 15615 12940 15660 12968
rect 13817 12931 13875 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16574 12968 16580 12980
rect 16535 12940 16580 12968
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 7926 12900 7932 12912
rect 3936 12872 5120 12900
rect 7852 12872 7932 12900
rect 3936 12860 3942 12872
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 3970 12764 3976 12776
rect 3931 12736 3976 12764
rect 3970 12724 3976 12736
rect 4028 12764 4034 12776
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4028 12736 4353 12764
rect 4028 12724 4034 12736
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 4341 12727 4399 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7098 12773 7104 12776
rect 7092 12764 7104 12773
rect 7059 12736 7104 12764
rect 7092 12727 7104 12736
rect 7156 12764 7162 12776
rect 7852 12764 7880 12872
rect 7926 12860 7932 12872
rect 7984 12860 7990 12912
rect 9677 12903 9735 12909
rect 9677 12869 9689 12903
rect 9723 12900 9735 12903
rect 9950 12900 9956 12912
rect 9723 12872 9956 12900
rect 9723 12869 9735 12872
rect 9677 12863 9735 12869
rect 9950 12860 9956 12872
rect 10008 12900 10014 12912
rect 10597 12903 10655 12909
rect 10008 12872 10364 12900
rect 10008 12860 10014 12872
rect 10336 12841 10364 12872
rect 10597 12869 10609 12903
rect 10643 12900 10655 12903
rect 15562 12900 15568 12912
rect 10643 12872 11928 12900
rect 15475 12872 15568 12900
rect 10643 12869 10655 12872
rect 10597 12863 10655 12869
rect 10321 12835 10379 12841
rect 7156 12736 7880 12764
rect 7944 12804 8432 12832
rect 7098 12724 7104 12727
rect 7156 12724 7162 12736
rect 3881 12699 3939 12705
rect 3881 12696 3893 12699
rect 3804 12668 3893 12696
rect 3881 12665 3893 12668
rect 3927 12665 3939 12699
rect 3881 12659 3939 12665
rect 6086 12656 6092 12708
rect 6144 12696 6150 12708
rect 7944 12696 7972 12804
rect 8202 12764 8208 12776
rect 6144 12668 7972 12696
rect 8036 12736 8208 12764
rect 6144 12656 6150 12668
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2777 12631 2835 12637
rect 2777 12628 2789 12631
rect 2648 12600 2789 12628
rect 2648 12588 2654 12600
rect 2777 12597 2789 12600
rect 2823 12597 2835 12631
rect 2777 12591 2835 12597
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 8036 12628 8064 12736
rect 8202 12724 8208 12736
rect 8260 12764 8266 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 8260 12736 8309 12764
rect 8260 12724 8266 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8404 12764 8432 12804
rect 10321 12801 10333 12835
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11900 12841 11928 12872
rect 15562 12860 15568 12872
rect 15620 12900 15626 12912
rect 15838 12900 15844 12912
rect 15620 12872 15844 12900
rect 15620 12860 15626 12872
rect 15838 12860 15844 12872
rect 15896 12860 15902 12912
rect 11149 12835 11207 12841
rect 11149 12832 11161 12835
rect 10836 12804 11161 12832
rect 10836 12792 10842 12804
rect 11149 12801 11161 12804
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12801 11943 12835
rect 12066 12832 12072 12844
rect 11979 12804 12072 12832
rect 11885 12795 11943 12801
rect 12066 12792 12072 12804
rect 12124 12832 12130 12844
rect 12124 12804 12572 12832
rect 12124 12792 12130 12804
rect 12544 12776 12572 12804
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 13998 12832 14004 12844
rect 13872 12804 14004 12832
rect 13872 12792 13878 12804
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 15344 12804 16221 12832
rect 15344 12792 15350 12804
rect 16209 12801 16221 12804
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 10686 12764 10692 12776
rect 8404 12736 10692 12764
rect 8297 12727 8355 12733
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 10962 12764 10968 12776
rect 10923 12736 10968 12764
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 11296 12736 12265 12764
rect 11296 12724 11302 12736
rect 12253 12733 12265 12736
rect 12299 12764 12311 12767
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 12299 12736 12449 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 12710 12773 12716 12776
rect 12704 12764 12716 12773
rect 12671 12736 12716 12764
rect 12704 12727 12716 12736
rect 12768 12764 12774 12776
rect 13262 12764 13268 12776
rect 12768 12736 13268 12764
rect 12710 12724 12716 12727
rect 12768 12724 12774 12736
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13722 12724 13728 12776
rect 13780 12764 13786 12776
rect 14182 12764 14188 12776
rect 13780 12736 14188 12764
rect 13780 12724 13786 12736
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14452 12767 14510 12773
rect 14452 12733 14464 12767
rect 14498 12764 14510 12767
rect 14734 12764 14740 12776
rect 14498 12736 14740 12764
rect 14498 12733 14510 12736
rect 14452 12727 14510 12733
rect 14734 12724 14740 12736
rect 14792 12764 14798 12776
rect 15304 12764 15332 12792
rect 14792 12736 15332 12764
rect 14792 12724 14798 12736
rect 15378 12724 15384 12776
rect 15436 12764 15442 12776
rect 16025 12767 16083 12773
rect 16025 12764 16037 12767
rect 15436 12736 16037 12764
rect 15436 12724 15442 12736
rect 16025 12733 16037 12736
rect 16071 12764 16083 12767
rect 16574 12764 16580 12776
rect 16071 12736 16580 12764
rect 16071 12733 16083 12736
rect 16025 12727 16083 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 8542 12699 8600 12705
rect 8542 12696 8554 12699
rect 8220 12668 8554 12696
rect 8220 12640 8248 12668
rect 8542 12665 8554 12668
rect 8588 12665 8600 12699
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 8542 12659 8600 12665
rect 9784 12668 11069 12696
rect 8202 12628 8208 12640
rect 6880 12600 8064 12628
rect 8115 12600 8208 12628
rect 6880 12588 6886 12600
rect 8202 12588 8208 12600
rect 8260 12588 8266 12640
rect 9784 12637 9812 12668
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11606 12696 11612 12708
rect 11057 12659 11115 12665
rect 11440 12668 11612 12696
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12597 9827 12631
rect 9769 12591 9827 12597
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10042 12628 10048 12640
rect 9916 12600 10048 12628
rect 9916 12588 9922 12600
rect 10042 12588 10048 12600
rect 10100 12628 10106 12640
rect 10137 12631 10195 12637
rect 10137 12628 10149 12631
rect 10100 12600 10149 12628
rect 10100 12588 10106 12600
rect 10137 12597 10149 12600
rect 10183 12597 10195 12631
rect 10137 12591 10195 12597
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 11440 12637 11468 12668
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 11425 12631 11483 12637
rect 10284 12600 10329 12628
rect 10284 12588 10290 12600
rect 11425 12597 11437 12631
rect 11471 12597 11483 12631
rect 11425 12591 11483 12597
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11756 12600 11805 12628
rect 11756 12588 11762 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 11793 12591 11851 12597
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 13722 12628 13728 12640
rect 12299 12600 13728 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 16117 12631 16175 12637
rect 16117 12597 16129 12631
rect 16163 12628 16175 12631
rect 16298 12628 16304 12640
rect 16163 12600 16304 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 3421 12427 3479 12433
rect 3421 12393 3433 12427
rect 3467 12424 3479 12427
rect 3510 12424 3516 12436
rect 3467 12396 3516 12424
rect 3467 12393 3479 12396
rect 3421 12387 3479 12393
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 4246 12424 4252 12436
rect 3660 12396 4252 12424
rect 3660 12384 3666 12396
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 6822 12424 6828 12436
rect 5644 12396 6828 12424
rect 5644 12356 5672 12396
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 7340 12396 7573 12424
rect 7340 12384 7346 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 7561 12387 7619 12393
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 10226 12424 10232 12436
rect 9539 12396 10232 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 11057 12427 11115 12433
rect 11057 12424 11069 12427
rect 10836 12396 11069 12424
rect 10836 12384 10842 12396
rect 11057 12393 11069 12396
rect 11103 12424 11115 12427
rect 11422 12424 11428 12436
rect 11103 12396 11428 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 12986 12424 12992 12436
rect 12667 12396 12992 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 15252 12396 15301 12424
rect 15252 12384 15258 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15746 12424 15752 12436
rect 15707 12396 15752 12424
rect 15289 12387 15347 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 5896 12359 5954 12365
rect 5896 12356 5908 12359
rect 2056 12328 5672 12356
rect 2056 12300 2084 12328
rect 2038 12288 2044 12300
rect 1999 12260 2044 12288
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2308 12291 2366 12297
rect 2308 12257 2320 12291
rect 2354 12288 2366 12291
rect 3050 12288 3056 12300
rect 2354 12260 3056 12288
rect 2354 12257 2366 12260
rect 2308 12251 2366 12257
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 4172 12297 4200 12328
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 4246 12248 4252 12300
rect 4304 12288 4310 12300
rect 5644 12297 5672 12328
rect 5736 12328 5908 12356
rect 4413 12291 4471 12297
rect 4413 12288 4425 12291
rect 4304 12260 4425 12288
rect 4304 12248 4310 12260
rect 4413 12257 4425 12260
rect 4459 12257 4471 12291
rect 4413 12251 4471 12257
rect 5629 12291 5687 12297
rect 5629 12257 5641 12291
rect 5675 12257 5687 12291
rect 5629 12251 5687 12257
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 5736 12220 5764 12328
rect 5896 12325 5908 12328
rect 5942 12356 5954 12359
rect 7190 12356 7196 12368
rect 5942 12328 7196 12356
rect 5942 12325 5954 12328
rect 5896 12319 5954 12325
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 9309 12359 9367 12365
rect 9309 12325 9321 12359
rect 9355 12356 9367 12359
rect 9766 12356 9772 12368
rect 9355 12328 9772 12356
rect 9355 12325 9367 12328
rect 9309 12319 9367 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9950 12365 9956 12368
rect 9944 12356 9956 12365
rect 9911 12328 9956 12356
rect 9944 12319 9956 12328
rect 9950 12316 9956 12319
rect 10008 12316 10014 12368
rect 13992 12359 14050 12365
rect 13992 12325 14004 12359
rect 14038 12356 14050 12359
rect 15562 12356 15568 12368
rect 14038 12328 15568 12356
rect 14038 12325 14050 12328
rect 13992 12319 14050 12325
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 6236 12260 7481 12288
rect 6236 12248 6242 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 9490 12288 9496 12300
rect 8619 12260 9496 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 9490 12248 9496 12260
rect 9548 12248 9554 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 11146 12288 11152 12300
rect 9723 12260 11152 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11422 12297 11428 12300
rect 11416 12288 11428 12297
rect 11335 12260 11428 12288
rect 11416 12251 11428 12260
rect 11480 12288 11486 12300
rect 12250 12288 12256 12300
rect 11480 12260 12256 12288
rect 11422 12248 11428 12251
rect 11480 12248 11486 12260
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 12986 12288 12992 12300
rect 12947 12260 12992 12288
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 13722 12288 13728 12300
rect 13683 12260 13728 12288
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14274 12248 14280 12300
rect 14332 12288 14338 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14332 12260 15669 12288
rect 14332 12248 14338 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 5316 12192 5764 12220
rect 7745 12223 7803 12229
rect 5316 12180 5322 12192
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8202 12220 8208 12232
rect 7791 12192 8208 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12768 12192 13093 12220
rect 12768 12180 12774 12192
rect 13081 12189 13093 12192
rect 13127 12189 13139 12223
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 13081 12183 13139 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15120 12192 15853 12220
rect 15120 12161 15148 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 15105 12155 15163 12161
rect 6564 12124 9168 12152
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 6564 12084 6592 12124
rect 7006 12084 7012 12096
rect 5132 12056 6592 12084
rect 6967 12056 7012 12084
rect 5132 12044 5138 12056
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7156 12056 7201 12084
rect 7156 12044 7162 12056
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 8757 12087 8815 12093
rect 8757 12084 8769 12087
rect 8720 12056 8769 12084
rect 8720 12044 8726 12056
rect 8757 12053 8769 12056
rect 8803 12084 8815 12087
rect 8846 12084 8852 12096
rect 8803 12056 8852 12084
rect 8803 12053 8815 12056
rect 8757 12047 8815 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 9140 12084 9168 12124
rect 15105 12121 15117 12155
rect 15151 12152 15163 12155
rect 15194 12152 15200 12164
rect 15151 12124 15200 12152
rect 15151 12121 15163 12124
rect 15105 12115 15163 12121
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 10594 12084 10600 12096
rect 9140 12056 10600 12084
rect 10594 12044 10600 12056
rect 10652 12044 10658 12096
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12066 12084 12072 12096
rect 11848 12056 12072 12084
rect 11848 12044 11854 12056
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 16209 12087 16267 12093
rect 16209 12053 16221 12087
rect 16255 12084 16267 12087
rect 16298 12084 16304 12096
rect 16255 12056 16304 12084
rect 16255 12053 16267 12056
rect 16209 12047 16267 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2314 11880 2320 11892
rect 1627 11852 2320 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2314 11840 2320 11852
rect 2372 11840 2378 11892
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3605 11883 3663 11889
rect 3605 11880 3617 11883
rect 3292 11852 3617 11880
rect 3292 11840 3298 11852
rect 3605 11849 3617 11852
rect 3651 11849 3663 11883
rect 3605 11843 3663 11849
rect 4985 11883 5043 11889
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 6178 11880 6184 11892
rect 5031 11852 6184 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7432 11852 8033 11880
rect 7432 11840 7438 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 8021 11843 8079 11849
rect 8849 11883 8907 11889
rect 8849 11849 8861 11883
rect 8895 11880 8907 11883
rect 9950 11880 9956 11892
rect 8895 11852 9956 11880
rect 8895 11849 8907 11852
rect 8849 11843 8907 11849
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 11698 11880 11704 11892
rect 10183 11852 11704 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 13078 11880 13084 11892
rect 12483 11852 13084 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 8386 11812 8392 11824
rect 4028 11784 8392 11812
rect 4028 11772 4034 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 9030 11772 9036 11824
rect 9088 11812 9094 11824
rect 10965 11815 11023 11821
rect 9088 11784 10640 11812
rect 9088 11772 9094 11784
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 3050 11704 3056 11716
rect 3108 11744 3114 11756
rect 4062 11744 4068 11756
rect 3108 11716 4068 11744
rect 3108 11704 3114 11716
rect 4062 11704 4068 11716
rect 4120 11744 4126 11756
rect 4157 11747 4215 11753
rect 4157 11744 4169 11747
rect 4120 11716 4169 11744
rect 4120 11704 4126 11716
rect 4157 11713 4169 11716
rect 4203 11713 4215 11747
rect 4157 11707 4215 11713
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4525 11747 4583 11753
rect 4525 11744 4537 11747
rect 4304 11716 4537 11744
rect 4304 11704 4310 11716
rect 4525 11713 4537 11716
rect 4571 11744 4583 11747
rect 5074 11744 5080 11756
rect 4571 11716 5080 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 7006 11744 7012 11756
rect 5675 11716 7012 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8662 11744 8668 11756
rect 8623 11716 8668 11744
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 8904 11716 9321 11744
rect 8904 11704 8910 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 9493 11747 9551 11753
rect 9493 11713 9505 11747
rect 9539 11744 9551 11747
rect 9582 11744 9588 11756
rect 9539 11716 9588 11744
rect 9539 11713 9551 11716
rect 9493 11707 9551 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 10612 11753 10640 11784
rect 10965 11781 10977 11815
rect 11011 11812 11023 11815
rect 11146 11812 11152 11824
rect 11011 11784 11152 11812
rect 11011 11781 11023 11784
rect 10965 11775 11023 11781
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 11900 11812 11928 11840
rect 11440 11784 11928 11812
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11713 10655 11747
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10597 11707 10655 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11440 11753 11468 11784
rect 13722 11772 13728 11824
rect 13780 11812 13786 11824
rect 13780 11784 14964 11812
rect 13780 11772 13786 11784
rect 11425 11747 11483 11753
rect 11425 11713 11437 11747
rect 11471 11713 11483 11747
rect 11425 11707 11483 11713
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11744 11667 11747
rect 11790 11744 11796 11756
rect 11655 11716 11796 11744
rect 11655 11713 11667 11716
rect 11609 11707 11667 11713
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12584 11716 13001 11744
rect 12584 11704 12590 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 14734 11744 14740 11756
rect 14695 11716 14740 11744
rect 12989 11707 13047 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 14936 11753 14964 11784
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2777 11679 2835 11685
rect 2777 11676 2789 11679
rect 2372 11648 2789 11676
rect 2372 11636 2378 11648
rect 2777 11645 2789 11648
rect 2823 11676 2835 11679
rect 3418 11676 3424 11688
rect 2823 11648 3424 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3878 11636 3884 11688
rect 3936 11676 3942 11688
rect 6822 11676 6828 11688
rect 3936 11648 6828 11676
rect 3936 11636 3942 11648
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 12894 11676 12900 11688
rect 7156 11648 12900 11676
rect 7156 11636 7162 11648
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 14001 11679 14059 11685
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14090 11676 14096 11688
rect 14047 11648 14096 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14090 11636 14096 11648
rect 14148 11676 14154 11688
rect 15194 11685 15200 11688
rect 15188 11676 15200 11685
rect 14148 11648 14412 11676
rect 15155 11648 15200 11676
rect 14148 11636 14154 11648
rect 1486 11608 1492 11620
rect 1399 11580 1492 11608
rect 1486 11568 1492 11580
rect 1544 11608 1550 11620
rect 2869 11611 2927 11617
rect 2869 11608 2881 11611
rect 1544 11580 2881 11608
rect 1544 11568 1550 11580
rect 2869 11577 2881 11580
rect 2915 11608 2927 11611
rect 2958 11608 2964 11620
rect 2915 11580 2964 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 3513 11611 3571 11617
rect 3513 11577 3525 11611
rect 3559 11608 3571 11611
rect 3973 11611 4031 11617
rect 3973 11608 3985 11611
rect 3559 11580 3985 11608
rect 3559 11577 3571 11580
rect 3513 11571 3571 11577
rect 3973 11577 3985 11580
rect 4019 11608 4031 11611
rect 4890 11608 4896 11620
rect 4019 11580 4896 11608
rect 4019 11577 4031 11580
rect 3973 11571 4031 11577
rect 4890 11568 4896 11580
rect 4948 11608 4954 11620
rect 5074 11608 5080 11620
rect 4948 11580 5080 11608
rect 4948 11568 4954 11580
rect 5074 11568 5080 11580
rect 5132 11568 5138 11620
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 7374 11608 7380 11620
rect 6788 11580 7380 11608
rect 6788 11568 6794 11580
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 8481 11611 8539 11617
rect 8481 11577 8493 11611
rect 8527 11608 8539 11611
rect 9674 11608 9680 11620
rect 8527 11580 9680 11608
rect 8527 11577 8539 11580
rect 8481 11571 8539 11577
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 9861 11611 9919 11617
rect 9861 11577 9873 11611
rect 9907 11608 9919 11611
rect 10870 11608 10876 11620
rect 9907 11580 10876 11608
rect 9907 11577 9919 11580
rect 9861 11571 9919 11577
rect 10870 11568 10876 11580
rect 10928 11608 10934 11620
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 10928 11580 11345 11608
rect 10928 11568 10934 11580
rect 11333 11577 11345 11580
rect 11379 11577 11391 11611
rect 14182 11608 14188 11620
rect 11333 11571 11391 11577
rect 11624 11580 14188 11608
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 2087 11512 2421 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4246 11540 4252 11552
rect 4111 11512 4252 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 5350 11540 5356 11552
rect 5311 11512 5356 11540
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5500 11512 5545 11540
rect 5500 11500 5506 11512
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7064 11512 8401 11540
rect 7064 11500 7070 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 9217 11543 9275 11549
rect 9217 11509 9229 11543
rect 9263 11540 9275 11543
rect 9490 11540 9496 11552
rect 9263 11512 9496 11540
rect 9263 11509 9275 11512
rect 9217 11503 9275 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 10042 11540 10048 11552
rect 9955 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11540 10106 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10100 11512 10517 11540
rect 10100 11500 10106 11512
rect 10505 11509 10517 11512
rect 10551 11540 10563 11543
rect 11624 11540 11652 11580
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 14384 11552 14412 11648
rect 15188 11639 15200 11648
rect 15194 11636 15200 11639
rect 15252 11636 15258 11688
rect 14461 11611 14519 11617
rect 14461 11577 14473 11611
rect 14507 11608 14519 11611
rect 15286 11608 15292 11620
rect 14507 11580 15292 11608
rect 14507 11577 14519 11580
rect 14461 11571 14519 11577
rect 15286 11568 15292 11580
rect 15344 11568 15350 11620
rect 10551 11512 11652 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 11756 11512 12817 11540
rect 11756 11500 11762 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 14090 11540 14096 11552
rect 12952 11512 12997 11540
rect 14051 11512 14096 11540
rect 12952 11500 12958 11512
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14553 11543 14611 11549
rect 14553 11540 14565 11543
rect 14424 11512 14565 11540
rect 14424 11500 14430 11512
rect 14553 11509 14565 11512
rect 14599 11509 14611 11543
rect 14553 11503 14611 11509
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 15252 11512 16313 11540
rect 15252 11500 15258 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1946 11296 1952 11348
rect 2004 11336 2010 11348
rect 2317 11339 2375 11345
rect 2317 11336 2329 11339
rect 2004 11308 2329 11336
rect 2004 11296 2010 11308
rect 2317 11305 2329 11308
rect 2363 11305 2375 11339
rect 2317 11299 2375 11305
rect 4709 11339 4767 11345
rect 4709 11305 4721 11339
rect 4755 11336 4767 11339
rect 5350 11336 5356 11348
rect 4755 11308 5356 11336
rect 4755 11305 4767 11308
rect 4709 11299 4767 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 6822 11296 6828 11348
rect 6880 11336 6886 11348
rect 6880 11308 8616 11336
rect 6880 11296 6886 11308
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11268 1915 11271
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 1903 11240 2789 11268
rect 1903 11237 1915 11240
rect 1857 11231 1915 11237
rect 2777 11237 2789 11240
rect 2823 11268 2835 11271
rect 2958 11268 2964 11280
rect 2823 11240 2964 11268
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 2958 11228 2964 11240
rect 3016 11268 3022 11280
rect 3602 11268 3608 11280
rect 3016 11240 3608 11268
rect 3016 11228 3022 11240
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 7282 11268 7288 11280
rect 4120 11240 7288 11268
rect 4120 11228 4126 11240
rect 7282 11228 7288 11240
rect 7340 11228 7346 11280
rect 2133 11203 2191 11209
rect 2133 11169 2145 11203
rect 2179 11200 2191 11203
rect 2314 11200 2320 11212
rect 2179 11172 2320 11200
rect 2179 11169 2191 11172
rect 2133 11163 2191 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 6730 11209 6736 11212
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 2731 11172 3157 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 3145 11169 3157 11172
rect 3191 11169 3203 11203
rect 3145 11163 3203 11169
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5537 11203 5595 11209
rect 5537 11200 5549 11203
rect 5123 11172 5549 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5537 11169 5549 11172
rect 5583 11169 5595 11203
rect 6724 11200 6736 11209
rect 6691 11172 6736 11200
rect 5537 11163 5595 11169
rect 6724 11163 6736 11172
rect 6730 11160 6736 11163
rect 6788 11160 6794 11212
rect 8202 11209 8208 11212
rect 8196 11200 8208 11209
rect 7852 11172 8208 11200
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3050 11132 3056 11144
rect 3007 11104 3056 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3050 11092 3056 11104
rect 3108 11132 3114 11144
rect 3694 11132 3700 11144
rect 3108 11104 3700 11132
rect 3108 11092 3114 11104
rect 3694 11092 3700 11104
rect 3752 11092 3758 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11101 5227 11135
rect 5169 11095 5227 11101
rect 4617 11067 4675 11073
rect 4617 11033 4629 11067
rect 4663 11064 4675 11067
rect 4982 11064 4988 11076
rect 4663 11036 4988 11064
rect 4663 11033 4675 11036
rect 4617 11027 4675 11033
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4632 10996 4660 11027
rect 4982 11024 4988 11036
rect 5040 11064 5046 11076
rect 5184 11064 5212 11095
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 6454 11132 6460 11144
rect 5316 11104 5361 11132
rect 6415 11104 6460 11132
rect 5316 11092 5322 11104
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 7852 11073 7880 11172
rect 8196 11163 8208 11172
rect 8202 11160 8208 11163
rect 8260 11160 8266 11212
rect 8588 11200 8616 11308
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8720 11308 9321 11336
rect 8720 11296 8726 11308
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 9309 11299 9367 11305
rect 9600 11308 10977 11336
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 9600 11268 9628 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 11701 11339 11759 11345
rect 11701 11305 11713 11339
rect 11747 11336 11759 11339
rect 12894 11336 12900 11348
rect 11747 11308 12900 11336
rect 11747 11305 11759 11308
rect 11701 11299 11759 11305
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13265 11339 13323 11345
rect 13265 11305 13277 11339
rect 13311 11336 13323 11339
rect 13906 11336 13912 11348
rect 13311 11308 13912 11336
rect 13311 11305 13323 11308
rect 13265 11299 13323 11305
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 14148 11308 14657 11336
rect 14148 11296 14154 11308
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 14645 11299 14703 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 9272 11240 9628 11268
rect 9677 11271 9735 11277
rect 9272 11228 9278 11240
rect 9677 11237 9689 11271
rect 9723 11268 9735 11271
rect 17218 11268 17224 11280
rect 9723 11240 17224 11268
rect 9723 11237 9735 11240
rect 9677 11231 9735 11237
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 11238 11200 11244 11212
rect 8588 11172 11244 11200
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 11900 11172 12081 11200
rect 11900 11144 11928 11172
rect 12069 11169 12081 11172
rect 12115 11169 12127 11203
rect 12069 11163 12127 11169
rect 12434 11160 12440 11212
rect 12492 11200 12498 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 12492 11172 13645 11200
rect 12492 11160 12498 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 17494 11200 17500 11212
rect 13633 11163 13691 11169
rect 14108 11172 17500 11200
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11132 11667 11135
rect 11882 11132 11888 11144
rect 11655 11104 11888 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 5040 11036 5212 11064
rect 7837 11067 7895 11073
rect 5040 11024 5046 11036
rect 7837 11033 7849 11067
rect 7883 11033 7895 11067
rect 7837 11027 7895 11033
rect 4028 10968 4660 10996
rect 4028 10956 4034 10968
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 7944 10996 7972 11095
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12161 11135 12219 11141
rect 12161 11132 12173 11135
rect 12032 11104 12173 11132
rect 12032 11092 12038 11104
rect 12161 11101 12173 11104
rect 12207 11101 12219 11135
rect 12161 11095 12219 11101
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 13722 11132 13728 11144
rect 12308 11104 12353 11132
rect 13683 11104 13728 11132
rect 12308 11092 12314 11104
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13906 11132 13912 11144
rect 13867 11104 13912 11132
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 9214 11064 9220 11076
rect 8996 11036 9220 11064
rect 8996 11024 9002 11036
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 9401 11067 9459 11073
rect 9401 11064 9413 11067
rect 9324 11036 9413 11064
rect 8294 10996 8300 11008
rect 6512 10968 8300 10996
rect 6512 10956 6518 10968
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 9324 10996 9352 11036
rect 9401 11033 9413 11036
rect 9447 11064 9459 11067
rect 10410 11064 10416 11076
rect 9447 11036 10416 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 10410 11024 10416 11036
rect 10468 11064 10474 11076
rect 14108 11064 14136 11172
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 14734 11132 14740 11144
rect 14695 11104 14740 11132
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11132 14979 11135
rect 15562 11132 15568 11144
rect 14967 11104 15568 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 14274 11064 14280 11076
rect 10468 11036 14136 11064
rect 14235 11036 14280 11064
rect 10468 11024 10474 11036
rect 14274 11024 14280 11036
rect 14332 11024 14338 11076
rect 8628 10968 9352 10996
rect 8628 10956 8634 10968
rect 9490 10956 9496 11008
rect 9548 10996 9554 11008
rect 12618 10996 12624 11008
rect 9548 10968 12624 10996
rect 9548 10956 9554 10968
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 5077 10795 5135 10801
rect 1636 10764 3924 10792
rect 1636 10752 1642 10764
rect 3896 10668 3924 10764
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5442 10792 5448 10804
rect 5123 10764 5448 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 7006 10792 7012 10804
rect 5951 10764 7012 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 7006 10752 7012 10764
rect 7064 10752 7070 10804
rect 10873 10795 10931 10801
rect 7484 10764 9628 10792
rect 7098 10724 7104 10736
rect 4908 10696 7104 10724
rect 4908 10668 4936 10696
rect 7098 10684 7104 10696
rect 7156 10684 7162 10736
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 3936 10628 4721 10656
rect 3936 10616 3942 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4890 10656 4896 10668
rect 4803 10628 4896 10656
rect 4709 10619 4767 10625
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5316 10628 5641 10656
rect 5316 10616 5322 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 1765 10591 1823 10597
rect 1765 10557 1777 10591
rect 1811 10588 1823 10591
rect 1854 10588 1860 10600
rect 1811 10560 1860 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 2032 10591 2090 10597
rect 2032 10557 2044 10591
rect 2078 10588 2090 10591
rect 2590 10588 2596 10600
rect 2078 10560 2596 10588
rect 2078 10557 2090 10560
rect 2032 10551 2090 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 4157 10591 4215 10597
rect 4157 10588 4169 10591
rect 3660 10560 4169 10588
rect 3660 10548 3666 10560
rect 4157 10557 4169 10560
rect 4203 10588 4215 10591
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 4203 10560 5549 10588
rect 4203 10557 4215 10560
rect 4157 10551 4215 10557
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 6564 10588 6592 10619
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 7484 10665 7512 10764
rect 9600 10736 9628 10764
rect 10873 10761 10885 10795
rect 10919 10792 10931 10795
rect 11698 10792 11704 10804
rect 10919 10764 11704 10792
rect 10919 10761 10931 10764
rect 10873 10755 10931 10761
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 13722 10792 13728 10804
rect 12759 10764 13728 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 14792 10764 15025 10792
rect 14792 10752 14798 10764
rect 15013 10761 15025 10764
rect 15059 10761 15071 10795
rect 15013 10755 15071 10761
rect 9582 10684 9588 10736
rect 9640 10724 9646 10736
rect 9640 10696 13492 10724
rect 9640 10684 9646 10696
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 6788 10628 7481 10656
rect 6788 10616 6794 10628
rect 7469 10625 7481 10628
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9456 10628 9873 10656
rect 9456 10616 9462 10628
rect 9861 10625 9873 10628
rect 9907 10656 9919 10659
rect 10594 10656 10600 10668
rect 9907 10628 10600 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 10594 10616 10600 10628
rect 10652 10616 10658 10668
rect 10704 10665 10732 10696
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 12250 10656 12256 10668
rect 11563 10628 12256 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 12250 10616 12256 10628
rect 12308 10616 12314 10668
rect 13262 10656 13268 10668
rect 13223 10628 13268 10656
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 6564 10560 8248 10588
rect 5537 10551 5595 10557
rect 8220 10532 8248 10560
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 10318 10588 10324 10600
rect 8352 10560 8397 10588
rect 8496 10560 10324 10588
rect 8352 10548 8358 10560
rect 3973 10523 4031 10529
rect 3973 10489 3985 10523
rect 4019 10520 4031 10523
rect 4338 10520 4344 10532
rect 4019 10492 4344 10520
rect 4019 10489 4031 10492
rect 3973 10483 4031 10489
rect 4338 10480 4344 10492
rect 4396 10520 4402 10532
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 4396 10492 5457 10520
rect 4396 10480 4402 10492
rect 5445 10489 5457 10492
rect 5491 10489 5503 10523
rect 5445 10483 5503 10489
rect 6273 10523 6331 10529
rect 6273 10489 6285 10523
rect 6319 10520 6331 10523
rect 7193 10523 7251 10529
rect 6319 10492 6868 10520
rect 6319 10489 6331 10492
rect 6273 10483 6331 10489
rect 1486 10412 1492 10464
rect 1544 10452 1550 10464
rect 2314 10452 2320 10464
rect 1544 10424 2320 10452
rect 1544 10412 1550 10424
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3789 10455 3847 10461
rect 3789 10421 3801 10455
rect 3835 10452 3847 10455
rect 3878 10452 3884 10464
rect 3835 10424 3884 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 4246 10452 4252 10464
rect 4207 10424 4252 10452
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 4614 10452 4620 10464
rect 4575 10424 4620 10452
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 6840 10461 6868 10492
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 7653 10523 7711 10529
rect 7653 10520 7665 10523
rect 7239 10492 7665 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 7653 10489 7665 10492
rect 7699 10489 7711 10523
rect 7653 10483 7711 10489
rect 8202 10480 8208 10532
rect 8260 10520 8266 10532
rect 8496 10520 8524 10560
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10413 10591 10471 10597
rect 10413 10557 10425 10591
rect 10459 10588 10471 10591
rect 10778 10588 10784 10600
rect 10459 10560 10784 10588
rect 10459 10557 10471 10560
rect 10413 10551 10471 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 11204 10560 13185 10588
rect 11204 10548 11210 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 8260 10492 8524 10520
rect 8564 10523 8622 10529
rect 8260 10480 8266 10492
rect 8564 10489 8576 10523
rect 8610 10520 8622 10523
rect 8662 10520 8668 10532
rect 8610 10492 8668 10520
rect 8610 10489 8622 10492
rect 8564 10483 8622 10489
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 10870 10520 10876 10532
rect 9088 10492 10876 10520
rect 9088 10480 9094 10492
rect 10870 10480 10876 10492
rect 10928 10480 10934 10532
rect 11241 10523 11299 10529
rect 11241 10489 11253 10523
rect 11287 10520 11299 10523
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 11287 10492 12081 10520
rect 11287 10489 11299 10492
rect 11241 10483 11299 10489
rect 12069 10489 12081 10492
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 6825 10455 6883 10461
rect 6420 10424 6465 10452
rect 6420 10412 6426 10424
rect 6825 10421 6837 10455
rect 6871 10421 6883 10455
rect 7282 10452 7288 10464
rect 7243 10424 7288 10452
rect 6825 10415 6883 10421
rect 7282 10412 7288 10424
rect 7340 10452 7346 10464
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7340 10424 7941 10452
rect 7340 10412 7346 10424
rect 7929 10421 7941 10424
rect 7975 10421 7987 10455
rect 7929 10415 7987 10421
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9766 10452 9772 10464
rect 9723 10424 9772 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10410 10412 10416 10464
rect 10468 10452 10474 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10468 10424 10517 10452
rect 10468 10412 10474 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 10594 10412 10600 10464
rect 10652 10452 10658 10464
rect 11330 10452 11336 10464
rect 10652 10424 11336 10452
rect 10652 10412 10658 10424
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 11974 10452 11980 10464
rect 11839 10424 11980 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 13081 10455 13139 10461
rect 13081 10452 13093 10455
rect 12952 10424 13093 10452
rect 12952 10412 12958 10424
rect 13081 10421 13093 10424
rect 13127 10421 13139 10455
rect 13464 10452 13492 10696
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 15565 10659 15623 10665
rect 15565 10656 15577 10659
rect 14884 10628 15577 10656
rect 14884 10616 14890 10628
rect 15565 10625 15577 10628
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 13538 10548 13544 10600
rect 13596 10588 13602 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 13596 10560 13641 10588
rect 14660 10560 15485 10588
rect 13596 10548 13602 10560
rect 14660 10532 14688 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 13808 10523 13866 10529
rect 13808 10489 13820 10523
rect 13854 10520 13866 10523
rect 13906 10520 13912 10532
rect 13854 10492 13912 10520
rect 13854 10489 13866 10492
rect 13808 10483 13866 10489
rect 13906 10480 13912 10492
rect 13964 10520 13970 10532
rect 14366 10520 14372 10532
rect 13964 10492 14372 10520
rect 13964 10480 13970 10492
rect 14366 10480 14372 10492
rect 14424 10480 14430 10532
rect 14642 10480 14648 10532
rect 14700 10480 14706 10532
rect 14734 10480 14740 10532
rect 14792 10520 14798 10532
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 14792 10492 15393 10520
rect 14792 10480 14798 10492
rect 15381 10489 15393 10492
rect 15427 10489 15439 10523
rect 15381 10483 15439 10489
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 13464 10424 14933 10452
rect 13081 10415 13139 10421
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 3694 10248 3700 10260
rect 3655 10220 3700 10248
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 4672 10220 5549 10248
rect 4672 10208 4678 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 5537 10211 5595 10217
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 9398 10248 9404 10260
rect 6748 10220 9404 10248
rect 1949 10183 2007 10189
rect 1949 10149 1961 10183
rect 1995 10180 2007 10183
rect 2498 10180 2504 10192
rect 1995 10152 2504 10180
rect 1995 10149 2007 10152
rect 1949 10143 2007 10149
rect 2498 10140 2504 10152
rect 2556 10140 2562 10192
rect 4332 10183 4390 10189
rect 4332 10149 4344 10183
rect 4378 10180 4390 10183
rect 4890 10180 4896 10192
rect 4378 10152 4896 10180
rect 4378 10149 4390 10152
rect 4332 10143 4390 10149
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 6748 10180 6776 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9674 10248 9680 10260
rect 9635 10220 9680 10248
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10870 10248 10876 10260
rect 10831 10220 10876 10248
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 12250 10248 12256 10260
rect 11388 10220 12256 10248
rect 11388 10208 11394 10220
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12897 10251 12955 10257
rect 12897 10217 12909 10251
rect 12943 10217 12955 10251
rect 14366 10248 14372 10260
rect 14327 10220 14372 10248
rect 12897 10211 12955 10217
rect 6288 10152 6776 10180
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 1762 10112 1768 10124
rect 1719 10084 1768 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 1762 10072 1768 10084
rect 1820 10072 1826 10124
rect 2584 10115 2642 10121
rect 2584 10081 2596 10115
rect 2630 10112 2642 10115
rect 3050 10112 3056 10124
rect 2630 10084 3056 10112
rect 2630 10081 2642 10084
rect 2584 10075 2642 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 3970 10072 3976 10124
rect 4028 10112 4034 10124
rect 6288 10112 6316 10152
rect 6822 10140 6828 10192
rect 6880 10140 6886 10192
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 8481 10183 8539 10189
rect 7156 10152 7972 10180
rect 7156 10140 7162 10152
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 4028 10084 6316 10112
rect 6380 10084 6745 10112
rect 4028 10072 4034 10084
rect 6380 10056 6408 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 6840 10112 6868 10140
rect 7653 10115 7711 10121
rect 6840 10084 6960 10112
rect 6733 10075 6791 10081
rect 1854 10004 1860 10056
rect 1912 10044 1918 10056
rect 2317 10047 2375 10053
rect 2317 10044 2329 10047
rect 1912 10016 2329 10044
rect 1912 10004 1918 10016
rect 2317 10013 2329 10016
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6362 10044 6368 10056
rect 6135 10016 6368 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 2332 9908 2360 10007
rect 4080 9908 4108 10007
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 6932 10053 6960 10084
rect 7653 10081 7665 10115
rect 7699 10112 7711 10115
rect 7699 10084 7880 10112
rect 7699 10081 7711 10084
rect 7653 10075 7711 10081
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6696 10016 6837 10044
rect 6696 10004 6702 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 7742 10044 7748 10056
rect 7703 10016 7748 10044
rect 6917 10007 6975 10013
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 5626 9936 5632 9988
rect 5684 9976 5690 9988
rect 7285 9979 7343 9985
rect 7285 9976 7297 9979
rect 5684 9948 7297 9976
rect 5684 9936 5690 9948
rect 7285 9945 7297 9948
rect 7331 9945 7343 9979
rect 7852 9976 7880 10084
rect 7944 10053 7972 10152
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 9030 10180 9036 10192
rect 8527 10152 9036 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 9030 10140 9036 10152
rect 9088 10140 9094 10192
rect 9125 10183 9183 10189
rect 9125 10149 9137 10183
rect 9171 10180 9183 10183
rect 10226 10180 10232 10192
rect 9171 10152 10232 10180
rect 9171 10149 9183 10152
rect 9125 10143 9183 10149
rect 10226 10140 10232 10152
rect 10284 10140 10290 10192
rect 11790 10189 11796 10192
rect 11784 10180 11796 10189
rect 11751 10152 11796 10180
rect 11784 10143 11796 10152
rect 11790 10140 11796 10143
rect 11848 10140 11854 10192
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12342 10180 12348 10192
rect 11940 10152 12348 10180
rect 11940 10140 11946 10152
rect 12342 10140 12348 10152
rect 12400 10140 12406 10192
rect 12912 10180 12940 10211
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14642 10248 14648 10260
rect 14603 10220 14648 10248
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 14792 10220 14841 10248
rect 14792 10208 14798 10220
rect 14829 10217 14841 10220
rect 14875 10217 14887 10251
rect 14829 10211 14887 10217
rect 13262 10189 13268 10192
rect 13256 10180 13268 10189
rect 12912 10152 13268 10180
rect 13256 10143 13268 10152
rect 13262 10140 13268 10143
rect 13320 10140 13326 10192
rect 8665 10115 8723 10121
rect 8665 10081 8677 10115
rect 8711 10112 8723 10115
rect 9674 10112 9680 10124
rect 8711 10084 9680 10112
rect 8711 10081 8723 10084
rect 8665 10075 8723 10081
rect 9674 10072 9680 10084
rect 9732 10112 9738 10124
rect 9858 10112 9864 10124
rect 9732 10084 9864 10112
rect 9732 10072 9738 10084
rect 9858 10072 9864 10084
rect 9916 10072 9922 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 10008 10084 10149 10112
rect 10008 10072 10014 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 10836 10084 11437 10112
rect 10836 10072 10842 10084
rect 11425 10081 11437 10084
rect 11471 10112 11483 10115
rect 12158 10112 12164 10124
rect 11471 10084 12164 10112
rect 11471 10081 11483 10084
rect 11425 10075 11483 10081
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 13538 10112 13544 10124
rect 13035 10084 13544 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8202 10044 8208 10056
rect 7975 10016 8208 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9214 10044 9220 10056
rect 9175 10016 9220 10044
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 10042 10044 10048 10056
rect 9447 10016 10048 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 8754 9976 8760 9988
rect 7852 9948 8248 9976
rect 8715 9948 8760 9976
rect 7285 9939 7343 9945
rect 5442 9908 5448 9920
rect 2332 9880 4108 9908
rect 5403 9880 5448 9908
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 6273 9911 6331 9917
rect 6273 9877 6285 9911
rect 6319 9908 6331 9911
rect 6638 9908 6644 9920
rect 6319 9880 6644 9908
rect 6319 9877 6331 9880
rect 6273 9871 6331 9877
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 8220 9917 8248 9948
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 11072 9976 11100 10007
rect 9824 9948 11100 9976
rect 9824 9936 9830 9948
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 8846 9908 8852 9920
rect 8251 9880 8852 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 10505 9911 10563 9917
rect 10505 9908 10517 9911
rect 9916 9880 10517 9908
rect 9916 9868 9922 9880
rect 10505 9877 10517 9880
rect 10551 9877 10563 9911
rect 11532 9908 11560 10007
rect 12526 9908 12532 9920
rect 11532 9880 12532 9908
rect 10505 9871 10563 9877
rect 12526 9868 12532 9880
rect 12584 9908 12590 9920
rect 13004 9908 13032 10075
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 12584 9880 13032 9908
rect 12584 9868 12590 9880
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 8202 9704 8208 9716
rect 4120 9676 8064 9704
rect 8163 9676 8208 9704
rect 4120 9664 4126 9676
rect 3786 9596 3792 9648
rect 3844 9636 3850 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 3844 9608 3985 9636
rect 3844 9596 3850 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 3973 9599 4031 9605
rect 5350 9596 5356 9648
rect 5408 9636 5414 9648
rect 6822 9636 6828 9648
rect 5408 9608 6828 9636
rect 5408 9596 5414 9608
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 8036 9636 8064 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9490 9704 9496 9716
rect 8312 9676 9496 9704
rect 8312 9636 8340 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 10962 9704 10968 9716
rect 9732 9676 10968 9704
rect 9732 9664 9738 9676
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 11848 9676 12112 9704
rect 11848 9664 11854 9676
rect 8036 9608 8340 9636
rect 8478 9596 8484 9648
rect 8536 9596 8542 9648
rect 10137 9639 10195 9645
rect 10137 9605 10149 9639
rect 10183 9605 10195 9639
rect 10137 9599 10195 9605
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4212 9540 4537 9568
rect 4212 9528 4218 9540
rect 4525 9537 4537 9540
rect 4571 9568 4583 9571
rect 5442 9568 5448 9580
rect 4571 9540 5448 9568
rect 4571 9537 4583 9540
rect 4525 9531 4583 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 5718 9568 5724 9580
rect 5583 9540 5724 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 8496 9568 8524 9596
rect 8220 9540 8524 9568
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 1964 9432 1992 9463
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 4304 9472 4353 9500
rect 4304 9460 4310 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 5626 9500 5632 9512
rect 4479 9472 5632 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 5902 9500 5908 9512
rect 5863 9472 5908 9500
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 6454 9432 6460 9444
rect 1964 9404 4936 9432
rect 4908 9373 4936 9404
rect 5828 9404 6460 9432
rect 5828 9376 5856 9404
rect 6454 9392 6460 9404
rect 6512 9432 6518 9444
rect 6840 9432 6868 9463
rect 6512 9404 6868 9432
rect 7092 9435 7150 9441
rect 6512 9392 6518 9404
rect 7092 9401 7104 9435
rect 7138 9432 7150 9435
rect 7190 9432 7196 9444
rect 7138 9404 7196 9432
rect 7138 9401 7150 9404
rect 7092 9395 7150 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 8220 9432 8248 9540
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10152 9568 10180 9599
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10284 9608 10329 9636
rect 10284 9596 10290 9608
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11333 9639 11391 9645
rect 11333 9636 11345 9639
rect 11296 9608 11345 9636
rect 11296 9596 11302 9608
rect 11333 9605 11345 9608
rect 11379 9636 11391 9639
rect 11379 9608 12020 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 11992 9580 12020 9608
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10008 9540 10793 9568
rect 10008 9528 10014 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 11974 9568 11980 9580
rect 11887 9540 11980 9568
rect 10781 9531 10839 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12084 9577 12112 9676
rect 12894 9664 12900 9716
rect 12952 9704 12958 9716
rect 13633 9707 13691 9713
rect 13633 9704 13645 9707
rect 12952 9676 13645 9704
rect 12952 9664 12958 9676
rect 13633 9673 13645 9676
rect 13679 9673 13691 9707
rect 13633 9667 13691 9673
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 12537 9636
rect 12492 9596 12498 9608
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13354 9636 13360 9648
rect 13044 9608 13360 9636
rect 13044 9596 13050 9608
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 13081 9571 13139 9577
rect 12115 9540 13032 9568
rect 12115 9537 12127 9540
rect 12069 9531 12127 9537
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 9024 9503 9082 9509
rect 9024 9469 9036 9503
rect 9070 9500 9082 9503
rect 9766 9500 9772 9512
rect 9070 9472 9772 9500
rect 9070 9469 9082 9472
rect 9024 9463 9082 9469
rect 7576 9404 8248 9432
rect 8772 9432 8800 9463
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 11146 9460 11152 9512
rect 11204 9500 11210 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 11204 9472 12909 9500
rect 11204 9460 11210 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 13004 9500 13032 9540
rect 13081 9537 13093 9571
rect 13127 9568 13139 9571
rect 13262 9568 13268 9580
rect 13127 9540 13268 9568
rect 13127 9537 13139 9540
rect 13081 9531 13139 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 15102 9568 15108 9580
rect 14323 9540 15108 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14292 9500 14320 9531
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 13004 9472 14320 9500
rect 12897 9463 12955 9469
rect 8772 9404 9168 9432
rect 4893 9367 4951 9373
rect 4893 9333 4905 9367
rect 4939 9333 4951 9367
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 4893 9327 4951 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 5721 9367 5779 9373
rect 5408 9336 5453 9364
rect 5408 9324 5414 9336
rect 5721 9333 5733 9367
rect 5767 9364 5779 9367
rect 5810 9364 5816 9376
rect 5767 9336 5816 9364
rect 5767 9333 5779 9336
rect 5721 9327 5779 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 7576 9364 7604 9404
rect 6236 9336 7604 9364
rect 6236 9324 6242 9336
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8202 9364 8208 9376
rect 7708 9336 8208 9364
rect 7708 9324 7714 9336
rect 8202 9324 8208 9336
rect 8260 9364 8266 9376
rect 8297 9367 8355 9373
rect 8297 9364 8309 9367
rect 8260 9336 8309 9364
rect 8260 9324 8266 9336
rect 8297 9333 8309 9336
rect 8343 9333 8355 9367
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8297 9327 8355 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9140 9364 9168 9404
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 10689 9435 10747 9441
rect 10689 9432 10701 9435
rect 9456 9404 10701 9432
rect 9456 9392 9462 9404
rect 10689 9401 10701 9404
rect 10735 9401 10747 9435
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 10689 9395 10747 9401
rect 11532 9404 12817 9432
rect 9674 9364 9680 9376
rect 9140 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10597 9367 10655 9373
rect 10597 9364 10609 9367
rect 10468 9336 10609 9364
rect 10468 9324 10474 9336
rect 10597 9333 10609 9336
rect 10643 9333 10655 9367
rect 10597 9327 10655 9333
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11238 9364 11244 9376
rect 11195 9336 11244 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11532 9373 11560 9404
rect 12805 9401 12817 9404
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 13357 9435 13415 9441
rect 13357 9432 13369 9435
rect 13136 9404 13369 9432
rect 13136 9392 13142 9404
rect 13357 9401 13369 9404
rect 13403 9432 13415 9435
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 13403 9404 14105 9432
rect 13403 9401 13415 9404
rect 13357 9395 13415 9401
rect 14093 9401 14105 9404
rect 14139 9432 14151 9435
rect 16022 9432 16028 9444
rect 14139 9404 16028 9432
rect 14139 9401 14151 9404
rect 14093 9395 14151 9401
rect 16022 9392 16028 9404
rect 16080 9392 16086 9444
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9333 11575 9367
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 11517 9327 11575 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 13446 9364 13452 9376
rect 13407 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9364 13510 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13504 9336 14013 9364
rect 13504 9324 13510 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 14001 9327 14059 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 1857 9163 1915 9169
rect 1857 9160 1869 9163
rect 1820 9132 1869 9160
rect 1820 9120 1826 9132
rect 1857 9129 1869 9132
rect 1903 9129 1915 9163
rect 1857 9123 1915 9129
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2363 9132 2789 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 5718 9160 5724 9172
rect 5679 9132 5724 9160
rect 2777 9123 2835 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7742 9160 7748 9172
rect 7699 9132 7748 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8202 9160 8208 9172
rect 8159 9132 8208 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 9214 9160 9220 9172
rect 8803 9132 9220 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 10962 9160 10968 9172
rect 9548 9132 10968 9160
rect 9548 9120 9554 9132
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11146 9160 11152 9172
rect 11107 9132 11152 9160
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11940 9132 11989 9160
rect 11940 9120 11946 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 11977 9123 12035 9129
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 12526 9160 12532 9172
rect 12299 9132 12532 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 13044 9132 13093 9160
rect 13044 9120 13050 9132
rect 13081 9129 13093 9132
rect 13127 9160 13139 9163
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13127 9132 13737 9160
rect 13127 9129 13139 9132
rect 13081 9123 13139 9129
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 13814 9092 13820 9104
rect 4120 9064 10088 9092
rect 4120 9052 4126 9064
rect 2038 8984 2044 9036
rect 2096 9024 2102 9036
rect 2225 9027 2283 9033
rect 2225 9024 2237 9027
rect 2096 8996 2237 9024
rect 2096 8984 2102 8996
rect 2225 8993 2237 8996
rect 2271 8993 2283 9027
rect 2225 8987 2283 8993
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3510 9024 3516 9036
rect 3191 8996 3516 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 4608 9027 4666 9033
rect 4608 8993 4620 9027
rect 4654 9024 4666 9027
rect 5534 9024 5540 9036
rect 4654 8996 5540 9024
rect 4654 8993 4666 8996
rect 4608 8987 4666 8993
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 6069 9027 6127 9033
rect 6069 9024 6081 9027
rect 5776 8996 6081 9024
rect 5776 8984 5782 8996
rect 6069 8993 6081 8996
rect 6115 8993 6127 9027
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 6069 8987 6127 8993
rect 8018 8984 8024 8996
rect 8076 9024 8082 9036
rect 8478 9024 8484 9036
rect 8076 8996 8484 9024
rect 8076 8984 8082 8996
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 9024 8723 9027
rect 8938 9024 8944 9036
rect 8711 8996 8944 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 9122 9024 9128 9036
rect 9083 8996 9128 9024
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 9950 9033 9956 9036
rect 9944 9024 9956 9033
rect 9416 8996 9956 9024
rect 2498 8956 2504 8968
rect 2459 8928 2504 8956
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 3234 8956 3240 8968
rect 3195 8928 3240 8956
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3418 8956 3424 8968
rect 3379 8928 3424 8956
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 5810 8956 5816 8968
rect 5723 8928 5816 8956
rect 4341 8919 4399 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 4356 8888 4384 8919
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 9416 8965 9444 8996
rect 9944 8987 9956 8996
rect 9950 8984 9956 8987
rect 10008 8984 10014 9036
rect 10060 9024 10088 9064
rect 10796 9064 13820 9092
rect 10796 9024 10824 9064
rect 13814 9052 13820 9064
rect 13872 9092 13878 9104
rect 14734 9092 14740 9104
rect 13872 9064 14740 9092
rect 13872 9052 13878 9064
rect 14734 9052 14740 9064
rect 14792 9052 14798 9104
rect 10060 8996 10824 9024
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 11204 8996 11529 9024
rect 11204 8984 11210 8996
rect 11517 8993 11529 8996
rect 11563 8993 11575 9027
rect 11517 8987 11575 8993
rect 11624 8996 12020 9024
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8925 9459 8959
rect 9674 8956 9680 8968
rect 9635 8928 9680 8956
rect 9401 8919 9459 8925
rect 1912 8860 4384 8888
rect 1912 8848 1918 8860
rect 4356 8820 4384 8860
rect 5828 8820 5856 8916
rect 7190 8888 7196 8900
rect 7103 8860 7196 8888
rect 7190 8848 7196 8860
rect 7248 8888 7254 8900
rect 8220 8888 8248 8919
rect 7248 8860 8248 8888
rect 7248 8848 7254 8860
rect 4356 8792 5856 8820
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7285 8823 7343 8829
rect 7285 8820 7297 8823
rect 7156 8792 7297 8820
rect 7156 8780 7162 8792
rect 7285 8789 7297 8792
rect 7331 8789 7343 8823
rect 7285 8783 7343 8789
rect 7834 8780 7840 8832
rect 7892 8820 7898 8832
rect 8478 8820 8484 8832
rect 7892 8792 8484 8820
rect 7892 8780 7898 8792
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 9232 8820 9260 8919
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 11624 8965 11652 8996
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 10928 8928 11621 8956
rect 10928 8916 10934 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11790 8956 11796 8968
rect 11751 8928 11796 8956
rect 11609 8919 11667 8925
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 10962 8848 10968 8900
rect 11020 8888 11026 8900
rect 11882 8888 11888 8900
rect 11020 8860 11888 8888
rect 11020 8848 11026 8860
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 11992 8888 12020 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 13630 9024 13636 9036
rect 12492 8996 12537 9024
rect 13591 8996 13636 9024
rect 12492 8984 12498 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 12986 8916 12992 8968
rect 13044 8956 13050 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13044 8928 13829 8956
rect 13044 8916 13050 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 12529 8891 12587 8897
rect 12529 8888 12541 8891
rect 11992 8860 12541 8888
rect 12529 8857 12541 8860
rect 12575 8857 12587 8891
rect 12529 8851 12587 8857
rect 9858 8820 9864 8832
rect 9232 8792 9864 8820
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 10778 8820 10784 8832
rect 10100 8792 10784 8820
rect 10100 8780 10106 8792
rect 10778 8780 10784 8792
rect 10836 8820 10842 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10836 8792 11069 8820
rect 10836 8780 10842 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 13078 8820 13084 8832
rect 11296 8792 13084 8820
rect 11296 8780 11302 8792
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13262 8820 13268 8832
rect 13223 8792 13268 8820
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 3510 8616 3516 8628
rect 3471 8588 3516 8616
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5258 8616 5264 8628
rect 4939 8588 5264 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 5408 8588 5733 8616
rect 5408 8576 5414 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 6914 8616 6920 8628
rect 5721 8579 5779 8585
rect 5828 8588 6920 8616
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 5828 8548 5856 8588
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 9214 8616 9220 8628
rect 9175 8588 9220 8616
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 10321 8619 10379 8625
rect 10321 8585 10333 8619
rect 10367 8616 10379 8619
rect 11238 8616 11244 8628
rect 10367 8588 11244 8616
rect 10367 8585 10379 8588
rect 10321 8579 10379 8585
rect 11238 8576 11244 8588
rect 11296 8616 11302 8628
rect 12434 8616 12440 8628
rect 11296 8588 12440 8616
rect 11296 8576 11302 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 17218 8616 17224 8628
rect 12544 8588 17224 8616
rect 4212 8520 5856 8548
rect 4212 8508 4218 8520
rect 5902 8508 5908 8560
rect 5960 8548 5966 8560
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 5960 8520 7665 8548
rect 5960 8508 5966 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 7653 8511 7711 8517
rect 8389 8551 8447 8557
rect 8389 8517 8401 8551
rect 8435 8548 8447 8551
rect 9398 8548 9404 8560
rect 8435 8520 9404 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 9398 8508 9404 8520
rect 9456 8508 9462 8560
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 9548 8520 10548 8548
rect 9548 8508 9554 8520
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4433 8483 4491 8489
rect 4433 8480 4445 8483
rect 4065 8443 4123 8449
rect 4172 8452 4445 8480
rect 2124 8415 2182 8421
rect 2124 8381 2136 8415
rect 2170 8412 2182 8415
rect 3142 8412 3148 8424
rect 2170 8384 3148 8412
rect 2170 8381 2182 8384
rect 2124 8375 2182 8381
rect 3142 8372 3148 8384
rect 3200 8412 3206 8424
rect 4080 8412 4108 8443
rect 3200 8384 4108 8412
rect 3200 8372 3206 8384
rect 3418 8344 3424 8356
rect 3252 8316 3424 8344
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3252 8285 3280 8316
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4172 8344 4200 8452
rect 4433 8449 4445 8452
rect 4479 8480 4491 8483
rect 5537 8483 5595 8489
rect 4479 8452 5488 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 5074 8412 5080 8424
rect 4304 8384 5080 8412
rect 4304 8372 4310 8384
rect 5074 8372 5080 8384
rect 5132 8412 5138 8424
rect 5353 8415 5411 8421
rect 5353 8412 5365 8415
rect 5132 8384 5365 8412
rect 5132 8372 5138 8384
rect 5353 8381 5365 8384
rect 5399 8381 5411 8415
rect 5460 8412 5488 8452
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 6273 8483 6331 8489
rect 6273 8480 6285 8483
rect 5583 8452 6285 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 5810 8412 5816 8424
rect 5460 8384 5816 8412
rect 5353 8375 5411 8381
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 4019 8316 4200 8344
rect 4617 8347 4675 8353
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 5261 8347 5319 8353
rect 5261 8344 5273 8347
rect 4663 8316 5273 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 5261 8313 5273 8316
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 5920 8344 5948 8452
rect 6273 8449 6285 8452
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 6420 8452 7389 8480
rect 6420 8440 6426 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 8849 8483 8907 8489
rect 8849 8480 8861 8483
rect 8352 8452 8861 8480
rect 8352 8440 8358 8452
rect 8849 8449 8861 8452
rect 8895 8449 8907 8483
rect 8849 8443 8907 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8480 9091 8483
rect 9766 8480 9772 8492
rect 9079 8452 9168 8480
rect 9079 8449 9091 8452
rect 9033 8443 9091 8449
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8412 6147 8415
rect 7098 8412 7104 8424
rect 6135 8384 7104 8412
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7466 8412 7472 8424
rect 7331 8384 7472 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 7834 8412 7840 8424
rect 7795 8384 7840 8412
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 9140 8412 9168 8452
rect 9324 8452 9772 8480
rect 9324 8412 9352 8452
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10410 8480 10416 8492
rect 10091 8452 10416 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10520 8480 10548 8520
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10689 8551 10747 8557
rect 10689 8548 10701 8551
rect 10652 8520 10701 8548
rect 10652 8508 10658 8520
rect 10689 8517 10701 8520
rect 10735 8517 10747 8551
rect 11146 8548 11152 8560
rect 11059 8520 11152 8548
rect 10689 8511 10747 8517
rect 11072 8480 11100 8520
rect 11146 8508 11152 8520
rect 11204 8548 11210 8560
rect 11517 8551 11575 8557
rect 11517 8548 11529 8551
rect 11204 8520 11529 8548
rect 11204 8508 11210 8520
rect 11517 8517 11529 8520
rect 11563 8517 11575 8551
rect 11517 8511 11575 8517
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 12544 8548 12572 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 13446 8548 13452 8560
rect 11940 8520 12572 8548
rect 12820 8520 13452 8548
rect 11940 8508 11946 8520
rect 12820 8492 12848 8520
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 10520 8452 11100 8480
rect 9140 8384 9352 8412
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 9548 8384 9597 8412
rect 9548 8372 9554 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9916 8384 10517 8412
rect 9916 8372 9922 8384
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 11072 8412 11100 8452
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8449 11299 8483
rect 11241 8443 11299 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8480 11851 8483
rect 11974 8480 11980 8492
rect 11839 8452 11980 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 11072 8384 11161 8412
rect 10505 8375 10563 8381
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 5592 8316 5948 8344
rect 6181 8347 6239 8353
rect 5592 8304 5598 8316
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 8113 8347 8171 8353
rect 6227 8316 6868 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 3237 8279 3295 8285
rect 3237 8276 3249 8279
rect 2832 8248 3249 8276
rect 2832 8236 2838 8248
rect 3237 8245 3249 8248
rect 3283 8245 3295 8279
rect 3237 8239 3295 8245
rect 3329 8279 3387 8285
rect 3329 8245 3341 8279
rect 3375 8276 3387 8279
rect 3878 8276 3884 8288
rect 3375 8248 3884 8276
rect 3375 8245 3387 8248
rect 3329 8239 3387 8245
rect 3878 8236 3884 8248
rect 3936 8276 3942 8288
rect 5350 8276 5356 8288
rect 3936 8248 5356 8276
rect 3936 8236 3942 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 6638 8276 6644 8288
rect 6599 8248 6644 8276
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 6840 8285 6868 8316
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 8294 8344 8300 8356
rect 8159 8316 8300 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9030 8344 9036 8356
rect 8720 8316 9036 8344
rect 8720 8304 8726 8316
rect 9030 8304 9036 8316
rect 9088 8344 9094 8356
rect 9677 8347 9735 8353
rect 9677 8344 9689 8347
rect 9088 8316 9689 8344
rect 9088 8304 9094 8316
rect 9677 8313 9689 8316
rect 9723 8313 9735 8347
rect 11256 8344 11284 8443
rect 9677 8307 9735 8313
rect 10428 8316 11284 8344
rect 6825 8279 6883 8285
rect 6825 8245 6837 8279
rect 6871 8245 6883 8279
rect 7190 8276 7196 8288
rect 7151 8248 7196 8276
rect 6825 8239 6883 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 8205 8279 8263 8285
rect 8205 8245 8217 8279
rect 8251 8276 8263 8279
rect 8386 8276 8392 8288
rect 8251 8248 8392 8276
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 8754 8276 8760 8288
rect 8444 8248 8760 8276
rect 8444 8236 8450 8248
rect 8754 8236 8760 8248
rect 8812 8236 8818 8288
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 10428 8276 10456 8316
rect 9180 8248 10456 8276
rect 11057 8279 11115 8285
rect 9180 8236 9186 8248
rect 11057 8245 11069 8279
rect 11103 8276 11115 8279
rect 11808 8276 11836 8443
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12802 8480 12808 8492
rect 12492 8452 12808 8480
rect 12492 8440 12498 8452
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 13044 8452 13369 8480
rect 13044 8440 13050 8452
rect 13357 8449 13369 8452
rect 13403 8449 13415 8483
rect 13630 8480 13636 8492
rect 13591 8452 13636 8480
rect 13357 8443 13415 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 12584 8384 14197 8412
rect 12584 8372 12590 8384
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 16224 8412 16252 8443
rect 15620 8384 16252 8412
rect 15620 8372 15626 8384
rect 12618 8344 12624 8356
rect 12579 8316 12624 8344
rect 12618 8304 12624 8316
rect 12676 8344 12682 8356
rect 13173 8347 13231 8353
rect 13173 8344 13185 8347
rect 12676 8316 13185 8344
rect 12676 8304 12682 8316
rect 13173 8313 13185 8316
rect 13219 8313 13231 8347
rect 13173 8307 13231 8313
rect 13265 8347 13323 8353
rect 13265 8313 13277 8347
rect 13311 8344 13323 8347
rect 13446 8344 13452 8356
rect 13311 8316 13452 8344
rect 13311 8313 13323 8316
rect 13265 8307 13323 8313
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 14366 8304 14372 8356
rect 14424 8353 14430 8356
rect 14424 8347 14488 8353
rect 14424 8313 14442 8347
rect 14476 8313 14488 8347
rect 14424 8307 14488 8313
rect 14424 8304 14430 8307
rect 14642 8304 14648 8356
rect 14700 8344 14706 8356
rect 16025 8347 16083 8353
rect 16025 8344 16037 8347
rect 14700 8316 16037 8344
rect 14700 8304 14706 8316
rect 16025 8313 16037 8316
rect 16071 8313 16083 8347
rect 16025 8307 16083 8313
rect 11103 8248 11836 8276
rect 12805 8279 12863 8285
rect 11103 8245 11115 8248
rect 11057 8239 11115 8245
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 13078 8276 13084 8288
rect 12851 8248 13084 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 15562 8276 15568 8288
rect 15523 8248 15568 8276
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 15712 8248 15757 8276
rect 15712 8236 15718 8248
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 16172 8248 16217 8276
rect 16172 8236 16178 8248
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2682 8072 2688 8084
rect 2556 8044 2688 8072
rect 2556 8032 2562 8044
rect 2682 8032 2688 8044
rect 2740 8072 2746 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2740 8044 2789 8072
rect 2740 8032 2746 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 4157 8075 4215 8081
rect 4157 8072 4169 8075
rect 3283 8044 4169 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 4157 8041 4169 8044
rect 4203 8072 4215 8075
rect 5442 8072 5448 8084
rect 4203 8044 5448 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5592 8044 5825 8072
rect 5592 8032 5598 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 5813 8035 5871 8041
rect 5997 8075 6055 8081
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 7282 8072 7288 8084
rect 6043 8044 7288 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 7282 8032 7288 8044
rect 7340 8072 7346 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7340 8044 7481 8072
rect 7340 8032 7346 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 14553 8075 14611 8081
rect 7469 8035 7527 8041
rect 8772 8044 14504 8072
rect 1854 8004 1860 8016
rect 1412 7976 1860 8004
rect 1412 7945 1440 7976
rect 1854 7964 1860 7976
rect 1912 7964 1918 8016
rect 4700 8007 4758 8013
rect 4700 7973 4712 8007
rect 4746 8004 4758 8007
rect 6086 8004 6092 8016
rect 4746 7976 6092 8004
rect 4746 7973 4758 7976
rect 4700 7967 4758 7973
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 8294 8004 8300 8016
rect 6380 7976 8300 8004
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 1397 7899 1455 7905
rect 1664 7939 1722 7945
rect 1664 7905 1676 7939
rect 1710 7936 1722 7939
rect 2774 7936 2780 7948
rect 1710 7908 2780 7936
rect 1710 7905 1722 7908
rect 1664 7899 1722 7905
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3375 7908 3832 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3142 7760 3148 7812
rect 3200 7800 3206 7812
rect 3436 7800 3464 7831
rect 3804 7809 3832 7908
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 6380 7936 6408 7976
rect 8294 7964 8300 7976
rect 8352 7964 8358 8016
rect 4120 7908 6408 7936
rect 4120 7896 4126 7908
rect 6454 7896 6460 7948
rect 6512 7936 6518 7948
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6512 7908 6561 7936
rect 6512 7896 6518 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 6972 7908 7389 7936
rect 6972 7896 6978 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7466 7896 7472 7948
rect 7524 7936 7530 7948
rect 8021 7939 8079 7945
rect 8021 7936 8033 7939
rect 7524 7908 8033 7936
rect 7524 7896 7530 7908
rect 8021 7905 8033 7908
rect 8067 7936 8079 7939
rect 8772 7936 8800 8044
rect 10680 8007 10738 8013
rect 10680 7973 10692 8007
rect 10726 8004 10738 8007
rect 10778 8004 10784 8016
rect 10726 7976 10784 8004
rect 10726 7973 10738 7976
rect 10680 7967 10738 7973
rect 10778 7964 10784 7976
rect 10836 7964 10842 8016
rect 10870 7964 10876 8016
rect 10928 7964 10934 8016
rect 12888 8007 12946 8013
rect 12888 7973 12900 8007
rect 12934 8004 12946 8007
rect 12986 8004 12992 8016
rect 12934 7976 12992 8004
rect 12934 7973 12946 7976
rect 12888 7967 12946 7973
rect 12986 7964 12992 7976
rect 13044 7964 13050 8016
rect 14476 8004 14504 8044
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 15289 8075 15347 8081
rect 15289 8072 15301 8075
rect 14599 8044 15301 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 15289 8041 15301 8044
rect 15335 8041 15347 8075
rect 15289 8035 15347 8041
rect 15010 8004 15016 8016
rect 14476 7976 15016 8004
rect 15010 7964 15016 7976
rect 15068 8004 15074 8016
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 15068 7976 15761 8004
rect 15068 7964 15074 7976
rect 15749 7973 15761 7976
rect 15795 8004 15807 8007
rect 16758 8004 16764 8016
rect 15795 7976 16764 8004
rect 15795 7973 15807 7976
rect 15749 7967 15807 7973
rect 16758 7964 16764 7976
rect 16816 7964 16822 8016
rect 8067 7908 8800 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 9732 7908 10425 7936
rect 9732 7896 9738 7908
rect 10413 7905 10425 7908
rect 10459 7936 10471 7939
rect 10888 7936 10916 7964
rect 12526 7936 12532 7948
rect 10459 7908 12532 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 12526 7896 12532 7908
rect 12584 7936 12590 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12584 7908 12633 7936
rect 12584 7896 12590 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 14458 7936 14464 7948
rect 14419 7908 14464 7936
rect 12621 7899 12679 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 15105 7939 15163 7945
rect 15105 7905 15117 7939
rect 15151 7936 15163 7939
rect 15470 7936 15476 7948
rect 15151 7908 15476 7936
rect 15151 7905 15163 7908
rect 15105 7899 15163 7905
rect 15470 7896 15476 7908
rect 15528 7936 15534 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15528 7908 15669 7936
rect 15528 7896 15534 7908
rect 15657 7905 15669 7908
rect 15703 7936 15715 7939
rect 15838 7936 15844 7948
rect 15703 7908 15844 7936
rect 15703 7905 15715 7908
rect 15657 7899 15715 7905
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 3200 7772 3464 7800
rect 3789 7803 3847 7809
rect 3200 7760 3206 7772
rect 3789 7769 3801 7803
rect 3835 7800 3847 7803
rect 4154 7800 4160 7812
rect 3835 7772 4160 7800
rect 3835 7769 3847 7772
rect 3789 7763 3847 7769
rect 4154 7760 4160 7772
rect 4212 7760 4218 7812
rect 2866 7732 2872 7744
rect 2827 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4448 7732 4476 7831
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6362 7868 6368 7880
rect 6144 7840 6368 7868
rect 6144 7828 6150 7840
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 6871 7840 7573 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7561 7837 7573 7840
rect 7607 7868 7619 7871
rect 7650 7868 7656 7880
rect 7607 7840 7656 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 14366 7868 14372 7880
rect 14016 7840 14372 7868
rect 5552 7800 5580 7828
rect 5718 7800 5724 7812
rect 5552 7772 5724 7800
rect 5718 7760 5724 7772
rect 5776 7800 5782 7812
rect 6546 7800 6552 7812
rect 5776 7772 6552 7800
rect 5776 7760 5782 7772
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 5074 7732 5080 7744
rect 4448 7704 5080 7732
rect 5074 7692 5080 7704
rect 5132 7692 5138 7744
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6362 7732 6368 7744
rect 6227 7704 6368 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 7006 7732 7012 7744
rect 6967 7704 7012 7732
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 7837 7735 7895 7741
rect 7837 7732 7849 7735
rect 7248 7704 7849 7732
rect 7248 7692 7254 7704
rect 7837 7701 7849 7704
rect 7883 7701 7895 7735
rect 7837 7695 7895 7701
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 8720 7704 8861 7732
rect 8720 7692 8726 7704
rect 8849 7701 8861 7704
rect 8895 7701 8907 7735
rect 8849 7695 8907 7701
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 9214 7732 9220 7744
rect 9171 7704 9220 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 9214 7692 9220 7704
rect 9272 7732 9278 7744
rect 9490 7732 9496 7744
rect 9272 7704 9496 7732
rect 9272 7692 9278 7704
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 11790 7732 11796 7744
rect 11751 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14016 7741 14044 7840
rect 14366 7828 14372 7840
rect 14424 7868 14430 7880
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14424 7840 14657 7868
rect 14424 7828 14430 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 15930 7868 15936 7880
rect 15891 7840 15936 7868
rect 14645 7831 14703 7837
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 14093 7803 14151 7809
rect 14093 7769 14105 7803
rect 14139 7800 14151 7803
rect 16114 7800 16120 7812
rect 14139 7772 16120 7800
rect 14139 7769 14151 7772
rect 14093 7763 14151 7769
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 14001 7735 14059 7741
rect 14001 7732 14013 7735
rect 13964 7704 14013 7732
rect 13964 7692 13970 7704
rect 14001 7701 14013 7704
rect 14047 7701 14059 7735
rect 14001 7695 14059 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3513 7531 3571 7537
rect 3513 7528 3525 7531
rect 3292 7500 3525 7528
rect 3292 7488 3298 7500
rect 3513 7497 3525 7500
rect 3559 7497 3571 7531
rect 3513 7491 3571 7497
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 4338 7528 4344 7540
rect 4120 7500 4344 7528
rect 4120 7488 4126 7500
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5316 7500 5365 7528
rect 5316 7488 5322 7500
rect 5353 7497 5365 7500
rect 5399 7528 5411 7531
rect 6454 7528 6460 7540
rect 5399 7500 6460 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 8849 7531 8907 7537
rect 8849 7497 8861 7531
rect 8895 7528 8907 7531
rect 9122 7528 9128 7540
rect 8895 7500 9128 7528
rect 8895 7497 8907 7500
rect 8849 7491 8907 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 14642 7528 14648 7540
rect 13311 7500 14648 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 15010 7528 15016 7540
rect 14971 7500 15016 7528
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 2225 7463 2283 7469
rect 2225 7429 2237 7463
rect 2271 7460 2283 7463
rect 3326 7460 3332 7472
rect 2271 7432 3332 7460
rect 2271 7429 2283 7432
rect 2225 7423 2283 7429
rect 2792 7401 2820 7432
rect 3326 7420 3332 7432
rect 3384 7420 3390 7472
rect 8754 7420 8760 7472
rect 8812 7460 8818 7472
rect 9217 7463 9275 7469
rect 9217 7460 9229 7463
rect 8812 7432 9229 7460
rect 8812 7420 8818 7432
rect 9217 7429 9229 7432
rect 9263 7460 9275 7463
rect 11333 7463 11391 7469
rect 9263 7432 9904 7460
rect 9263 7429 9275 7432
rect 9217 7423 9275 7429
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 2961 7395 3019 7401
rect 2823 7364 2857 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3142 7392 3148 7404
rect 3007 7364 3148 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3200 7364 4077 7392
rect 3200 7352 3206 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 6362 7392 6368 7404
rect 6323 7364 6368 7392
rect 4065 7355 4123 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 6730 7392 6736 7404
rect 6595 7364 6736 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 9876 7401 9904 7432
rect 11333 7429 11345 7463
rect 11379 7460 11391 7463
rect 11882 7460 11888 7472
rect 11379 7432 11888 7460
rect 11379 7429 11391 7432
rect 11333 7423 11391 7429
rect 11882 7420 11888 7432
rect 11940 7420 11946 7472
rect 12437 7463 12495 7469
rect 12437 7429 12449 7463
rect 12483 7460 12495 7463
rect 14734 7460 14740 7472
rect 12483 7432 14740 7460
rect 12483 7429 12495 7432
rect 12437 7423 12495 7429
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 10318 7392 10324 7404
rect 10091 7364 10324 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 12342 7352 12348 7404
rect 12400 7352 12406 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12768 7364 13001 7392
rect 12768 7352 12774 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 13136 7364 13737 7392
rect 13136 7352 13142 7364
rect 13725 7361 13737 7364
rect 13771 7361 13783 7395
rect 13906 7392 13912 7404
rect 13867 7364 13912 7392
rect 13725 7355 13783 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 5902 7324 5908 7336
rect 5767 7296 5908 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5902 7284 5908 7296
rect 5960 7284 5966 7336
rect 6273 7327 6331 7333
rect 6273 7293 6285 7327
rect 6319 7324 6331 7327
rect 7006 7324 7012 7336
rect 6319 7296 7012 7324
rect 6319 7293 6331 7296
rect 6273 7287 6331 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 2685 7259 2743 7265
rect 2685 7225 2697 7259
rect 2731 7256 2743 7259
rect 3145 7259 3203 7265
rect 3145 7256 3157 7259
rect 2731 7228 3157 7256
rect 2731 7225 2743 7228
rect 2685 7219 2743 7225
rect 3145 7225 3157 7228
rect 3191 7225 3203 7259
rect 3145 7219 3203 7225
rect 3973 7259 4031 7265
rect 3973 7225 3985 7259
rect 4019 7256 4031 7259
rect 4019 7228 4844 7256
rect 4019 7225 4031 7228
rect 3973 7219 4031 7225
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2406 7188 2412 7200
rect 2363 7160 2412 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3878 7148 3884 7160
rect 3936 7188 3942 7200
rect 4816 7197 4844 7228
rect 5166 7216 5172 7268
rect 5224 7256 5230 7268
rect 6454 7256 6460 7268
rect 5224 7228 6460 7256
rect 5224 7216 5230 7228
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 3936 7160 4537 7188
rect 3936 7148 3942 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 4525 7151 4583 7157
rect 4801 7191 4859 7197
rect 4801 7157 4813 7191
rect 4847 7188 4859 7191
rect 5258 7188 5264 7200
rect 4847 7160 5264 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5552 7197 5580 7228
rect 6454 7216 6460 7228
rect 6512 7256 6518 7268
rect 7484 7256 7512 7287
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11296 7296 11529 7324
rect 11296 7284 11302 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 11606 7284 11612 7336
rect 11664 7324 11670 7336
rect 12360 7324 12388 7352
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 11664 7296 12909 7324
rect 11664 7284 11670 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 15562 7333 15568 7336
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13320 7296 13645 7324
rect 13320 7284 13326 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 15289 7327 15347 7333
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 15556 7324 15568 7333
rect 15523 7296 15568 7324
rect 15289 7287 15347 7293
rect 15556 7287 15568 7296
rect 7742 7265 7748 7268
rect 6512 7228 7512 7256
rect 6512 7216 6518 7228
rect 7736 7219 7748 7265
rect 7800 7256 7806 7268
rect 7800 7228 7836 7256
rect 7742 7216 7748 7219
rect 7800 7216 7806 7228
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11112 7228 12296 7256
rect 11112 7216 11118 7228
rect 5537 7191 5595 7197
rect 5537 7157 5549 7191
rect 5583 7157 5595 7191
rect 5537 7151 5595 7157
rect 5905 7191 5963 7197
rect 5905 7157 5917 7191
rect 5951 7188 5963 7191
rect 8294 7188 8300 7200
rect 5951 7160 8300 7188
rect 5951 7157 5963 7160
rect 5905 7151 5963 7157
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9766 7188 9772 7200
rect 9727 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 11664 7160 12081 7188
rect 11664 7148 11670 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12268 7188 12296 7228
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12805 7259 12863 7265
rect 12805 7256 12817 7259
rect 12400 7228 12817 7256
rect 12400 7216 12406 7228
rect 12805 7225 12817 7228
rect 12851 7225 12863 7259
rect 12805 7219 12863 7225
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 15304 7256 15332 7287
rect 15562 7284 15568 7287
rect 15620 7284 15626 7336
rect 15470 7256 15476 7268
rect 13964 7228 15476 7256
rect 13964 7216 13970 7228
rect 15470 7216 15476 7228
rect 15528 7216 15534 7268
rect 12526 7188 12532 7200
rect 12268 7160 12532 7188
rect 12069 7151 12127 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 16666 7188 16672 7200
rect 16627 7160 16672 7188
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 3605 6987 3663 6993
rect 3605 6953 3617 6987
rect 3651 6984 3663 6987
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 3651 6956 4077 6984
rect 3651 6953 3663 6956
rect 3605 6947 3663 6953
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 4525 6987 4583 6993
rect 4525 6984 4537 6987
rect 4396 6956 4537 6984
rect 4396 6944 4402 6956
rect 4525 6953 4537 6956
rect 4571 6953 4583 6987
rect 4525 6947 4583 6953
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7800 6956 7849 6984
rect 7800 6944 7806 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 7837 6947 7895 6953
rect 4433 6919 4491 6925
rect 4433 6885 4445 6919
rect 4479 6916 4491 6919
rect 4982 6916 4988 6928
rect 4479 6888 4988 6916
rect 4479 6885 4491 6888
rect 4433 6879 4491 6885
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 2866 6848 2872 6860
rect 2547 6820 2872 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2866 6808 2872 6820
rect 2924 6808 2930 6860
rect 3510 6848 3516 6860
rect 3471 6820 3516 6848
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 4448 6848 4476 6879
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 5994 6916 6000 6928
rect 5955 6888 6000 6916
rect 5994 6876 6000 6888
rect 6052 6876 6058 6928
rect 7852 6916 7880 6947
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 8444 6956 9229 6984
rect 8444 6944 8450 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 9217 6947 9275 6953
rect 9232 6916 9260 6947
rect 9766 6944 9772 6996
rect 9824 6984 9830 6996
rect 10505 6987 10563 6993
rect 10505 6984 10517 6987
rect 9824 6956 10517 6984
rect 9824 6944 9830 6956
rect 10505 6953 10517 6956
rect 10551 6953 10563 6987
rect 11606 6984 11612 6996
rect 10505 6947 10563 6953
rect 11072 6956 11612 6984
rect 10045 6919 10103 6925
rect 10045 6916 10057 6919
rect 7852 6888 8432 6916
rect 9232 6888 10057 6916
rect 3712 6820 4476 6848
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2774 6780 2780 6792
rect 2731 6752 2780 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6780 3111 6783
rect 3712 6780 3740 6820
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 5074 6848 5080 6860
rect 4948 6820 5080 6848
rect 4948 6808 4954 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 6730 6857 6736 6860
rect 6724 6848 6736 6857
rect 6288 6820 6736 6848
rect 3099 6752 3740 6780
rect 3789 6783 3847 6789
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3789 6749 3801 6783
rect 3835 6780 3847 6783
rect 3970 6780 3976 6792
rect 3835 6752 3976 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5350 6780 5356 6792
rect 4755 6752 5356 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 6288 6789 6316 6820
rect 6724 6811 6736 6820
rect 6730 6808 6736 6811
rect 6788 6808 6794 6860
rect 8404 6848 8432 6888
rect 10045 6885 10057 6888
rect 10091 6885 10103 6919
rect 11072 6916 11100 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12434 6984 12440 6996
rect 12400 6956 12440 6984
rect 12400 6944 12406 6956
rect 12434 6944 12440 6956
rect 12492 6944 12498 6996
rect 13814 6984 13820 6996
rect 13775 6956 13820 6984
rect 13814 6944 13820 6956
rect 13872 6984 13878 6996
rect 14277 6987 14335 6993
rect 14277 6984 14289 6987
rect 13872 6956 14289 6984
rect 13872 6944 13878 6956
rect 14277 6953 14289 6956
rect 14323 6953 14335 6987
rect 14277 6947 14335 6953
rect 10045 6879 10103 6885
rect 10152 6888 11100 6916
rect 11140 6919 11198 6925
rect 8404 6820 8524 6848
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6454 6780 6460 6792
rect 6415 6752 6460 6780
rect 6273 6743 6331 6749
rect 2038 6712 2044 6724
rect 1999 6684 2044 6712
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 4890 6672 4896 6724
rect 4948 6712 4954 6724
rect 5261 6715 5319 6721
rect 5261 6712 5273 6715
rect 4948 6684 5273 6712
rect 4948 6672 4954 6684
rect 5261 6681 5273 6684
rect 5307 6712 5319 6715
rect 5902 6712 5908 6724
rect 5307 6684 5908 6712
rect 5307 6681 5319 6684
rect 5261 6675 5319 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 6104 6712 6132 6743
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 8496 6789 8524 6820
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 10152 6848 10180 6888
rect 11140 6885 11152 6919
rect 11186 6916 11198 6919
rect 11790 6916 11796 6928
rect 11186 6888 11796 6916
rect 11186 6885 11198 6888
rect 11140 6879 11198 6885
rect 11790 6876 11796 6888
rect 11848 6876 11854 6928
rect 13556 6888 14780 6916
rect 8628 6820 10180 6848
rect 8628 6808 8634 6820
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 10284 6820 11928 6848
rect 10284 6808 10290 6820
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10318 6780 10324 6792
rect 10231 6752 10324 6780
rect 10137 6743 10195 6749
rect 6362 6712 6368 6724
rect 6104 6684 6368 6712
rect 6362 6672 6368 6684
rect 6420 6672 6426 6724
rect 8404 6712 8432 6743
rect 7392 6684 8432 6712
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3326 6644 3332 6656
rect 3191 6616 3332 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 5629 6647 5687 6653
rect 5629 6613 5641 6647
rect 5675 6644 5687 6647
rect 7392 6644 7420 6684
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 9677 6715 9735 6721
rect 9677 6712 9689 6715
rect 8996 6684 9689 6712
rect 8996 6672 9002 6684
rect 9677 6681 9689 6684
rect 9723 6681 9735 6715
rect 9677 6675 9735 6681
rect 5675 6616 7420 6644
rect 5675 6613 5687 6616
rect 5629 6607 5687 6613
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7616 6616 7941 6644
rect 7616 6604 7622 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 9214 6604 9220 6656
rect 9272 6644 9278 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9272 6616 9413 6644
rect 9272 6604 9278 6616
rect 9401 6613 9413 6616
rect 9447 6644 9459 6647
rect 10152 6644 10180 6743
rect 10318 6740 10324 6752
rect 10376 6780 10382 6792
rect 10376 6752 10824 6780
rect 10376 6740 10382 6752
rect 9447 6616 10180 6644
rect 10796 6644 10824 6752
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 11900 6780 11928 6820
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 13556 6848 13584 6888
rect 12032 6820 13584 6848
rect 13633 6851 13691 6857
rect 12032 6808 12038 6820
rect 13633 6817 13645 6851
rect 13679 6848 13691 6851
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 13679 6820 14381 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 14369 6817 14381 6820
rect 14415 6848 14427 6851
rect 14642 6848 14648 6860
rect 14415 6820 14648 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 13648 6780 13676 6811
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 14752 6848 14780 6888
rect 17586 6848 17592 6860
rect 14752 6820 17592 6848
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 14550 6780 14556 6792
rect 10928 6752 10973 6780
rect 11900 6752 13676 6780
rect 14511 6752 14556 6780
rect 10928 6740 10934 6752
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 14734 6780 14740 6792
rect 14695 6752 14740 6780
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 13078 6672 13084 6724
rect 13136 6712 13142 6724
rect 15194 6712 15200 6724
rect 13136 6684 15200 6712
rect 13136 6672 13142 6684
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 11974 6644 11980 6656
rect 10796 6616 11980 6644
rect 9447 6613 9459 6616
rect 9401 6607 9459 6613
rect 11974 6604 11980 6616
rect 12032 6644 12038 6656
rect 12253 6647 12311 6653
rect 12253 6644 12265 6647
rect 12032 6616 12265 6644
rect 12032 6604 12038 6616
rect 12253 6613 12265 6616
rect 12299 6613 12311 6647
rect 12253 6607 12311 6613
rect 13909 6647 13967 6653
rect 13909 6613 13921 6647
rect 13955 6644 13967 6647
rect 15746 6644 15752 6656
rect 13955 6616 15752 6644
rect 13955 6613 13967 6616
rect 13909 6607 13967 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 3050 6400 3056 6452
rect 3108 6440 3114 6452
rect 3237 6443 3295 6449
rect 3237 6440 3249 6443
rect 3108 6412 3249 6440
rect 3108 6400 3114 6412
rect 3237 6409 3249 6412
rect 3283 6440 3295 6443
rect 3602 6440 3608 6452
rect 3283 6412 3608 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4120 6412 6316 6440
rect 4120 6400 4126 6412
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 5166 6372 5172 6384
rect 4212 6344 5172 6372
rect 4212 6332 4218 6344
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 3142 6304 3148 6316
rect 2884 6276 3148 6304
rect 1854 6236 1860 6248
rect 1815 6208 1860 6236
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 2124 6171 2182 6177
rect 2124 6137 2136 6171
rect 2170 6168 2182 6171
rect 2884 6168 2912 6276
rect 3142 6264 3148 6276
rect 3200 6304 3206 6316
rect 3970 6304 3976 6316
rect 3200 6276 3976 6304
rect 3200 6264 3206 6276
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 4890 6304 4896 6316
rect 4847 6276 4896 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 6288 6304 6316 6412
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 7009 6443 7067 6449
rect 7009 6440 7021 6443
rect 6420 6412 7021 6440
rect 6420 6400 6426 6412
rect 7009 6409 7021 6412
rect 7055 6409 7067 6443
rect 12342 6440 12348 6452
rect 7009 6403 7067 6409
rect 7107 6412 12348 6440
rect 6641 6375 6699 6381
rect 6641 6341 6653 6375
rect 6687 6372 6699 6375
rect 6730 6372 6736 6384
rect 6687 6344 6736 6372
rect 6687 6341 6699 6344
rect 6641 6335 6699 6341
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 7107 6304 7135 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6440 12495 6443
rect 14458 6440 14464 6452
rect 12483 6412 14464 6440
rect 12483 6409 12495 6412
rect 12437 6403 12495 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 17678 6440 17684 6452
rect 14884 6412 17684 6440
rect 14884 6400 14890 6412
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 10468 6344 11989 6372
rect 10468 6332 10474 6344
rect 7650 6304 7656 6316
rect 5031 6276 5396 6304
rect 6288 6276 7135 6304
rect 7611 6276 7656 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5368 6248 5396 6276
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8938 6304 8944 6316
rect 8899 6276 8944 6304
rect 8938 6264 8944 6276
rect 8996 6264 9002 6316
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 11333 6307 11391 6313
rect 11333 6304 11345 6307
rect 9171 6276 9444 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4212 6208 4721 6236
rect 4212 6196 4218 6208
rect 4709 6205 4721 6208
rect 4755 6205 4767 6239
rect 5258 6236 5264 6248
rect 5219 6208 5264 6236
rect 4709 6199 4767 6205
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 5350 6196 5356 6248
rect 5408 6196 5414 6248
rect 5528 6239 5586 6245
rect 5528 6205 5540 6239
rect 5574 6236 5586 6239
rect 7668 6236 7696 6264
rect 9306 6236 9312 6248
rect 5574 6208 7696 6236
rect 9267 6208 9312 6236
rect 5574 6205 5586 6208
rect 5528 6199 5586 6205
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 9416 6236 9444 6276
rect 10765 6276 11345 6304
rect 9950 6236 9956 6248
rect 9416 6208 9956 6236
rect 9950 6196 9956 6208
rect 10008 6236 10014 6248
rect 10765 6236 10793 6276
rect 11333 6273 11345 6276
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 10008 6208 10793 6236
rect 10008 6196 10014 6208
rect 2170 6140 2912 6168
rect 2170 6137 2182 6140
rect 2124 6131 2182 6137
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 8849 6171 8907 6177
rect 4120 6140 8616 6168
rect 4120 6128 4126 6140
rect 3418 6100 3424 6112
rect 3379 6072 3424 6100
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 4341 6103 4399 6109
rect 4341 6100 4353 6103
rect 3927 6072 4353 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 4341 6069 4353 6072
rect 4387 6069 4399 6103
rect 7374 6100 7380 6112
rect 7335 6072 7380 6100
rect 4341 6063 4399 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7466 6060 7472 6112
rect 7524 6100 7530 6112
rect 7524 6072 7569 6100
rect 7524 6060 7530 6072
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7800 6072 7849 6100
rect 7800 6060 7806 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 8478 6100 8484 6112
rect 8439 6072 8484 6100
rect 7837 6063 7895 6069
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 8588 6100 8616 6140
rect 8849 6137 8861 6171
rect 8895 6168 8907 6171
rect 9398 6168 9404 6180
rect 8895 6140 9404 6168
rect 8895 6137 8907 6140
rect 8849 6131 8907 6137
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 9576 6171 9634 6177
rect 9576 6137 9588 6171
rect 9622 6168 9634 6171
rect 10318 6168 10324 6180
rect 9622 6140 10324 6168
rect 9622 6137 9634 6140
rect 9576 6131 9634 6137
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 10765 6168 10793 6208
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11149 6239 11207 6245
rect 11149 6236 11161 6239
rect 11112 6208 11161 6236
rect 11112 6196 11118 6208
rect 11149 6205 11161 6208
rect 11195 6205 11207 6239
rect 11149 6199 11207 6205
rect 11241 6239 11299 6245
rect 11241 6205 11253 6239
rect 11287 6236 11299 6239
rect 11422 6236 11428 6248
rect 11287 6208 11428 6236
rect 11287 6205 11299 6208
rect 11241 6199 11299 6205
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 11808 6168 11836 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 15194 6372 15200 6384
rect 15107 6344 15200 6372
rect 11977 6335 12035 6341
rect 15194 6332 15200 6344
rect 15252 6372 15258 6384
rect 15930 6372 15936 6384
rect 15252 6344 15936 6372
rect 15252 6332 15258 6344
rect 15930 6332 15936 6344
rect 15988 6332 15994 6384
rect 13078 6304 13084 6316
rect 13039 6276 13084 6304
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12544 6208 12817 6236
rect 12544 6168 12572 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 13817 6239 13875 6245
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 13906 6236 13912 6248
rect 13863 6208 13912 6236
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 12897 6171 12955 6177
rect 12897 6168 12909 6171
rect 10704 6140 10793 6168
rect 11164 6140 11376 6168
rect 11808 6140 12572 6168
rect 12636 6140 12909 6168
rect 10226 6100 10232 6112
rect 8588 6072 10232 6100
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10704 6109 10732 6140
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 10836 6072 10881 6100
rect 10836 6060 10842 6072
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11164 6100 11192 6140
rect 11020 6072 11192 6100
rect 11348 6100 11376 6140
rect 12161 6103 12219 6109
rect 12161 6100 12173 6103
rect 11348 6072 12173 6100
rect 11020 6060 11026 6072
rect 12161 6069 12173 6072
rect 12207 6100 12219 6103
rect 12636 6100 12664 6140
rect 12897 6137 12909 6140
rect 12943 6137 12955 6171
rect 12897 6131 12955 6137
rect 13078 6128 13084 6180
rect 13136 6168 13142 6180
rect 13832 6168 13860 6199
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 14084 6239 14142 6245
rect 14084 6205 14096 6239
rect 14130 6236 14142 6239
rect 14458 6236 14464 6248
rect 14130 6208 14464 6236
rect 14130 6205 14142 6208
rect 14084 6199 14142 6205
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 15856 6236 15884 6267
rect 14700 6208 15884 6236
rect 14700 6196 14706 6208
rect 16022 6196 16028 6248
rect 16080 6236 16086 6248
rect 16393 6239 16451 6245
rect 16393 6236 16405 6239
rect 16080 6208 16405 6236
rect 16080 6196 16086 6208
rect 16393 6205 16405 6208
rect 16439 6205 16451 6239
rect 16393 6199 16451 6205
rect 13136 6140 13860 6168
rect 13136 6128 13142 6140
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 15657 6171 15715 6177
rect 15657 6168 15669 6171
rect 14240 6140 15669 6168
rect 14240 6128 14246 6140
rect 15657 6137 15669 6140
rect 15703 6137 15715 6171
rect 15657 6131 15715 6137
rect 16660 6171 16718 6177
rect 16660 6137 16672 6171
rect 16706 6168 16718 6171
rect 17402 6168 17408 6180
rect 16706 6140 17408 6168
rect 16706 6137 16718 6140
rect 16660 6131 16718 6137
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 12207 6072 12664 6100
rect 12207 6069 12219 6072
rect 12161 6063 12219 6069
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14550 6100 14556 6112
rect 14332 6072 14556 6100
rect 14332 6060 14338 6072
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 15286 6100 15292 6112
rect 15247 6072 15292 6100
rect 15286 6060 15292 6072
rect 15344 6060 15350 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 17773 6103 17831 6109
rect 17773 6100 17785 6103
rect 15436 6072 17785 6100
rect 15436 6060 15442 6072
rect 17773 6069 17785 6072
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 3142 5896 3148 5908
rect 3103 5868 3148 5896
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 3605 5899 3663 5905
rect 3605 5896 3617 5899
rect 3568 5868 3617 5896
rect 3568 5856 3574 5868
rect 3605 5865 3617 5868
rect 3651 5865 3663 5899
rect 3605 5859 3663 5865
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4890 5896 4896 5908
rect 4764 5868 4896 5896
rect 4764 5856 4770 5868
rect 4890 5856 4896 5868
rect 4948 5896 4954 5908
rect 5258 5896 5264 5908
rect 4948 5868 5264 5896
rect 4948 5856 4954 5868
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5902 5896 5908 5908
rect 5592 5868 5908 5896
rect 5592 5856 5598 5868
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 6086 5896 6092 5908
rect 6047 5868 6092 5896
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7524 5868 7941 5896
rect 7524 5856 7530 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 8297 5899 8355 5905
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 8386 5896 8392 5908
rect 8343 5868 8392 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8536 5868 9137 5896
rect 8536 5856 8542 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9217 5899 9275 5905
rect 9217 5865 9229 5899
rect 9263 5896 9275 5899
rect 10778 5896 10784 5908
rect 9263 5868 10784 5896
rect 9263 5865 9275 5868
rect 9217 5859 9275 5865
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 11020 5868 11069 5896
rect 11020 5856 11026 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 14093 5899 14151 5905
rect 14093 5865 14105 5899
rect 14139 5896 14151 5899
rect 14182 5896 14188 5908
rect 14139 5868 14188 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14461 5899 14519 5905
rect 14461 5865 14473 5899
rect 14507 5896 14519 5899
rect 14734 5896 14740 5908
rect 14507 5868 14740 5896
rect 14507 5865 14519 5868
rect 14461 5859 14519 5865
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 17678 5856 17684 5908
rect 17736 5896 17742 5908
rect 17957 5899 18015 5905
rect 17957 5896 17969 5899
rect 17736 5868 17969 5896
rect 17736 5856 17742 5868
rect 17957 5865 17969 5868
rect 18003 5865 18015 5899
rect 17957 5859 18015 5865
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 6724 5831 6782 5837
rect 4120 5800 5396 5828
rect 4120 5788 4126 5800
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 1854 5760 1860 5772
rect 1811 5732 1860 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 2032 5763 2090 5769
rect 2032 5729 2044 5763
rect 2078 5760 2090 5763
rect 4080 5760 4108 5788
rect 5368 5772 5396 5800
rect 6724 5797 6736 5831
rect 6770 5828 6782 5831
rect 8202 5828 8208 5840
rect 6770 5800 8208 5828
rect 6770 5797 6782 5800
rect 6724 5791 6782 5797
rect 8202 5788 8208 5800
rect 8260 5828 8266 5840
rect 9674 5828 9680 5840
rect 8260 5800 8432 5828
rect 8260 5788 8266 5800
rect 4706 5760 4712 5772
rect 2078 5732 4108 5760
rect 4667 5732 4712 5760
rect 2078 5729 2090 5732
rect 2032 5723 2090 5729
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 4976 5763 5034 5769
rect 4976 5729 4988 5763
rect 5022 5760 5034 5763
rect 5258 5760 5264 5772
rect 5022 5732 5264 5760
rect 5022 5729 5034 5732
rect 4976 5723 5034 5729
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 8404 5760 8432 5800
rect 8588 5800 9680 5828
rect 5408 5732 7972 5760
rect 8404 5732 8524 5760
rect 5408 5720 5414 5732
rect 6454 5692 6460 5704
rect 6367 5664 6460 5692
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 4154 5556 4160 5568
rect 4115 5528 4160 5556
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 6472 5556 6500 5652
rect 7650 5584 7656 5636
rect 7708 5624 7714 5636
rect 7837 5627 7895 5633
rect 7837 5624 7849 5627
rect 7708 5596 7849 5624
rect 7708 5584 7714 5596
rect 7837 5593 7849 5596
rect 7883 5593 7895 5627
rect 7944 5624 7972 5732
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8496 5701 8524 5732
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8588 5624 8616 5800
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 9941 5837 9947 5840
rect 9933 5831 9947 5837
rect 9933 5828 9945 5831
rect 9902 5800 9945 5828
rect 9933 5797 9945 5800
rect 9933 5791 9947 5797
rect 9941 5788 9947 5791
rect 9999 5788 10005 5840
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 13078 5828 13084 5840
rect 11940 5800 13084 5828
rect 11940 5788 11946 5800
rect 9766 5760 9772 5772
rect 9416 5732 9772 5760
rect 9416 5704 9444 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 11146 5720 11152 5772
rect 11204 5720 11210 5772
rect 11238 5720 11244 5772
rect 11296 5760 11302 5772
rect 12636 5769 12664 5800
rect 13078 5788 13084 5800
rect 13136 5788 13142 5840
rect 15749 5831 15807 5837
rect 15749 5797 15761 5831
rect 15795 5828 15807 5831
rect 17865 5831 17923 5837
rect 17865 5828 17877 5831
rect 15795 5800 17877 5828
rect 15795 5797 15807 5800
rect 15749 5791 15807 5797
rect 17865 5797 17877 5800
rect 17911 5797 17923 5831
rect 17865 5791 17923 5797
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11296 5732 11529 5760
rect 11296 5720 11302 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 12621 5763 12679 5769
rect 12621 5729 12633 5763
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 12888 5763 12946 5769
rect 12888 5729 12900 5763
rect 12934 5760 12946 5763
rect 14550 5760 14556 5772
rect 12934 5732 14412 5760
rect 14463 5732 14556 5760
rect 12934 5729 12946 5732
rect 12888 5723 12946 5729
rect 9398 5692 9404 5704
rect 9311 5664 9404 5692
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 11164 5692 11192 5720
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11164 5664 11621 5692
rect 9677 5655 9735 5661
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 11793 5695 11851 5701
rect 11793 5661 11805 5695
rect 11839 5692 11851 5695
rect 11974 5692 11980 5704
rect 11839 5664 11980 5692
rect 11839 5661 11851 5664
rect 11793 5655 11851 5661
rect 7944 5596 8616 5624
rect 7837 5587 7895 5593
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 9692 5624 9720 5655
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 14384 5636 14412 5732
rect 14550 5720 14556 5732
rect 14608 5760 14614 5772
rect 14921 5763 14979 5769
rect 14921 5760 14933 5763
rect 14608 5732 14933 5760
rect 14608 5720 14614 5732
rect 14921 5729 14933 5732
rect 14967 5729 14979 5763
rect 14921 5723 14979 5729
rect 16292 5763 16350 5769
rect 16292 5729 16304 5763
rect 16338 5760 16350 5763
rect 16338 5732 17080 5760
rect 16338 5729 16350 5732
rect 16292 5723 16350 5729
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 9364 5596 9720 5624
rect 11149 5627 11207 5633
rect 9364 5584 9370 5596
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 11422 5624 11428 5636
rect 11195 5596 11428 5624
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 14660 5624 14688 5655
rect 15470 5652 15476 5704
rect 15528 5692 15534 5704
rect 16022 5692 16028 5704
rect 15528 5664 16028 5692
rect 15528 5652 15534 5664
rect 16022 5652 16028 5664
rect 16080 5652 16086 5704
rect 17052 5636 17080 5732
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 14424 5596 14688 5624
rect 14424 5584 14430 5596
rect 17034 5584 17040 5636
rect 17092 5624 17098 5636
rect 18064 5624 18092 5655
rect 17092 5596 18092 5624
rect 17092 5584 17098 5596
rect 6730 5556 6736 5568
rect 6472 5528 6736 5556
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7742 5556 7748 5568
rect 7156 5528 7748 5556
rect 7156 5516 7162 5528
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 12434 5556 12440 5568
rect 8803 5528 12440 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 13998 5556 14004 5568
rect 13911 5528 14004 5556
rect 13998 5516 14004 5528
rect 14056 5556 14062 5568
rect 14642 5556 14648 5568
rect 14056 5528 14648 5556
rect 14056 5516 14062 5528
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 17494 5556 17500 5568
rect 17455 5528 17500 5556
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5352 3755 5355
rect 3786 5352 3792 5364
rect 3743 5324 3792 5352
rect 3743 5321 3755 5324
rect 3697 5315 3755 5321
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 4798 5352 4804 5364
rect 4663 5324 4804 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4798 5312 4804 5324
rect 4856 5312 4862 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 5994 5352 6000 5364
rect 5951 5324 6000 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7650 5352 7656 5364
rect 6972 5324 7656 5352
rect 6972 5312 6978 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8202 5312 8208 5364
rect 8260 5352 8266 5364
rect 8849 5355 8907 5361
rect 8849 5352 8861 5355
rect 8260 5324 8861 5352
rect 8260 5312 8266 5324
rect 8849 5321 8861 5324
rect 8895 5321 8907 5355
rect 11146 5352 11152 5364
rect 11107 5324 11152 5352
rect 8849 5315 8907 5321
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11974 5352 11980 5364
rect 11256 5324 11980 5352
rect 3970 5244 3976 5296
rect 4028 5284 4034 5296
rect 6362 5284 6368 5296
rect 4028 5256 6368 5284
rect 4028 5244 4034 5256
rect 6362 5244 6368 5256
rect 6420 5244 6426 5296
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 8941 5287 8999 5293
rect 8941 5284 8953 5287
rect 8536 5256 8953 5284
rect 8536 5244 8542 5256
rect 8941 5253 8953 5256
rect 8987 5253 8999 5287
rect 8941 5247 8999 5253
rect 10321 5287 10379 5293
rect 10321 5253 10333 5287
rect 10367 5284 10379 5287
rect 10410 5284 10416 5296
rect 10367 5256 10416 5284
rect 10367 5253 10379 5256
rect 10321 5247 10379 5253
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4120 5188 4261 5216
rect 4120 5176 4126 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 5258 5216 5264 5228
rect 5219 5188 5264 5216
rect 4249 5179 4307 5185
rect 5258 5176 5264 5188
rect 5316 5176 5322 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6914 5216 6920 5228
rect 6595 5188 6920 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 8956 5216 8984 5247
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 11256 5284 11284 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 14090 5352 14096 5364
rect 13096 5324 14096 5352
rect 13096 5284 13124 5324
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 16853 5355 16911 5361
rect 14240 5324 16804 5352
rect 14240 5312 14246 5324
rect 10980 5256 11284 5284
rect 11624 5256 13124 5284
rect 16776 5284 16804 5324
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 17034 5352 17040 5364
rect 16899 5324 17040 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 17770 5352 17776 5364
rect 17731 5324 17776 5352
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 18138 5284 18144 5296
rect 16776 5256 18144 5284
rect 9674 5216 9680 5228
rect 8956 5188 9680 5216
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 10980 5225 11008 5256
rect 11624 5225 11652 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 10965 5219 11023 5225
rect 10965 5185 10977 5219
rect 11011 5185 11023 5219
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 10965 5179 11023 5185
rect 11072 5188 11621 5216
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2124 5151 2182 5157
rect 2124 5117 2136 5151
rect 2170 5148 2182 5151
rect 2682 5148 2688 5160
rect 2170 5120 2688 5148
rect 2170 5117 2182 5120
rect 2124 5111 2182 5117
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6638 5148 6644 5160
rect 5859 5120 6644 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 6730 5108 6736 5160
rect 6788 5148 6794 5160
rect 7282 5148 7288 5160
rect 6788 5120 7288 5148
rect 6788 5108 6794 5120
rect 7282 5108 7288 5120
rect 7340 5148 7346 5160
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 7340 5120 7481 5148
rect 7340 5108 7346 5120
rect 7469 5117 7481 5120
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7736 5151 7794 5157
rect 7736 5117 7748 5151
rect 7782 5148 7794 5151
rect 9398 5148 9404 5160
rect 7782 5120 9404 5148
rect 7782 5117 7794 5120
rect 7736 5111 7794 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 11072 5148 11100 5188
rect 11609 5185 11621 5188
rect 11655 5185 11667 5219
rect 11790 5216 11796 5228
rect 11751 5188 11796 5216
rect 11609 5179 11667 5185
rect 11790 5176 11796 5188
rect 11848 5176 11854 5228
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 15105 5219 15163 5225
rect 15105 5216 15117 5219
rect 14700 5188 15117 5216
rect 14700 5176 14706 5188
rect 15105 5185 15117 5188
rect 15151 5185 15163 5219
rect 15470 5216 15476 5228
rect 15431 5188 15476 5216
rect 15105 5179 15163 5185
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 16666 5176 16672 5228
rect 16724 5216 16730 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 16724 5188 17509 5216
rect 16724 5176 16730 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 13078 5148 13084 5160
rect 9968 5120 11100 5148
rect 13039 5120 13084 5148
rect 2958 5040 2964 5092
rect 3016 5080 3022 5092
rect 3513 5083 3571 5089
rect 3513 5080 3525 5083
rect 3016 5052 3525 5080
rect 3016 5040 3022 5052
rect 3513 5049 3525 5052
rect 3559 5080 3571 5083
rect 4157 5083 4215 5089
rect 4157 5080 4169 5083
rect 3559 5052 4169 5080
rect 3559 5049 3571 5052
rect 3513 5043 3571 5049
rect 4157 5049 4169 5052
rect 4203 5080 4215 5083
rect 5629 5083 5687 5089
rect 5629 5080 5641 5083
rect 4203 5052 5641 5080
rect 4203 5049 4215 5052
rect 4157 5043 4215 5049
rect 5629 5049 5641 5052
rect 5675 5049 5687 5083
rect 5629 5043 5687 5049
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 3237 5015 3295 5021
rect 3237 5012 3249 5015
rect 3108 4984 3249 5012
rect 3108 4972 3114 4984
rect 3237 4981 3249 4984
rect 3283 4981 3295 5015
rect 3237 4975 3295 4981
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 3694 5012 3700 5024
rect 3467 4984 3700 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 3694 4972 3700 4984
rect 3752 5012 3758 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 3752 4984 4077 5012
rect 3752 4972 3758 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 4065 4975 4123 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5534 5012 5540 5024
rect 5123 4984 5540 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 5644 5012 5672 5043
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 9968 5089 9996 5120
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13170 5108 13176 5160
rect 13228 5148 13234 5160
rect 14921 5151 14979 5157
rect 14921 5148 14933 5151
rect 13228 5120 14933 5148
rect 13228 5108 13234 5120
rect 14921 5117 14933 5120
rect 14967 5117 14979 5151
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 14921 5111 14979 5117
rect 15580 5120 19073 5148
rect 9953 5083 10011 5089
rect 9953 5080 9965 5083
rect 6880 5052 9965 5080
rect 6880 5040 6886 5052
rect 9953 5049 9965 5052
rect 9999 5049 10011 5083
rect 9953 5043 10011 5049
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 11054 5080 11060 5092
rect 10468 5052 11060 5080
rect 10468 5040 10474 5052
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 13348 5083 13406 5089
rect 11563 5052 12296 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 12268 5024 12296 5052
rect 13348 5049 13360 5083
rect 13394 5080 13406 5083
rect 13394 5052 13676 5080
rect 13394 5049 13406 5052
rect 13348 5043 13406 5049
rect 6270 5012 6276 5024
rect 5644 4984 6276 5012
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 6638 5012 6644 5024
rect 6411 4984 6644 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 8938 5012 8944 5024
rect 6788 4984 8944 5012
rect 6788 4972 6794 4984
rect 8938 4972 8944 4984
rect 8996 5012 9002 5024
rect 9582 5012 9588 5024
rect 8996 4984 9588 5012
rect 8996 4972 9002 4984
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 10100 4984 10149 5012
rect 10100 4972 10106 4984
rect 10137 4981 10149 4984
rect 10183 5012 10195 5015
rect 10689 5015 10747 5021
rect 10689 5012 10701 5015
rect 10183 4984 10701 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10689 4981 10701 4984
rect 10735 4981 10747 5015
rect 10689 4975 10747 4981
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 11146 5012 11152 5024
rect 10827 4984 11152 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 11977 5015 12035 5021
rect 11977 5012 11989 5015
rect 11940 4984 11989 5012
rect 11940 4972 11946 4984
rect 11977 4981 11989 4984
rect 12023 4981 12035 5015
rect 12250 5012 12256 5024
rect 12163 4984 12256 5012
rect 11977 4975 12035 4981
rect 12250 4972 12256 4984
rect 12308 5012 12314 5024
rect 13538 5012 13544 5024
rect 12308 4984 13544 5012
rect 12308 4972 12314 4984
rect 13538 4972 13544 4984
rect 13596 4972 13602 5024
rect 13648 5012 13676 5052
rect 13722 5040 13728 5092
rect 13780 5080 13786 5092
rect 15013 5083 15071 5089
rect 15013 5080 15025 5083
rect 13780 5052 15025 5080
rect 13780 5040 13786 5052
rect 15013 5049 15025 5052
rect 15059 5049 15071 5083
rect 15013 5043 15071 5049
rect 15194 5040 15200 5092
rect 15252 5080 15258 5092
rect 15580 5080 15608 5120
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 15746 5089 15752 5092
rect 15740 5080 15752 5089
rect 15252 5052 15608 5080
rect 15707 5052 15752 5080
rect 15252 5040 15258 5052
rect 15740 5043 15752 5052
rect 15804 5080 15810 5092
rect 16666 5080 16672 5092
rect 15804 5052 16672 5080
rect 15746 5040 15752 5043
rect 15804 5040 15810 5052
rect 16666 5040 16672 5052
rect 16724 5040 16730 5092
rect 17313 5083 17371 5089
rect 17313 5049 17325 5083
rect 17359 5080 17371 5083
rect 17770 5080 17776 5092
rect 17359 5052 17776 5080
rect 17359 5049 17371 5052
rect 17313 5043 17371 5049
rect 17770 5040 17776 5052
rect 17828 5040 17834 5092
rect 19337 5083 19395 5089
rect 19337 5049 19349 5083
rect 19383 5080 19395 5083
rect 19978 5080 19984 5092
rect 19383 5052 19984 5080
rect 19383 5049 19395 5052
rect 19337 5043 19395 5049
rect 19978 5040 19984 5052
rect 20036 5040 20042 5092
rect 13998 5012 14004 5024
rect 13648 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14458 5012 14464 5024
rect 14419 4984 14464 5012
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 16942 5012 16948 5024
rect 14608 4984 14653 5012
rect 16903 4984 16948 5012
rect 14608 4972 14614 4984
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17405 5015 17463 5021
rect 17405 5012 17417 5015
rect 17276 4984 17417 5012
rect 17276 4972 17282 4984
rect 17405 4981 17417 4984
rect 17451 5012 17463 5015
rect 18049 5015 18107 5021
rect 18049 5012 18061 5015
rect 17451 4984 18061 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 18049 4981 18061 4984
rect 18095 4981 18107 5015
rect 18049 4975 18107 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4777 2099 4811
rect 3418 4808 3424 4820
rect 3379 4780 3424 4808
rect 2041 4771 2099 4777
rect 1670 4700 1676 4752
rect 1728 4740 1734 4752
rect 1765 4743 1823 4749
rect 1765 4740 1777 4743
rect 1728 4712 1777 4740
rect 1728 4700 1734 4712
rect 1765 4709 1777 4712
rect 1811 4709 1823 4743
rect 1765 4703 1823 4709
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4672 1547 4675
rect 2056 4672 2084 4771
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5997 4811 6055 4817
rect 5997 4808 6009 4811
rect 5316 4780 6009 4808
rect 5316 4768 5322 4780
rect 5997 4777 6009 4780
rect 6043 4777 6055 4811
rect 5997 4771 6055 4777
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 7374 4808 7380 4820
rect 7331 4780 7380 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 8113 4811 8171 4817
rect 8113 4777 8125 4811
rect 8159 4808 8171 4811
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 8159 4780 10333 4808
rect 8159 4777 8171 4780
rect 8113 4771 8171 4777
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 10321 4771 10379 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 12437 4811 12495 4817
rect 12437 4808 12449 4811
rect 11940 4780 12449 4808
rect 11940 4768 11946 4780
rect 12437 4777 12449 4780
rect 12483 4777 12495 4811
rect 12437 4771 12495 4777
rect 12897 4811 12955 4817
rect 12897 4777 12909 4811
rect 12943 4808 12955 4811
rect 13170 4808 13176 4820
rect 12943 4780 13176 4808
rect 12943 4777 12955 4780
rect 12897 4771 12955 4777
rect 13170 4768 13176 4780
rect 13228 4768 13234 4820
rect 13722 4808 13728 4820
rect 13683 4780 13728 4808
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 15194 4808 15200 4820
rect 14476 4780 15200 4808
rect 3326 4740 3332 4752
rect 3287 4712 3332 4740
rect 3326 4700 3332 4712
rect 3384 4700 3390 4752
rect 14476 4740 14504 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15344 4780 15669 4808
rect 15344 4768 15350 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 16117 4811 16175 4817
rect 16117 4777 16129 4811
rect 16163 4777 16175 4811
rect 16117 4771 16175 4777
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 16942 4808 16948 4820
rect 16623 4780 16948 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 4540 4712 14504 4740
rect 1535 4644 2084 4672
rect 2409 4675 2467 4681
rect 1535 4641 1547 4644
rect 1489 4635 1547 4641
rect 2409 4641 2421 4675
rect 2455 4641 2467 4675
rect 2409 4635 2467 4641
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 3142 4672 3148 4684
rect 2547 4644 3148 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 1394 4564 1400 4616
rect 1452 4604 1458 4616
rect 2424 4604 2452 4635
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 1452 4576 2452 4604
rect 2685 4607 2743 4613
rect 1452 4564 1458 4576
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 2774 4604 2780 4616
rect 2731 4576 2780 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 3602 4604 3608 4616
rect 3563 4576 3608 4604
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 4540 4536 4568 4712
rect 14550 4700 14556 4752
rect 14608 4740 14614 4752
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 14608 4712 15761 4740
rect 14608 4700 14614 4712
rect 15749 4709 15761 4712
rect 15795 4709 15807 4743
rect 16132 4740 16160 4771
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17313 4811 17371 4817
rect 17313 4777 17325 4811
rect 17359 4808 17371 4811
rect 17494 4808 17500 4820
rect 17359 4780 17500 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 17405 4743 17463 4749
rect 17405 4740 17417 4743
rect 16132 4712 17417 4740
rect 15749 4703 15807 4709
rect 17405 4709 17417 4712
rect 17451 4709 17463 4743
rect 17405 4703 17463 4709
rect 4617 4675 4675 4681
rect 4617 4641 4629 4675
rect 4663 4672 4675 4675
rect 4706 4672 4712 4684
rect 4663 4644 4712 4672
rect 4663 4641 4675 4644
rect 4617 4635 4675 4641
rect 4706 4632 4712 4644
rect 4764 4632 4770 4684
rect 4884 4675 4942 4681
rect 4884 4641 4896 4675
rect 4930 4672 4942 4675
rect 5442 4672 5448 4684
rect 4930 4644 5448 4672
rect 4930 4641 4942 4644
rect 4884 4635 4942 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7650 4672 7656 4684
rect 6972 4644 7656 4672
rect 6972 4632 6978 4644
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8478 4672 8484 4684
rect 8439 4644 8484 4672
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10778 4672 10784 4684
rect 10336 4644 10784 4672
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7064 4576 7757 4604
rect 7064 4564 7070 4576
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4604 7987 4607
rect 8202 4604 8208 4616
rect 7975 4576 8208 4604
rect 7975 4573 7987 4576
rect 7929 4567 7987 4573
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8570 4604 8576 4616
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 8754 4604 8760 4616
rect 8715 4576 8760 4604
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 10336 4604 10364 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 11112 4644 11621 4672
rect 11112 4632 11118 4644
rect 11609 4641 11621 4644
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4672 11759 4675
rect 11974 4672 11980 4684
rect 11747 4644 11980 4672
rect 11747 4641 11759 4644
rect 11701 4635 11759 4641
rect 9784 4576 10364 4604
rect 3007 4508 4568 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 6178 4496 6184 4548
rect 6236 4536 6242 4548
rect 9214 4536 9220 4548
rect 6236 4508 9220 4536
rect 6236 4496 6242 4508
rect 9214 4496 9220 4508
rect 9272 4496 9278 4548
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 6914 4468 6920 4480
rect 4212 4440 6920 4468
rect 4212 4428 4218 4440
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7101 4471 7159 4477
rect 7101 4468 7113 4471
rect 7064 4440 7113 4468
rect 7064 4428 7070 4440
rect 7101 4437 7113 4440
rect 7147 4468 7159 4471
rect 9784 4468 9812 4576
rect 10410 4564 10416 4616
rect 10468 4604 10474 4616
rect 10468 4576 10513 4604
rect 10468 4564 10474 4576
rect 9861 4539 9919 4545
rect 9861 4505 9873 4539
rect 9907 4536 9919 4539
rect 11624 4536 11652 4635
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13630 4632 13636 4684
rect 13688 4672 13694 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13688 4644 14105 4672
rect 13688 4632 13694 4644
rect 14093 4641 14105 4644
rect 14139 4672 14151 4675
rect 14274 4672 14280 4684
rect 14139 4644 14280 4672
rect 14139 4641 14151 4644
rect 14093 4635 14151 4641
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 14467 4644 16497 4672
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 11848 4576 11893 4604
rect 11992 4576 12541 4604
rect 11848 4564 11854 4576
rect 11992 4536 12020 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12529 4567 12587 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 12860 4576 13369 4604
rect 12860 4564 12866 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 13357 4567 13415 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13814 4604 13820 4616
rect 13587 4576 13820 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14182 4604 14188 4616
rect 14143 4576 14188 4604
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 9907 4508 11192 4536
rect 11624 4508 12020 4536
rect 12069 4539 12127 4545
rect 9907 4505 9919 4508
rect 9861 4499 9919 4505
rect 7147 4440 9812 4468
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 10134 4428 10140 4480
rect 10192 4468 10198 4480
rect 10781 4471 10839 4477
rect 10781 4468 10793 4471
rect 10192 4440 10793 4468
rect 10192 4428 10198 4440
rect 10781 4437 10793 4440
rect 10827 4437 10839 4471
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 10781 4431 10839 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11164 4468 11192 4508
rect 12069 4505 12081 4539
rect 12115 4536 12127 4539
rect 14467 4536 14495 4644
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 19978 4672 19984 4684
rect 19939 4644 19984 4672
rect 16485 4635 16543 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 14550 4564 14556 4616
rect 14608 4604 14614 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 14608 4576 15853 4604
rect 14608 4564 14614 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4604 16819 4607
rect 17034 4604 17040 4616
rect 16807 4576 17040 4604
rect 16807 4573 16819 4576
rect 16761 4567 16819 4573
rect 17034 4564 17040 4576
rect 17092 4564 17098 4616
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 15746 4536 15752 4548
rect 12115 4508 14495 4536
rect 14568 4508 15752 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 12710 4468 12716 4480
rect 11164 4440 12716 4468
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 12894 4428 12900 4480
rect 12952 4468 12958 4480
rect 14568 4468 14596 4508
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 12952 4440 14596 4468
rect 14645 4471 14703 4477
rect 12952 4428 12958 4440
rect 14645 4437 14657 4471
rect 14691 4468 14703 4471
rect 15010 4468 15016 4480
rect 14691 4440 15016 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 15010 4428 15016 4440
rect 15068 4428 15074 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 16945 4471 17003 4477
rect 16945 4437 16957 4471
rect 16991 4468 17003 4471
rect 17126 4468 17132 4480
rect 16991 4440 17132 4468
rect 16991 4437 17003 4440
rect 16945 4431 17003 4437
rect 17126 4428 17132 4440
rect 17184 4428 17190 4480
rect 20165 4471 20223 4477
rect 20165 4437 20177 4471
rect 20211 4468 20223 4471
rect 20806 4468 20812 4480
rect 20211 4440 20812 4468
rect 20211 4437 20223 4440
rect 20165 4431 20223 4437
rect 20806 4428 20812 4440
rect 20864 4428 20870 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 2832 4236 3249 4264
rect 2832 4224 2838 4236
rect 3237 4233 3249 4236
rect 3283 4233 3295 4267
rect 3237 4227 3295 4233
rect 3252 4128 3280 4227
rect 4062 4224 4068 4276
rect 4120 4264 4126 4276
rect 6178 4264 6184 4276
rect 4120 4236 6184 4264
rect 4120 4224 4126 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6328 4236 6837 4264
rect 6328 4224 6334 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 4798 4156 4804 4208
rect 4856 4196 4862 4208
rect 5074 4196 5080 4208
rect 4856 4168 5080 4196
rect 4856 4156 4862 4168
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 5534 4156 5540 4208
rect 5592 4196 5598 4208
rect 6840 4196 6868 4227
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7193 4267 7251 4273
rect 7193 4264 7205 4267
rect 6972 4236 7205 4264
rect 6972 4224 6978 4236
rect 7193 4233 7205 4236
rect 7239 4233 7251 4267
rect 7193 4227 7251 4233
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 8478 4264 8484 4276
rect 8435 4236 8484 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 8478 4224 8484 4236
rect 8536 4224 8542 4276
rect 10137 4267 10195 4273
rect 10137 4233 10149 4267
rect 10183 4264 10195 4267
rect 10226 4264 10232 4276
rect 10183 4236 10232 4264
rect 10183 4233 10195 4236
rect 10137 4227 10195 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 11146 4264 11152 4276
rect 11107 4236 11152 4264
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11348 4236 11989 4264
rect 5592 4168 6776 4196
rect 6840 4168 6960 4196
rect 5592 4156 5598 4168
rect 3252 4100 3464 4128
rect 1854 4060 1860 4072
rect 1767 4032 1860 4060
rect 1854 4020 1860 4032
rect 1912 4060 1918 4072
rect 3326 4060 3332 4072
rect 1912 4032 3332 4060
rect 1912 4020 1918 4032
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3436 4060 3464 4100
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 4764 4100 6101 4128
rect 4764 4088 4770 4100
rect 6089 4097 6101 4100
rect 6135 4128 6147 4131
rect 6178 4128 6184 4140
rect 6135 4100 6184 4128
rect 6135 4097 6147 4100
rect 6089 4091 6147 4097
rect 6178 4088 6184 4100
rect 6236 4088 6242 4140
rect 6748 4128 6776 4168
rect 6932 4140 6960 4168
rect 8220 4168 8708 4196
rect 8220 4140 8248 4168
rect 6822 4128 6828 4140
rect 6748 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6914 4088 6920 4140
rect 6972 4088 6978 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 7024 4100 8033 4128
rect 3585 4063 3643 4069
rect 3585 4060 3597 4063
rect 3436 4032 3597 4060
rect 3585 4029 3597 4032
rect 3631 4029 3643 4063
rect 3585 4023 3643 4029
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 5353 4063 5411 4069
rect 5353 4060 5365 4063
rect 4120 4032 5365 4060
rect 4120 4020 4126 4032
rect 5353 4029 5365 4032
rect 5399 4060 5411 4063
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5399 4032 6009 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 5997 4029 6009 4032
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 2038 3952 2044 4004
rect 2096 4001 2102 4004
rect 2096 3995 2160 4001
rect 2096 3961 2114 3995
rect 2148 3961 2160 3995
rect 4154 3992 4160 4004
rect 2096 3955 2160 3961
rect 2424 3964 4160 3992
rect 2096 3952 2102 3955
rect 1118 3884 1124 3936
rect 1176 3924 1182 3936
rect 2424 3924 2452 3964
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 7024 4001 7052 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8202 4128 8208 4140
rect 8115 4100 8208 4128
rect 8021 4091 8079 4097
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7156 4032 7941 4060
rect 7156 4020 7162 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 8036 4060 8064 4091
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8680 4128 8708 4168
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 8812 4168 10732 4196
rect 8812 4156 8818 4168
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8680 4100 9045 4128
rect 9033 4097 9045 4100
rect 9079 4128 9091 4131
rect 9122 4128 9128 4140
rect 9079 4100 9128 4128
rect 9079 4097 9091 4100
rect 9033 4091 9091 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 10134 4128 10140 4140
rect 9324 4100 10140 4128
rect 9324 4060 9352 4100
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 10594 4128 10600 4140
rect 10555 4100 10600 4128
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 10704 4137 10732 4168
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11348 4196 11376 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 13630 4264 13636 4276
rect 11977 4227 12035 4233
rect 12176 4236 13636 4264
rect 11790 4196 11796 4208
rect 11112 4168 11376 4196
rect 11716 4168 11796 4196
rect 11112 4156 11118 4168
rect 11716 4137 11744 4168
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 8036 4032 9352 4060
rect 7929 4023 7987 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 11057 4063 11115 4069
rect 11057 4060 11069 4063
rect 9456 4032 11069 4060
rect 9456 4020 9462 4032
rect 11057 4029 11069 4032
rect 11103 4060 11115 4063
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11103 4032 11621 4060
rect 11103 4029 11115 4032
rect 11057 4023 11115 4029
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 7009 3995 7067 4001
rect 7009 3992 7021 3995
rect 4540 3964 7021 3992
rect 1176 3896 2452 3924
rect 1176 3884 1182 3896
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 4540 3924 4568 3964
rect 7009 3961 7021 3964
rect 7055 3961 7067 3995
rect 8570 3992 8576 4004
rect 7009 3955 7067 3961
rect 7576 3964 8576 3992
rect 4706 3924 4712 3936
rect 2556 3896 4568 3924
rect 4667 3896 4712 3924
rect 2556 3884 2562 3896
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6362 3924 6368 3936
rect 6052 3896 6368 3924
rect 6052 3884 6058 3896
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 6604 3896 7389 3924
rect 6604 3884 6610 3896
rect 7377 3893 7389 3896
rect 7423 3924 7435 3927
rect 7466 3924 7472 3936
rect 7423 3896 7472 3924
rect 7423 3893 7435 3896
rect 7377 3887 7435 3893
rect 7466 3884 7472 3896
rect 7524 3884 7530 3936
rect 7576 3933 7604 3964
rect 8570 3952 8576 3964
rect 8628 3952 8634 4004
rect 8849 3995 8907 4001
rect 8849 3992 8861 3995
rect 8680 3964 8861 3992
rect 7561 3927 7619 3933
rect 7561 3893 7573 3927
rect 7607 3893 7619 3927
rect 7561 3887 7619 3893
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 8680 3924 8708 3964
rect 8849 3961 8861 3964
rect 8895 3992 8907 3995
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 8895 3964 9229 3992
rect 8895 3961 8907 3964
rect 8849 3955 8907 3961
rect 9217 3961 9229 3964
rect 9263 3992 9275 3995
rect 10042 3992 10048 4004
rect 9263 3964 10048 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 10042 3952 10048 3964
rect 10100 3952 10106 4004
rect 10134 3952 10140 4004
rect 10192 3992 10198 4004
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 10192 3964 11529 3992
rect 10192 3952 10198 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 11624 3992 11652 4023
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12176 4069 12204 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 14366 4264 14372 4276
rect 13872 4236 14372 4264
rect 13872 4224 13878 4236
rect 14366 4224 14372 4236
rect 14424 4264 14430 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14424 4236 15025 4264
rect 14424 4224 14430 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 12250 4156 12256 4208
rect 12308 4196 12314 4208
rect 12621 4199 12679 4205
rect 12621 4196 12633 4199
rect 12308 4168 12633 4196
rect 12308 4156 12314 4168
rect 12621 4165 12633 4168
rect 12667 4196 12679 4199
rect 13262 4196 13268 4208
rect 12667 4168 13268 4196
rect 12667 4165 12679 4168
rect 12621 4159 12679 4165
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 12802 4128 12808 4140
rect 12763 4100 12808 4128
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 15010 4088 15016 4140
rect 15068 4128 15074 4140
rect 22646 4128 22652 4140
rect 15068 4100 22652 4128
rect 15068 4088 15074 4100
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 12032 4032 12173 4060
rect 12032 4020 12038 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 13630 4060 13636 4072
rect 13591 4032 13636 4060
rect 12161 4023 12219 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 12802 3992 12808 4004
rect 11624 3964 12808 3992
rect 11517 3955 11575 3961
rect 8536 3896 8708 3924
rect 8757 3927 8815 3933
rect 8536 3884 8542 3896
rect 8757 3893 8769 3927
rect 8803 3924 8815 3927
rect 8938 3924 8944 3936
rect 8803 3896 8944 3924
rect 8803 3893 8815 3896
rect 8757 3887 8815 3893
rect 8938 3884 8944 3896
rect 8996 3924 9002 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 8996 3896 9413 3924
rect 8996 3884 9002 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10870 3924 10876 3936
rect 10551 3896 10876 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11532 3924 11560 3955
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 13906 4001 13912 4004
rect 13900 3992 13912 4001
rect 13867 3964 13912 3992
rect 13900 3955 13912 3964
rect 13906 3952 13912 3955
rect 13964 3952 13970 4004
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 15028 3992 15056 4088
rect 17126 4060 17132 4072
rect 17087 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 14332 3964 15056 3992
rect 17405 3995 17463 4001
rect 14332 3952 14338 3964
rect 17405 3961 17417 3995
rect 17451 3992 17463 3995
rect 18046 3992 18052 4004
rect 17451 3964 18052 3992
rect 17451 3961 17463 3964
rect 17405 3955 17463 3961
rect 18046 3952 18052 3964
rect 18104 3952 18110 4004
rect 11882 3924 11888 3936
rect 11532 3896 11888 3924
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 13814 3924 13820 3936
rect 12308 3896 13820 3924
rect 12308 3884 12314 3896
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 198 3680 204 3732
rect 256 3720 262 3732
rect 2774 3720 2780 3732
rect 256 3692 2780 3720
rect 256 3680 262 3692
rect 2774 3680 2780 3692
rect 2832 3680 2838 3732
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 3476 3692 5396 3720
rect 3476 3680 3482 3692
rect 1940 3655 1998 3661
rect 1940 3621 1952 3655
rect 1986 3652 1998 3655
rect 3050 3652 3056 3664
rect 1986 3624 3056 3652
rect 1986 3621 1998 3624
rect 1940 3615 1998 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 3326 3612 3332 3664
rect 3384 3652 3390 3664
rect 3384 3624 4568 3652
rect 3384 3612 3390 3624
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 1762 3584 1768 3596
rect 1719 3556 1768 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 3513 3587 3571 3593
rect 3513 3584 3525 3587
rect 2832 3556 3525 3584
rect 2832 3544 2838 3556
rect 3513 3553 3525 3556
rect 3559 3553 3571 3587
rect 3513 3547 3571 3553
rect 3602 3544 3608 3596
rect 3660 3584 3666 3596
rect 4540 3593 4568 3624
rect 4706 3612 4712 3664
rect 4764 3661 4770 3664
rect 4764 3655 4828 3661
rect 4764 3621 4782 3655
rect 4816 3621 4828 3655
rect 4764 3615 4828 3621
rect 4764 3612 4770 3615
rect 4890 3612 4896 3664
rect 4948 3612 4954 3664
rect 5368 3652 5396 3692
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5500 3692 5917 3720
rect 5500 3680 5506 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 5997 3723 6055 3729
rect 5997 3689 6009 3723
rect 6043 3720 6055 3723
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 6043 3692 7205 3720
rect 6043 3689 6055 3692
rect 5997 3683 6055 3689
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 7699 3692 8953 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 8941 3683 8999 3689
rect 5626 3652 5632 3664
rect 5368 3624 5632 3652
rect 5626 3612 5632 3624
rect 5684 3612 5690 3664
rect 5920 3652 5948 3683
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10042 3720 10048 3732
rect 9907 3692 10048 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 10321 3723 10379 3729
rect 10321 3689 10333 3723
rect 10367 3720 10379 3723
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10367 3692 10701 3720
rect 10367 3689 10379 3692
rect 10321 3683 10379 3689
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11517 3723 11575 3729
rect 11517 3720 11529 3723
rect 10928 3692 11529 3720
rect 10928 3680 10934 3692
rect 11517 3689 11529 3692
rect 11563 3689 11575 3723
rect 13078 3720 13084 3732
rect 11517 3683 11575 3689
rect 12084 3692 13084 3720
rect 5920 3624 7236 3652
rect 4525 3587 4583 3593
rect 3660 3556 3705 3584
rect 3660 3544 3666 3556
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4908 3584 4936 3612
rect 6362 3584 6368 3596
rect 4571 3556 4936 3584
rect 6323 3556 6368 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 6730 3584 6736 3596
rect 6503 3556 6736 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7208 3584 7236 3624
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 8110 3652 8116 3664
rect 7524 3624 8116 3652
rect 7524 3612 7530 3624
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 10134 3652 10140 3664
rect 8220 3624 10140 3652
rect 7208 3556 7420 3584
rect 7392 3525 7420 3556
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8021 3587 8079 3593
rect 8021 3584 8033 3587
rect 7708 3556 8033 3584
rect 7708 3544 7714 3556
rect 8021 3553 8033 3556
rect 8067 3553 8079 3587
rect 8220 3584 8248 3624
rect 10134 3612 10140 3624
rect 10192 3612 10198 3664
rect 10229 3655 10287 3661
rect 10229 3621 10241 3655
rect 10275 3652 10287 3655
rect 10962 3652 10968 3664
rect 10275 3624 10968 3652
rect 10275 3621 10287 3624
rect 10229 3615 10287 3621
rect 10962 3612 10968 3624
rect 11020 3612 11026 3664
rect 8846 3584 8852 3596
rect 8021 3547 8079 3553
rect 8128 3556 8248 3584
rect 8807 3556 8852 3584
rect 3697 3519 3755 3525
rect 3697 3485 3709 3519
rect 3743 3485 3755 3519
rect 3697 3479 3755 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 7285 3519 7343 3525
rect 7285 3485 7297 3519
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 8128 3516 8156 3556
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9401 3587 9459 3593
rect 9401 3584 9413 3587
rect 8996 3556 9413 3584
rect 8996 3544 9002 3556
rect 9401 3553 9413 3556
rect 9447 3584 9459 3587
rect 11057 3587 11115 3593
rect 9447 3556 10272 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 7377 3479 7435 3485
rect 7944 3488 8156 3516
rect 3712 3448 3740 3479
rect 3068 3420 3740 3448
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 3068 3389 3096 3420
rect 6178 3408 6184 3460
rect 6236 3448 6242 3460
rect 6564 3448 6592 3479
rect 6822 3448 6828 3460
rect 6236 3420 6592 3448
rect 6783 3420 6828 3448
rect 6236 3408 6242 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7300 3448 7328 3479
rect 6972 3420 7328 3448
rect 6972 3408 6978 3420
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 2096 3352 3065 3380
rect 2096 3340 2102 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7944 3380 7972 3488
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8260 3488 8305 3516
rect 8260 3476 8266 3488
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9033 3519 9091 3525
rect 9033 3516 9045 3519
rect 8812 3488 9045 3516
rect 8812 3476 8818 3488
rect 9033 3485 9045 3488
rect 9079 3516 9091 3519
rect 10042 3516 10048 3528
rect 9079 3488 10048 3516
rect 9079 3485 9091 3488
rect 9033 3479 9091 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 8481 3451 8539 3457
rect 8481 3417 8493 3451
rect 8527 3448 8539 3451
rect 10134 3448 10140 3460
rect 8527 3420 10140 3448
rect 8527 3417 8539 3420
rect 8481 3411 8539 3417
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 10244 3448 10272 3556
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11422 3584 11428 3596
rect 11103 3556 11428 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11422 3544 11428 3556
rect 11480 3544 11486 3596
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10376 3488 10425 3516
rect 10376 3476 10382 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11698 3516 11704 3528
rect 11379 3488 11704 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11164 3448 11192 3479
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12084 3516 12112 3692
rect 13078 3680 13084 3692
rect 13136 3720 13142 3732
rect 13630 3720 13636 3732
rect 13136 3692 13636 3720
rect 13136 3680 13142 3692
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14182 3720 14188 3732
rect 13955 3692 14188 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 12161 3655 12219 3661
rect 12161 3621 12173 3655
rect 12207 3652 12219 3655
rect 15562 3652 15568 3664
rect 12207 3624 15568 3652
rect 12207 3621 12219 3624
rect 12161 3615 12219 3621
rect 15562 3612 15568 3624
rect 15620 3652 15626 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15620 3624 16037 3652
rect 15620 3612 15626 3624
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 16025 3615 16083 3621
rect 12517 3544 12523 3596
rect 12575 3584 12581 3596
rect 12575 3556 12620 3584
rect 12575 3544 12581 3556
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 15473 3587 15531 3593
rect 14332 3556 14377 3584
rect 14332 3544 14338 3556
rect 15473 3553 15485 3587
rect 15519 3584 15531 3587
rect 15654 3584 15660 3596
rect 15519 3556 15660 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 18046 3584 18052 3596
rect 18007 3556 18052 3584
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 12253 3519 12311 3525
rect 12253 3516 12265 3519
rect 11848 3488 12265 3516
rect 11848 3476 11854 3488
rect 12253 3485 12265 3488
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 13872 3488 14381 3516
rect 13872 3476 13878 3488
rect 14369 3485 14381 3488
rect 14415 3485 14427 3519
rect 14369 3479 14427 3485
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3485 14519 3519
rect 14461 3479 14519 3485
rect 15749 3519 15807 3525
rect 15749 3485 15761 3519
rect 15795 3516 15807 3519
rect 16390 3516 16396 3528
rect 15795 3488 16396 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 12161 3451 12219 3457
rect 12161 3448 12173 3451
rect 10244 3420 12173 3448
rect 12161 3417 12173 3420
rect 12207 3417 12219 3451
rect 12161 3411 12219 3417
rect 13633 3451 13691 3457
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 13906 3448 13912 3460
rect 13679 3420 13912 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 13906 3408 13912 3420
rect 13964 3448 13970 3460
rect 14476 3448 14504 3479
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 20162 3448 20168 3460
rect 13964 3420 14504 3448
rect 18156 3420 20168 3448
rect 13964 3408 13970 3420
rect 6788 3352 7972 3380
rect 6788 3340 6794 3352
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9766 3380 9772 3392
rect 8168 3352 9772 3380
rect 8168 3340 8174 3352
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 13354 3380 13360 3392
rect 11940 3352 13360 3380
rect 11940 3340 11946 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 13817 3383 13875 3389
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 13998 3380 14004 3392
rect 13863 3352 14004 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 13998 3340 14004 3352
rect 14056 3380 14062 3392
rect 14274 3380 14280 3392
rect 14056 3352 14280 3380
rect 14056 3340 14062 3352
rect 14274 3340 14280 3352
rect 14332 3380 14338 3392
rect 18156 3380 18184 3420
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 14332 3352 18184 3380
rect 18233 3383 18291 3389
rect 14332 3340 14338 3352
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18966 3380 18972 3392
rect 18279 3352 18972 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 18966 3340 18972 3352
rect 19024 3340 19030 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 3602 3176 3608 3188
rect 2832 3148 2877 3176
rect 3563 3148 3608 3176
rect 2832 3136 2838 3148
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3176 4767 3179
rect 4890 3176 4896 3188
rect 4755 3148 4896 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 7098 3176 7104 3188
rect 5000 3148 7104 3176
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 5000 3108 5028 3148
rect 7098 3136 7104 3148
rect 7156 3136 7162 3188
rect 8478 3176 8484 3188
rect 7576 3148 8484 3176
rect 5534 3108 5540 3120
rect 1728 3080 5028 3108
rect 5092 3080 5540 3108
rect 1728 3068 1734 3080
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 1636 3012 2421 3040
rect 1636 3000 1642 3012
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2682 3040 2688 3052
rect 2639 3012 2688 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2682 3000 2688 3012
rect 2740 3040 2746 3052
rect 3050 3040 3056 3052
rect 2740 3012 3056 3040
rect 2740 3000 2746 3012
rect 3050 3000 3056 3012
rect 3108 3040 3114 3052
rect 3329 3043 3387 3049
rect 3329 3040 3341 3043
rect 3108 3012 3341 3040
rect 3108 3000 3114 3012
rect 3329 3009 3341 3012
rect 3375 3040 3387 3043
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3375 3012 4169 3040
rect 3375 3009 3387 3012
rect 3329 3003 3387 3009
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 2317 2975 2375 2981
rect 2317 2972 2329 2975
rect 1544 2944 2329 2972
rect 1544 2932 1550 2944
rect 2317 2941 2329 2944
rect 2363 2941 2375 2975
rect 4246 2972 4252 2984
rect 2317 2935 2375 2941
rect 3160 2944 4252 2972
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 2590 2904 2596 2916
rect 1719 2876 2596 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 2590 2864 2596 2876
rect 2648 2864 2654 2916
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1946 2836 1952 2848
rect 1907 2808 1952 2836
rect 1946 2796 1952 2808
rect 2004 2796 2010 2848
rect 3050 2796 3056 2848
rect 3108 2836 3114 2848
rect 3160 2845 3188 2944
rect 4246 2932 4252 2944
rect 4304 2932 4310 2984
rect 5092 2981 5120 3080
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 7576 3108 7604 3148
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 8812 3148 8953 3176
rect 8812 3136 8818 3148
rect 8941 3145 8953 3148
rect 8987 3145 8999 3179
rect 9306 3176 9312 3188
rect 8941 3139 8999 3145
rect 9048 3148 9312 3176
rect 5960 3080 6408 3108
rect 5960 3068 5966 3080
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5442 3040 5448 3052
rect 5399 3012 5448 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 6086 3040 6092 3052
rect 6043 3012 6092 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6178 3000 6184 3052
rect 6236 3040 6242 3052
rect 6380 3049 6408 3080
rect 6932 3080 7604 3108
rect 6365 3043 6423 3049
rect 6236 3012 6281 3040
rect 6236 3000 6242 3012
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 5077 2975 5135 2981
rect 5077 2941 5089 2975
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 5169 2975 5227 2981
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5534 2972 5540 2984
rect 5215 2944 5540 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 6932 2972 6960 3080
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7340 3012 7573 3040
rect 7340 3000 7346 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 5684 2944 6960 2972
rect 7009 2975 7067 2981
rect 5684 2932 5690 2944
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7466 2972 7472 2984
rect 7055 2944 7472 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7828 2975 7886 2981
rect 7828 2972 7840 2975
rect 7760 2944 7840 2972
rect 7760 2916 7788 2944
rect 7828 2941 7840 2944
rect 7874 2972 7886 2975
rect 8202 2972 8208 2984
rect 7874 2944 8208 2972
rect 7874 2941 7886 2944
rect 7828 2935 7886 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8956 2972 8984 3139
rect 9048 3049 9076 3148
rect 9306 3136 9312 3148
rect 9364 3176 9370 3188
rect 10410 3176 10416 3188
rect 9364 3148 10272 3176
rect 10371 3148 10416 3176
rect 9364 3136 9370 3148
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3009 9091 3043
rect 10244 3040 10272 3148
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 11790 3176 11796 3188
rect 10520 3148 11796 3176
rect 10520 3049 10548 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12526 3176 12532 3188
rect 11931 3148 12532 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12526 3136 12532 3148
rect 12584 3176 12590 3188
rect 13814 3176 13820 3188
rect 12584 3148 12931 3176
rect 13775 3148 13820 3176
rect 12584 3136 12590 3148
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3077 12495 3111
rect 12437 3071 12495 3077
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10244 3012 10517 3040
rect 9033 3003 9091 3009
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 9289 2975 9347 2981
rect 9289 2972 9301 2975
rect 8956 2944 9301 2972
rect 9289 2941 9301 2944
rect 9335 2941 9347 2975
rect 9289 2935 9347 2941
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 12066 2972 12072 2984
rect 10100 2944 12072 2972
rect 10100 2932 10106 2944
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 12452 2972 12480 3071
rect 12903 3040 12931 3148
rect 13814 3136 13820 3148
rect 13872 3176 13878 3188
rect 18233 3179 18291 3185
rect 13872 3148 16068 3176
rect 13872 3136 13878 3148
rect 15286 3108 15292 3120
rect 14200 3080 15292 3108
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12903 3012 13001 3040
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13265 2975 13323 2981
rect 13265 2972 13277 2975
rect 12452 2944 13277 2972
rect 13265 2941 13277 2944
rect 13311 2941 13323 2975
rect 13265 2935 13323 2941
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14200 2972 14228 3080
rect 15286 3068 15292 3080
rect 15344 3068 15350 3120
rect 14277 3043 14335 3049
rect 14277 3009 14289 3043
rect 14323 3040 14335 3043
rect 14323 3012 14964 3040
rect 14323 3009 14335 3012
rect 14277 3003 14335 3009
rect 14047 2944 14228 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 14936 2981 14964 3012
rect 16040 2984 16068 3148
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 22186 3176 22192 3188
rect 18279 3148 22192 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 16209 3111 16267 3117
rect 16209 3077 16221 3111
rect 16255 3108 16267 3111
rect 16574 3108 16580 3120
rect 16255 3080 16580 3108
rect 16255 3077 16267 3080
rect 16209 3071 16267 3077
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 17405 3111 17463 3117
rect 17405 3077 17417 3111
rect 17451 3108 17463 3111
rect 17954 3108 17960 3120
rect 17451 3080 17960 3108
rect 17451 3077 17463 3080
rect 17405 3071 17463 3077
rect 17954 3068 17960 3080
rect 18012 3068 18018 3120
rect 18138 3068 18144 3120
rect 18196 3108 18202 3120
rect 18417 3111 18475 3117
rect 18417 3108 18429 3111
rect 18196 3080 18429 3108
rect 18196 3068 18202 3080
rect 18417 3077 18429 3080
rect 18463 3077 18475 3111
rect 18417 3071 18475 3077
rect 18785 3111 18843 3117
rect 18785 3077 18797 3111
rect 18831 3108 18843 3111
rect 19426 3108 19432 3120
rect 18831 3080 19432 3108
rect 18831 3077 18843 3080
rect 18785 3071 18843 3077
rect 19426 3068 19432 3080
rect 19484 3068 19490 3120
rect 19613 3111 19671 3117
rect 19613 3077 19625 3111
rect 19659 3108 19671 3111
rect 20346 3108 20352 3120
rect 19659 3080 20352 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 20346 3068 20352 3080
rect 20404 3068 20410 3120
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 16172 3012 19809 3040
rect 16172 3000 16178 3012
rect 14553 2975 14611 2981
rect 14553 2972 14565 2975
rect 14424 2944 14565 2972
rect 14424 2932 14430 2944
rect 14553 2941 14565 2944
rect 14599 2941 14611 2975
rect 14553 2935 14611 2941
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 15289 2975 15347 2981
rect 15289 2941 15301 2975
rect 15335 2972 15347 2975
rect 15378 2972 15384 2984
rect 15335 2944 15384 2972
rect 15335 2941 15347 2944
rect 15289 2935 15347 2941
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 15620 2944 15669 2972
rect 15620 2932 15626 2944
rect 15657 2941 15669 2944
rect 15703 2941 15715 2975
rect 16022 2972 16028 2984
rect 15935 2944 16028 2972
rect 15657 2935 15715 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16390 2972 16396 2984
rect 16351 2944 16396 2972
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 16758 2972 16764 2984
rect 16719 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 17218 2972 17224 2984
rect 17179 2944 17224 2972
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 17586 2972 17592 2984
rect 17368 2944 17592 2972
rect 17368 2932 17374 2944
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 17770 2932 17776 2984
rect 17828 2972 17834 2984
rect 18046 2972 18052 2984
rect 17828 2944 18052 2972
rect 17828 2932 17834 2944
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18601 2975 18659 2981
rect 18601 2972 18613 2975
rect 18196 2944 18613 2972
rect 18196 2932 18202 2944
rect 18601 2941 18613 2944
rect 18647 2941 18659 2975
rect 19058 2972 19064 2984
rect 19019 2944 19064 2972
rect 18601 2935 18659 2941
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19444 2981 19472 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 19797 3003 19855 3009
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2941 19487 2975
rect 20180 2972 20208 3000
rect 20349 2975 20407 2981
rect 20349 2972 20361 2975
rect 20180 2944 20361 2972
rect 19429 2935 19487 2941
rect 20349 2941 20361 2944
rect 20395 2941 20407 2975
rect 20349 2935 20407 2941
rect 3973 2907 4031 2913
rect 3973 2873 3985 2907
rect 4019 2904 4031 2907
rect 4338 2904 4344 2916
rect 4019 2876 4344 2904
rect 4019 2873 4031 2876
rect 3973 2867 4031 2873
rect 4338 2864 4344 2876
rect 4396 2904 4402 2916
rect 4433 2907 4491 2913
rect 4433 2904 4445 2907
rect 4396 2876 4445 2904
rect 4396 2864 4402 2876
rect 4433 2873 4445 2876
rect 4479 2873 4491 2907
rect 4433 2867 4491 2873
rect 5350 2864 5356 2916
rect 5408 2904 5414 2916
rect 5905 2907 5963 2913
rect 5905 2904 5917 2907
rect 5408 2876 5917 2904
rect 5408 2864 5414 2876
rect 5905 2873 5917 2876
rect 5951 2873 5963 2907
rect 5905 2867 5963 2873
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 6825 2907 6883 2913
rect 6825 2904 6837 2907
rect 6788 2876 6837 2904
rect 6788 2864 6794 2876
rect 6825 2873 6837 2876
rect 6871 2873 6883 2907
rect 6825 2867 6883 2873
rect 7285 2907 7343 2913
rect 7285 2873 7297 2907
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 3145 2839 3203 2845
rect 3145 2836 3157 2839
rect 3108 2808 3157 2836
rect 3108 2796 3114 2808
rect 3145 2805 3157 2808
rect 3191 2805 3203 2839
rect 3145 2799 3203 2805
rect 3237 2839 3295 2845
rect 3237 2805 3249 2839
rect 3283 2836 3295 2839
rect 3694 2836 3700 2848
rect 3283 2808 3700 2836
rect 3283 2805 3295 2808
rect 3237 2799 3295 2805
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 4065 2839 4123 2845
rect 4065 2805 4077 2839
rect 4111 2836 4123 2839
rect 4154 2836 4160 2848
rect 4111 2808 4160 2836
rect 4111 2805 4123 2808
rect 4065 2799 4123 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 6914 2836 6920 2848
rect 5583 2808 6920 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7300 2836 7328 2867
rect 7742 2864 7748 2916
rect 7800 2864 7806 2916
rect 8864 2876 9260 2904
rect 8864 2836 8892 2876
rect 7300 2808 8892 2836
rect 9232 2836 9260 2876
rect 10134 2864 10140 2916
rect 10192 2904 10198 2916
rect 10318 2904 10324 2916
rect 10192 2876 10324 2904
rect 10192 2864 10198 2876
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 10750 2907 10808 2913
rect 10750 2904 10762 2907
rect 10652 2876 10762 2904
rect 10652 2864 10658 2876
rect 10750 2873 10762 2876
rect 10796 2873 10808 2907
rect 10750 2867 10808 2873
rect 11146 2864 11152 2916
rect 11204 2904 11210 2916
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 11204 2876 12909 2904
rect 11204 2864 11210 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 13541 2907 13599 2913
rect 13541 2873 13553 2907
rect 13587 2904 13599 2907
rect 13906 2904 13912 2916
rect 13587 2876 13912 2904
rect 13587 2873 13599 2876
rect 13541 2867 13599 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 17034 2904 17040 2916
rect 16592 2876 17040 2904
rect 12710 2836 12716 2848
rect 9232 2808 12716 2836
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 12802 2796 12808 2848
rect 12860 2836 12866 2848
rect 14734 2836 14740 2848
rect 12860 2808 12905 2836
rect 14695 2808 14740 2836
rect 12860 2796 12866 2808
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 15105 2839 15163 2845
rect 15105 2805 15117 2839
rect 15151 2836 15163 2839
rect 15194 2836 15200 2848
rect 15151 2808 15200 2836
rect 15151 2805 15163 2808
rect 15105 2799 15163 2805
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2836 15531 2839
rect 15654 2836 15660 2848
rect 15519 2808 15660 2836
rect 15519 2805 15531 2808
rect 15473 2799 15531 2805
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 15841 2839 15899 2845
rect 15841 2805 15853 2839
rect 15887 2836 15899 2839
rect 16114 2836 16120 2848
rect 15887 2808 16120 2836
rect 15887 2805 15899 2808
rect 15841 2799 15899 2805
rect 16114 2796 16120 2808
rect 16172 2796 16178 2848
rect 16592 2845 16620 2876
rect 17034 2864 17040 2876
rect 17092 2864 17098 2916
rect 19886 2904 19892 2916
rect 19260 2876 19892 2904
rect 16577 2839 16635 2845
rect 16577 2805 16589 2839
rect 16623 2805 16635 2839
rect 16577 2799 16635 2805
rect 16945 2839 17003 2845
rect 16945 2805 16957 2839
rect 16991 2836 17003 2839
rect 17494 2836 17500 2848
rect 16991 2808 17500 2836
rect 16991 2805 17003 2808
rect 16945 2799 17003 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 17773 2839 17831 2845
rect 17773 2805 17785 2839
rect 17819 2836 17831 2839
rect 18138 2836 18144 2848
rect 17819 2808 18144 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 19260 2845 19288 2876
rect 19886 2864 19892 2876
rect 19944 2864 19950 2916
rect 19245 2839 19303 2845
rect 19245 2805 19257 2839
rect 19291 2805 19303 2839
rect 19245 2799 19303 2805
rect 20533 2839 20591 2845
rect 20533 2805 20545 2839
rect 20579 2836 20591 2839
rect 21266 2836 21272 2848
rect 20579 2808 21272 2836
rect 20579 2805 20591 2808
rect 20533 2799 20591 2805
rect 21266 2796 21272 2808
rect 21324 2796 21330 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1394 2632 1400 2644
rect 1355 2604 1400 2632
rect 1394 2592 1400 2604
rect 1452 2592 1458 2644
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 1946 2632 1952 2644
rect 1903 2604 1952 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2225 2635 2283 2641
rect 2225 2601 2237 2635
rect 2271 2601 2283 2635
rect 2590 2632 2596 2644
rect 2551 2604 2596 2632
rect 2225 2595 2283 2601
rect 1765 2567 1823 2573
rect 1765 2533 1777 2567
rect 1811 2564 1823 2567
rect 2240 2564 2268 2595
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 3694 2632 3700 2644
rect 3655 2604 3700 2632
rect 3694 2592 3700 2604
rect 3752 2592 3758 2644
rect 4154 2592 4160 2644
rect 4212 2632 4218 2644
rect 4709 2635 4767 2641
rect 4709 2632 4721 2635
rect 4212 2604 4721 2632
rect 4212 2592 4218 2604
rect 4709 2601 4721 2604
rect 4755 2632 4767 2635
rect 5074 2632 5080 2644
rect 4755 2604 5080 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5534 2632 5540 2644
rect 5495 2604 5540 2632
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 6086 2592 6092 2644
rect 6144 2632 6150 2644
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 6144 2604 6377 2632
rect 6144 2592 6150 2604
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8846 2632 8852 2644
rect 8067 2604 8852 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 10318 2632 10324 2644
rect 10279 2604 10324 2632
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 10594 2632 10600 2644
rect 10468 2604 10600 2632
rect 10468 2592 10474 2604
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 10962 2632 10968 2644
rect 10923 2604 10968 2632
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11471 2604 11897 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 11885 2601 11897 2604
rect 11931 2632 11943 2635
rect 11974 2632 11980 2644
rect 11931 2604 11980 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 14090 2592 14096 2644
rect 14148 2632 14154 2644
rect 14369 2635 14427 2641
rect 14369 2632 14381 2635
rect 14148 2604 14381 2632
rect 14148 2592 14154 2604
rect 14369 2601 14381 2604
rect 14415 2601 14427 2635
rect 14369 2595 14427 2601
rect 15197 2635 15255 2641
rect 15197 2601 15209 2635
rect 15243 2632 15255 2635
rect 15378 2632 15384 2644
rect 15243 2604 15384 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 15896 2604 15945 2632
rect 15896 2592 15902 2604
rect 15933 2601 15945 2604
rect 15979 2601 15991 2635
rect 15933 2595 15991 2601
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 16117 2635 16175 2641
rect 16117 2632 16129 2635
rect 16080 2604 16129 2632
rect 16080 2592 16086 2604
rect 16117 2601 16129 2604
rect 16163 2601 16175 2635
rect 16117 2595 16175 2601
rect 16669 2635 16727 2641
rect 16669 2601 16681 2635
rect 16715 2632 16727 2635
rect 16758 2632 16764 2644
rect 16715 2604 16764 2632
rect 16715 2601 16727 2604
rect 16669 2595 16727 2601
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 17218 2632 17224 2644
rect 17175 2604 17224 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 17310 2592 17316 2644
rect 17368 2632 17374 2644
rect 17405 2635 17463 2641
rect 17405 2632 17417 2635
rect 17368 2604 17417 2632
rect 17368 2592 17374 2604
rect 17405 2601 17417 2604
rect 17451 2601 17463 2635
rect 17405 2595 17463 2601
rect 17957 2635 18015 2641
rect 17957 2601 17969 2635
rect 18003 2632 18015 2635
rect 18046 2632 18052 2644
rect 18003 2604 18052 2632
rect 18003 2601 18015 2604
rect 17957 2595 18015 2601
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 18969 2635 19027 2641
rect 18969 2601 18981 2635
rect 19015 2632 19027 2635
rect 19058 2632 19064 2644
rect 19015 2604 19064 2632
rect 19015 2601 19027 2604
rect 18969 2595 19027 2601
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 1811 2536 2268 2564
rect 1811 2533 1823 2536
rect 1765 2527 1823 2533
rect 2682 2524 2688 2576
rect 2740 2524 2746 2576
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 7929 2567 7987 2573
rect 7929 2564 7941 2567
rect 7156 2536 7941 2564
rect 7156 2524 7162 2536
rect 7929 2533 7941 2536
rect 7975 2564 7987 2567
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 7975 2536 8493 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 8481 2533 8493 2536
rect 8527 2564 8539 2567
rect 9398 2564 9404 2576
rect 8527 2536 9404 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 9398 2524 9404 2536
rect 9456 2524 9462 2576
rect 10226 2564 10232 2576
rect 9784 2536 10232 2564
rect 2700 2496 2728 2524
rect 2700 2468 2820 2496
rect 2038 2428 2044 2440
rect 1999 2400 2044 2428
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 2792 2437 2820 2468
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4985 2499 5043 2505
rect 4985 2496 4997 2499
rect 4120 2468 4997 2496
rect 4120 2456 4126 2468
rect 4985 2465 4997 2468
rect 5031 2496 5043 2499
rect 5718 2496 5724 2508
rect 5031 2468 5724 2496
rect 5031 2465 5043 2468
rect 4985 2459 5043 2465
rect 5718 2456 5724 2468
rect 5776 2496 5782 2508
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5776 2468 5917 2496
rect 5776 2456 5782 2468
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 6638 2456 6644 2508
rect 6696 2496 6702 2508
rect 7653 2499 7711 2505
rect 7653 2496 7665 2499
rect 6696 2468 7665 2496
rect 6696 2456 6702 2468
rect 7653 2465 7665 2468
rect 7699 2496 7711 2499
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7699 2468 8401 2496
rect 7699 2465 7711 2468
rect 7653 2459 7711 2465
rect 8389 2465 8401 2468
rect 8435 2496 8447 2499
rect 9784 2496 9812 2536
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10796 2564 10824 2592
rect 11333 2567 11391 2573
rect 11333 2564 11345 2567
rect 10796 2536 11345 2564
rect 11333 2533 11345 2536
rect 11379 2533 11391 2567
rect 11333 2527 11391 2533
rect 12710 2524 12716 2576
rect 12768 2564 12774 2576
rect 12768 2536 13584 2564
rect 12768 2524 12774 2536
rect 8435 2468 9812 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10413 2499 10471 2505
rect 10413 2496 10425 2499
rect 10008 2468 10425 2496
rect 10008 2456 10014 2468
rect 10413 2465 10425 2468
rect 10459 2465 10471 2499
rect 10413 2459 10471 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 13556 2505 13584 2536
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12492 2468 12633 2496
rect 12492 2456 12498 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 13173 2499 13231 2505
rect 13173 2496 13185 2499
rect 12943 2468 13185 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 13173 2465 13185 2468
rect 13219 2465 13231 2499
rect 13173 2459 13231 2465
rect 13541 2499 13599 2505
rect 13541 2465 13553 2499
rect 13587 2465 13599 2499
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 13541 2459 13599 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 15565 2499 15623 2505
rect 15565 2465 15577 2499
rect 15611 2496 15623 2499
rect 15856 2496 15884 2592
rect 15611 2468 15884 2496
rect 15611 2465 15623 2468
rect 15565 2459 15623 2465
rect 2685 2431 2743 2437
rect 2685 2397 2697 2431
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2397 2835 2431
rect 5997 2431 6055 2437
rect 5997 2428 6009 2431
rect 2777 2391 2835 2397
rect 5184 2400 6009 2428
rect 2700 2360 2728 2391
rect 2866 2360 2872 2372
rect 2700 2332 2872 2360
rect 2866 2320 2872 2332
rect 2924 2360 2930 2372
rect 3237 2363 3295 2369
rect 3237 2360 3249 2363
rect 2924 2332 3249 2360
rect 2924 2320 2930 2332
rect 3237 2329 3249 2332
rect 3283 2329 3295 2363
rect 3237 2323 3295 2329
rect 5184 2304 5212 2400
rect 5997 2397 6009 2400
rect 6043 2397 6055 2431
rect 6178 2428 6184 2440
rect 6139 2400 6184 2428
rect 5997 2391 6055 2397
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 7800 2400 8585 2428
rect 7800 2388 7806 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 10594 2428 10600 2440
rect 10555 2400 10600 2428
rect 8573 2391 8631 2397
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 5350 2292 5356 2304
rect 5311 2264 5356 2292
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 8588 2292 8616 2391
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11256 2400 11529 2428
rect 9953 2363 10011 2369
rect 9953 2329 9965 2363
rect 9999 2360 10011 2363
rect 11146 2360 11152 2372
rect 9999 2332 11152 2360
rect 9999 2329 10011 2332
rect 9953 2323 10011 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 11256 2292 11284 2400
rect 11517 2397 11529 2400
rect 11563 2428 11575 2431
rect 11698 2428 11704 2440
rect 11563 2400 11704 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 8588 2264 11284 2292
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 13320 2264 13369 2292
rect 13320 2252 13326 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13722 2292 13728 2304
rect 13683 2264 13728 2292
rect 13357 2255 13415 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14093 2295 14151 2301
rect 14093 2261 14105 2295
rect 14139 2292 14151 2295
rect 14274 2292 14280 2304
rect 14139 2264 14280 2292
rect 14139 2261 14151 2264
rect 14093 2255 14151 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 6638 2088 6644 2100
rect 2096 2060 6644 2088
rect 2096 2048 2102 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 15746 2048 15752 2100
rect 15804 2088 15810 2100
rect 21726 2088 21732 2100
rect 15804 2060 21732 2088
rect 15804 2048 15810 2060
rect 21726 2048 21732 2060
rect 21784 2048 21790 2100
rect 658 1980 664 2032
rect 716 2020 722 2032
rect 6546 2020 6552 2032
rect 716 1992 6552 2020
rect 716 1980 722 1992
rect 6546 1980 6552 1992
rect 6604 1980 6610 2032
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 2780 20544 2832 20596
rect 2872 20476 2924 20528
rect 7104 20544 7156 20596
rect 7748 20544 7800 20596
rect 10784 20544 10836 20596
rect 6276 20451 6328 20460
rect 6276 20417 6285 20451
rect 6285 20417 6319 20451
rect 6319 20417 6328 20451
rect 6276 20408 6328 20417
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 2136 20383 2188 20392
rect 2136 20349 2145 20383
rect 2145 20349 2179 20383
rect 2179 20349 2188 20383
rect 2136 20340 2188 20349
rect 4528 20340 4580 20392
rect 8944 20340 8996 20392
rect 5540 20204 5592 20256
rect 6828 20272 6880 20324
rect 13268 20272 13320 20324
rect 21824 20272 21876 20324
rect 6552 20204 6604 20256
rect 7012 20204 7064 20256
rect 9588 20247 9640 20256
rect 9588 20213 9597 20247
rect 9597 20213 9631 20247
rect 9631 20213 9640 20247
rect 9588 20204 9640 20213
rect 13728 20204 13780 20256
rect 19524 20204 19576 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 4528 20043 4580 20052
rect 4528 20009 4537 20043
rect 4537 20009 4571 20043
rect 4571 20009 4580 20043
rect 4528 20000 4580 20009
rect 6828 20043 6880 20052
rect 6828 20009 6837 20043
rect 6837 20009 6871 20043
rect 6871 20009 6880 20043
rect 6828 20000 6880 20009
rect 7748 20043 7800 20052
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 8300 20000 8352 20052
rect 9588 20000 9640 20052
rect 12624 20000 12676 20052
rect 13084 20000 13136 20052
rect 13268 20043 13320 20052
rect 13268 20009 13277 20043
rect 13277 20009 13311 20043
rect 13311 20009 13320 20043
rect 13268 20000 13320 20009
rect 13728 20043 13780 20052
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 8668 19932 8720 19984
rect 11980 19932 12032 19984
rect 17224 20000 17276 20052
rect 2228 19907 2280 19916
rect 2228 19873 2237 19907
rect 2237 19873 2271 19907
rect 2271 19873 2280 19907
rect 2228 19864 2280 19873
rect 4160 19864 4212 19916
rect 6276 19864 6328 19916
rect 7012 19864 7064 19916
rect 9312 19864 9364 19916
rect 11060 19864 11112 19916
rect 12164 19864 12216 19916
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 21364 19932 21416 19984
rect 2780 19796 2832 19848
rect 4804 19796 4856 19848
rect 4896 19796 4948 19848
rect 7380 19796 7432 19848
rect 8116 19839 8168 19848
rect 2872 19728 2924 19780
rect 6184 19728 6236 19780
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 7288 19660 7340 19712
rect 8116 19805 8125 19839
rect 8125 19805 8159 19839
rect 8159 19805 8168 19839
rect 8116 19796 8168 19805
rect 9680 19703 9732 19712
rect 9680 19669 9689 19703
rect 9689 19669 9723 19703
rect 9723 19669 9732 19703
rect 9680 19660 9732 19669
rect 10324 19660 10376 19712
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 12440 19660 12492 19669
rect 12900 19660 12952 19712
rect 14556 19660 14608 19712
rect 16028 19660 16080 19712
rect 16580 19864 16632 19916
rect 20904 19728 20956 19780
rect 18788 19660 18840 19712
rect 19156 19660 19208 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1676 19499 1728 19508
rect 1676 19465 1685 19499
rect 1685 19465 1719 19499
rect 1719 19465 1728 19499
rect 1676 19456 1728 19465
rect 2228 19456 2280 19508
rect 1768 19320 1820 19372
rect 2872 19363 2924 19372
rect 2872 19329 2881 19363
rect 2881 19329 2915 19363
rect 2915 19329 2924 19363
rect 2872 19320 2924 19329
rect 4896 19456 4948 19508
rect 6276 19456 6328 19508
rect 4712 19388 4764 19440
rect 2504 19252 2556 19304
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 2780 19252 2832 19261
rect 4712 19295 4764 19304
rect 2596 19184 2648 19236
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 6920 19320 6972 19372
rect 8116 19456 8168 19508
rect 8668 19363 8720 19372
rect 8668 19329 8677 19363
rect 8677 19329 8711 19363
rect 8711 19329 8720 19363
rect 8668 19320 8720 19329
rect 6184 19295 6236 19304
rect 6184 19261 6193 19295
rect 6193 19261 6227 19295
rect 6227 19261 6236 19295
rect 6184 19252 6236 19261
rect 7288 19295 7340 19304
rect 4804 19184 4856 19236
rect 5080 19184 5132 19236
rect 7288 19261 7322 19295
rect 7322 19261 7340 19295
rect 7288 19252 7340 19261
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 9036 19184 9088 19236
rect 10324 19252 10376 19304
rect 11060 19456 11112 19508
rect 12164 19499 12216 19508
rect 12164 19465 12173 19499
rect 12173 19465 12207 19499
rect 12207 19465 12216 19499
rect 12164 19456 12216 19465
rect 15384 19456 15436 19508
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12716 19252 12768 19304
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 11428 19184 11480 19236
rect 13452 19184 13504 19236
rect 14280 19252 14332 19304
rect 14740 19252 14792 19304
rect 15384 19252 15436 19304
rect 15660 19295 15712 19304
rect 15660 19261 15669 19295
rect 15669 19261 15703 19295
rect 15703 19261 15712 19295
rect 15660 19252 15712 19261
rect 15936 19252 15988 19304
rect 16856 19252 16908 19304
rect 17500 19295 17552 19304
rect 17500 19261 17509 19295
rect 17509 19261 17543 19295
rect 17543 19261 17552 19295
rect 17500 19252 17552 19261
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 18788 19295 18840 19304
rect 18788 19261 18797 19295
rect 18797 19261 18831 19295
rect 18831 19261 18840 19295
rect 18788 19252 18840 19261
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19524 19295 19576 19304
rect 19524 19261 19533 19295
rect 19533 19261 19567 19295
rect 19567 19261 19576 19295
rect 19524 19252 19576 19261
rect 7380 19116 7432 19168
rect 9312 19116 9364 19168
rect 13544 19116 13596 19168
rect 14372 19184 14424 19236
rect 14924 19184 14976 19236
rect 15752 19116 15804 19168
rect 16304 19184 16356 19236
rect 17224 19227 17276 19236
rect 17224 19193 17233 19227
rect 17233 19193 17267 19227
rect 17267 19193 17276 19227
rect 17224 19184 17276 19193
rect 16764 19116 16816 19168
rect 17684 19159 17736 19168
rect 17684 19125 17693 19159
rect 17693 19125 17727 19159
rect 17727 19125 17736 19159
rect 17684 19116 17736 19125
rect 18144 19116 18196 19168
rect 18604 19159 18656 19168
rect 18604 19125 18613 19159
rect 18613 19125 18647 19159
rect 18647 19125 18656 19159
rect 18604 19116 18656 19125
rect 19064 19116 19116 19168
rect 19984 19184 20036 19236
rect 20444 19116 20496 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 1124 18844 1176 18896
rect 4620 18912 4672 18964
rect 4804 18912 4856 18964
rect 8484 18912 8536 18964
rect 9680 18912 9732 18964
rect 12256 18955 12308 18964
rect 12256 18921 12265 18955
rect 12265 18921 12299 18955
rect 12299 18921 12308 18955
rect 12256 18912 12308 18921
rect 12808 18912 12860 18964
rect 2136 18844 2188 18896
rect 5724 18844 5776 18896
rect 6368 18844 6420 18896
rect 7380 18844 7432 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 4712 18776 4764 18828
rect 6920 18819 6972 18828
rect 6920 18785 6929 18819
rect 6929 18785 6963 18819
rect 6963 18785 6972 18819
rect 6920 18776 6972 18785
rect 8760 18776 8812 18828
rect 10876 18776 10928 18828
rect 11704 18776 11756 18828
rect 12440 18844 12492 18896
rect 15936 18912 15988 18964
rect 14740 18844 14792 18896
rect 4252 18708 4304 18760
rect 9312 18751 9364 18760
rect 664 18572 716 18624
rect 2688 18572 2740 18624
rect 3976 18572 4028 18624
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 10692 18708 10744 18760
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 12348 18751 12400 18760
rect 11428 18708 11480 18717
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 13912 18776 13964 18828
rect 15200 18776 15252 18828
rect 18420 18844 18472 18896
rect 6000 18640 6052 18692
rect 4896 18572 4948 18624
rect 12440 18640 12492 18692
rect 16856 18776 16908 18828
rect 19524 18844 19576 18896
rect 17500 18708 17552 18760
rect 22284 18708 22336 18760
rect 8944 18572 8996 18624
rect 11244 18572 11296 18624
rect 11796 18615 11848 18624
rect 11796 18581 11805 18615
rect 11805 18581 11839 18615
rect 11839 18581 11848 18615
rect 11796 18572 11848 18581
rect 12808 18572 12860 18624
rect 14096 18572 14148 18624
rect 15384 18615 15436 18624
rect 15384 18581 15393 18615
rect 15393 18581 15427 18615
rect 15427 18581 15436 18615
rect 15384 18572 15436 18581
rect 15660 18572 15712 18624
rect 16304 18572 16356 18624
rect 18052 18572 18104 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1584 18368 1636 18420
rect 2504 18368 2556 18420
rect 1952 18343 2004 18352
rect 1952 18309 1961 18343
rect 1961 18309 1995 18343
rect 1995 18309 2004 18343
rect 1952 18300 2004 18309
rect 3976 18411 4028 18420
rect 3976 18377 3985 18411
rect 3985 18377 4019 18411
rect 4019 18377 4028 18411
rect 4252 18411 4304 18420
rect 3976 18368 4028 18377
rect 4252 18377 4261 18411
rect 4261 18377 4295 18411
rect 4295 18377 4304 18411
rect 4252 18368 4304 18377
rect 4804 18368 4856 18420
rect 10140 18368 10192 18420
rect 10876 18411 10928 18420
rect 10876 18377 10885 18411
rect 10885 18377 10919 18411
rect 10919 18377 10928 18411
rect 10876 18368 10928 18377
rect 7748 18300 7800 18352
rect 2596 18275 2648 18284
rect 2596 18241 2605 18275
rect 2605 18241 2639 18275
rect 2639 18241 2648 18275
rect 2596 18232 2648 18241
rect 4896 18275 4948 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 4896 18241 4905 18275
rect 4905 18241 4939 18275
rect 4939 18241 4948 18275
rect 4896 18232 4948 18241
rect 5540 18275 5592 18284
rect 5540 18241 5549 18275
rect 5549 18241 5583 18275
rect 5583 18241 5592 18275
rect 5540 18232 5592 18241
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 9956 18232 10008 18284
rect 12164 18300 12216 18352
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 12348 18368 12400 18420
rect 14096 18368 14148 18420
rect 17776 18368 17828 18420
rect 12440 18300 12492 18352
rect 14464 18300 14516 18352
rect 19156 18300 19208 18352
rect 5080 18164 5132 18216
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 11244 18207 11296 18216
rect 11244 18173 11253 18207
rect 11253 18173 11287 18207
rect 11287 18173 11296 18207
rect 11244 18164 11296 18173
rect 11796 18164 11848 18216
rect 12440 18207 12492 18216
rect 12440 18173 12456 18207
rect 12456 18173 12490 18207
rect 12490 18173 12492 18207
rect 12440 18164 12492 18173
rect 2780 18096 2832 18148
rect 5264 18096 5316 18148
rect 6276 18096 6328 18148
rect 10784 18096 10836 18148
rect 12532 18096 12584 18148
rect 1400 18071 1452 18080
rect 1400 18037 1409 18071
rect 1409 18037 1443 18071
rect 1443 18037 1452 18071
rect 1400 18028 1452 18037
rect 4436 18028 4488 18080
rect 5356 18028 5408 18080
rect 8852 18071 8904 18080
rect 8852 18037 8861 18071
rect 8861 18037 8895 18071
rect 8895 18037 8904 18071
rect 8852 18028 8904 18037
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 9680 18028 9732 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 4344 17824 4396 17876
rect 5264 17824 5316 17876
rect 5356 17824 5408 17876
rect 9220 17824 9272 17876
rect 1768 17756 1820 17808
rect 2780 17799 2832 17808
rect 2780 17765 2789 17799
rect 2789 17765 2823 17799
rect 2823 17765 2832 17799
rect 2780 17756 2832 17765
rect 1860 17688 1912 17740
rect 2504 17731 2556 17740
rect 2504 17697 2513 17731
rect 2513 17697 2547 17731
rect 2547 17697 2556 17731
rect 2504 17688 2556 17697
rect 8852 17756 8904 17808
rect 2964 17552 3016 17604
rect 3056 17552 3108 17604
rect 6460 17688 6512 17740
rect 9128 17731 9180 17740
rect 9128 17697 9137 17731
rect 9137 17697 9171 17731
rect 9171 17697 9180 17731
rect 9128 17688 9180 17697
rect 4804 17620 4856 17672
rect 6552 17620 6604 17672
rect 7380 17620 7432 17672
rect 10692 17756 10744 17808
rect 14004 17824 14056 17876
rect 12072 17756 12124 17808
rect 9772 17688 9824 17740
rect 9956 17731 10008 17740
rect 9956 17697 9990 17731
rect 9990 17697 10008 17731
rect 9956 17688 10008 17697
rect 11060 17688 11112 17740
rect 3148 17484 3200 17536
rect 7104 17484 7156 17536
rect 9588 17484 9640 17536
rect 11244 17688 11296 17740
rect 12440 17688 12492 17740
rect 13360 17688 13412 17740
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1676 17280 1728 17332
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 4068 17280 4120 17332
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 4896 17280 4948 17332
rect 6460 17187 6512 17196
rect 3976 17076 4028 17128
rect 4068 17076 4120 17128
rect 4804 17076 4856 17128
rect 6460 17153 6469 17187
rect 6469 17153 6503 17187
rect 6503 17153 6512 17187
rect 6460 17144 6512 17153
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 8116 17144 8168 17196
rect 6736 17008 6788 17060
rect 6920 17076 6972 17128
rect 7380 17076 7432 17128
rect 8208 17076 8260 17128
rect 7196 17008 7248 17060
rect 8116 17008 8168 17060
rect 2136 16940 2188 16992
rect 2964 16983 3016 16992
rect 2964 16949 2973 16983
rect 2973 16949 3007 16983
rect 3007 16949 3016 16983
rect 2964 16940 3016 16949
rect 3424 16940 3476 16992
rect 6644 16940 6696 16992
rect 7380 16940 7432 16992
rect 9772 17280 9824 17332
rect 9956 17280 10008 17332
rect 12072 17187 12124 17196
rect 9588 17076 9640 17128
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 10324 17076 10376 17128
rect 12900 17076 12952 17128
rect 14188 17076 14240 17128
rect 17960 17008 18012 17060
rect 11336 16940 11388 16992
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 11888 16940 11940 16992
rect 15476 16940 15528 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2964 16736 3016 16788
rect 1860 16668 1912 16720
rect 3240 16668 3292 16720
rect 4896 16736 4948 16788
rect 6920 16736 6972 16788
rect 7104 16779 7156 16788
rect 7104 16745 7113 16779
rect 7113 16745 7147 16779
rect 7147 16745 7156 16779
rect 7104 16736 7156 16745
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 10600 16736 10652 16788
rect 11336 16779 11388 16788
rect 6828 16668 6880 16720
rect 7288 16668 7340 16720
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 11520 16736 11572 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 2136 16643 2188 16652
rect 2136 16609 2145 16643
rect 2145 16609 2179 16643
rect 2179 16609 2188 16643
rect 2136 16600 2188 16609
rect 4252 16600 4304 16652
rect 5264 16600 5316 16652
rect 4804 16532 4856 16584
rect 7380 16575 7432 16584
rect 4896 16464 4948 16516
rect 5080 16464 5132 16516
rect 3516 16396 3568 16448
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 6736 16507 6788 16516
rect 6736 16473 6745 16507
rect 6745 16473 6779 16507
rect 6779 16473 6788 16507
rect 6736 16464 6788 16473
rect 7196 16396 7248 16448
rect 10048 16600 10100 16652
rect 10232 16600 10284 16652
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 8208 16532 8260 16541
rect 10324 16575 10376 16584
rect 10324 16541 10333 16575
rect 10333 16541 10367 16575
rect 10367 16541 10376 16575
rect 10324 16532 10376 16541
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 10692 16532 10744 16584
rect 11152 16464 11204 16516
rect 12072 16532 12124 16584
rect 12532 16532 12584 16584
rect 10508 16396 10560 16448
rect 10876 16396 10928 16448
rect 11244 16396 11296 16448
rect 12532 16396 12584 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 1400 16056 1452 16108
rect 4068 16192 4120 16244
rect 5264 16192 5316 16244
rect 6828 16192 6880 16244
rect 7196 16124 7248 16176
rect 8852 16192 8904 16244
rect 9864 16192 9916 16244
rect 11796 16192 11848 16244
rect 11980 16192 12032 16244
rect 3516 15988 3568 16040
rect 5724 15988 5776 16040
rect 2872 15920 2924 15972
rect 4620 15920 4672 15972
rect 8668 15920 8720 15972
rect 2688 15852 2740 15904
rect 8208 15852 8260 15904
rect 11428 16056 11480 16108
rect 12624 16056 12676 16108
rect 11244 15988 11296 16040
rect 12532 15988 12584 16040
rect 8852 15852 8904 15904
rect 14096 15920 14148 15972
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 11152 15852 11204 15904
rect 14648 15852 14700 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 4252 15648 4304 15700
rect 4344 15648 4396 15700
rect 8668 15691 8720 15700
rect 8668 15657 8677 15691
rect 8677 15657 8711 15691
rect 8711 15657 8720 15691
rect 8668 15648 8720 15657
rect 9036 15648 9088 15700
rect 10600 15648 10652 15700
rect 10968 15648 11020 15700
rect 11060 15648 11112 15700
rect 12624 15691 12676 15700
rect 5540 15580 5592 15632
rect 2320 15512 2372 15564
rect 3424 15512 3476 15564
rect 4160 15512 4212 15564
rect 7288 15580 7340 15632
rect 7380 15580 7432 15632
rect 7748 15580 7800 15632
rect 8208 15580 8260 15632
rect 9956 15580 10008 15632
rect 10140 15580 10192 15632
rect 10692 15580 10744 15632
rect 6920 15512 6972 15564
rect 7196 15512 7248 15564
rect 1768 15444 1820 15496
rect 4620 15487 4672 15496
rect 4620 15453 4629 15487
rect 4629 15453 4663 15487
rect 4663 15453 4672 15487
rect 4620 15444 4672 15453
rect 7288 15487 7340 15496
rect 7288 15453 7297 15487
rect 7297 15453 7331 15487
rect 7331 15453 7340 15487
rect 7288 15444 7340 15453
rect 8668 15444 8720 15496
rect 9036 15444 9088 15496
rect 7196 15351 7248 15360
rect 7196 15317 7205 15351
rect 7205 15317 7239 15351
rect 7239 15317 7248 15351
rect 7196 15308 7248 15317
rect 10416 15444 10468 15496
rect 11428 15580 11480 15632
rect 11704 15580 11756 15632
rect 12624 15657 12633 15691
rect 12633 15657 12667 15691
rect 12667 15657 12676 15691
rect 12624 15648 12676 15657
rect 13268 15648 13320 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 12532 15512 12584 15564
rect 13268 15512 13320 15564
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 11060 15444 11112 15496
rect 14188 15419 14240 15428
rect 10968 15308 11020 15360
rect 14188 15385 14197 15419
rect 14197 15385 14231 15419
rect 14231 15385 14240 15419
rect 14188 15376 14240 15385
rect 14004 15308 14056 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 5540 15104 5592 15156
rect 6644 15104 6696 15156
rect 8944 15147 8996 15156
rect 5724 15036 5776 15088
rect 2872 15011 2924 15020
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 3884 14968 3936 15020
rect 7196 14968 7248 15020
rect 8944 15113 8953 15147
rect 8953 15113 8987 15147
rect 8987 15113 8996 15147
rect 8944 15104 8996 15113
rect 9220 15036 9272 15088
rect 9864 15104 9916 15156
rect 11060 15104 11112 15156
rect 11244 15104 11296 15156
rect 6920 14900 6972 14952
rect 9128 14968 9180 15020
rect 9036 14900 9088 14952
rect 9496 15011 9548 15020
rect 9496 14977 9505 15011
rect 9505 14977 9539 15011
rect 9539 14977 9548 15011
rect 9496 14968 9548 14977
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 10876 14968 10928 15020
rect 13176 15104 13228 15156
rect 14556 15104 14608 15156
rect 14188 15079 14240 15088
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 10416 14900 10468 14952
rect 3792 14832 3844 14884
rect 3332 14764 3384 14816
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 6368 14807 6420 14816
rect 3608 14764 3660 14773
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 9220 14832 9272 14884
rect 10692 14832 10744 14884
rect 10968 14832 11020 14884
rect 11888 14832 11940 14884
rect 7012 14764 7064 14816
rect 8484 14764 8536 14816
rect 10784 14764 10836 14816
rect 11060 14764 11112 14816
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11244 14764 11296 14773
rect 11336 14764 11388 14816
rect 14188 15045 14197 15079
rect 14197 15045 14231 15079
rect 14231 15045 14240 15079
rect 14188 15036 14240 15045
rect 12532 14968 12584 15020
rect 13268 14968 13320 15020
rect 13544 14900 13596 14952
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 14096 14900 14148 14952
rect 14648 14943 14700 14952
rect 14648 14909 14682 14943
rect 14682 14909 14700 14943
rect 14648 14900 14700 14909
rect 13452 14832 13504 14884
rect 13728 14875 13780 14884
rect 13728 14841 13737 14875
rect 13737 14841 13771 14875
rect 13771 14841 13780 14875
rect 13728 14832 13780 14841
rect 13084 14764 13136 14816
rect 13176 14764 13228 14816
rect 18788 14832 18840 14884
rect 15292 14764 15344 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2780 14560 2832 14612
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 6368 14560 6420 14612
rect 9036 14603 9088 14612
rect 2136 14467 2188 14476
rect 2136 14433 2145 14467
rect 2145 14433 2179 14467
rect 2179 14433 2188 14467
rect 2136 14424 2188 14433
rect 3884 14424 3936 14476
rect 7656 14424 7708 14476
rect 2320 14356 2372 14408
rect 5540 14399 5592 14408
rect 2044 14288 2096 14340
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 6920 14331 6972 14340
rect 6920 14297 6929 14331
rect 6929 14297 6963 14331
rect 6963 14297 6972 14331
rect 9036 14569 9045 14603
rect 9045 14569 9079 14603
rect 9079 14569 9088 14603
rect 9036 14560 9088 14569
rect 9680 14560 9732 14612
rect 10876 14560 10928 14612
rect 10968 14560 11020 14612
rect 13084 14603 13136 14612
rect 9220 14467 9272 14476
rect 9220 14433 9229 14467
rect 9229 14433 9263 14467
rect 9263 14433 9272 14467
rect 9220 14424 9272 14433
rect 9404 14424 9456 14476
rect 6920 14288 6972 14297
rect 9864 14424 9916 14476
rect 10324 14424 10376 14476
rect 10784 14492 10836 14544
rect 11336 14535 11388 14544
rect 11336 14501 11345 14535
rect 11345 14501 11379 14535
rect 11379 14501 11388 14535
rect 11336 14492 11388 14501
rect 12808 14492 12860 14544
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 13176 14560 13228 14612
rect 13728 14560 13780 14612
rect 14188 14560 14240 14612
rect 15568 14560 15620 14612
rect 22744 14560 22796 14612
rect 13452 14535 13504 14544
rect 10600 14424 10652 14476
rect 10876 14467 10928 14476
rect 10876 14433 10885 14467
rect 10885 14433 10919 14467
rect 10919 14433 10928 14467
rect 10876 14424 10928 14433
rect 11704 14424 11756 14476
rect 12532 14424 12584 14476
rect 11980 14356 12032 14408
rect 13452 14501 13461 14535
rect 13461 14501 13495 14535
rect 13495 14501 13504 14535
rect 13452 14492 13504 14501
rect 14556 14535 14608 14544
rect 14556 14501 14565 14535
rect 14565 14501 14599 14535
rect 14599 14501 14608 14535
rect 14556 14492 14608 14501
rect 14372 14424 14424 14476
rect 11244 14288 11296 14340
rect 13176 14288 13228 14340
rect 4068 14220 4120 14272
rect 7012 14263 7064 14272
rect 7012 14229 7021 14263
rect 7021 14229 7055 14263
rect 7055 14229 7064 14263
rect 7012 14220 7064 14229
rect 10232 14263 10284 14272
rect 10232 14229 10241 14263
rect 10241 14229 10275 14263
rect 10275 14229 10284 14263
rect 10232 14220 10284 14229
rect 10784 14220 10836 14272
rect 11980 14220 12032 14272
rect 12624 14220 12676 14272
rect 13084 14220 13136 14272
rect 13728 14399 13780 14408
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15108 14220 15160 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 2780 14059 2832 14068
rect 2780 14025 2789 14059
rect 2789 14025 2823 14059
rect 2823 14025 2832 14059
rect 3332 14059 3384 14068
rect 2780 14016 2832 14025
rect 3332 14025 3341 14059
rect 3341 14025 3375 14059
rect 3375 14025 3384 14059
rect 3332 14016 3384 14025
rect 3608 14016 3660 14068
rect 9312 14059 9364 14068
rect 3884 13923 3936 13932
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2320 13855 2372 13864
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 2504 13812 2556 13864
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 5816 13880 5868 13932
rect 7196 13880 7248 13932
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 11152 14016 11204 14068
rect 12900 14016 12952 14068
rect 13176 14016 13228 14068
rect 13544 14059 13596 14068
rect 13544 14025 13553 14059
rect 13553 14025 13587 14059
rect 13587 14025 13596 14059
rect 13544 14016 13596 14025
rect 8944 13880 8996 13932
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 11060 13880 11112 13932
rect 4804 13812 4856 13864
rect 5632 13812 5684 13864
rect 5724 13855 5776 13864
rect 5724 13821 5733 13855
rect 5733 13821 5767 13855
rect 5767 13821 5776 13855
rect 5724 13812 5776 13821
rect 6092 13812 6144 13864
rect 7840 13812 7892 13864
rect 8024 13812 8076 13864
rect 9864 13855 9916 13864
rect 2964 13676 3016 13728
rect 3884 13676 3936 13728
rect 4068 13676 4120 13728
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 7104 13719 7156 13728
rect 7104 13685 7113 13719
rect 7113 13685 7147 13719
rect 7147 13685 7156 13719
rect 7104 13676 7156 13685
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 10232 13812 10284 13864
rect 9496 13744 9548 13796
rect 10692 13787 10744 13796
rect 10692 13753 10701 13787
rect 10701 13753 10735 13787
rect 10735 13753 10744 13787
rect 10692 13744 10744 13753
rect 10784 13744 10836 13796
rect 13268 13812 13320 13864
rect 13452 13880 13504 13932
rect 14464 14016 14516 14068
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 15752 13948 15804 14000
rect 15108 13923 15160 13932
rect 13544 13812 13596 13864
rect 13636 13812 13688 13864
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 14372 13812 14424 13864
rect 15568 13812 15620 13864
rect 12808 13744 12860 13796
rect 11520 13676 11572 13728
rect 12716 13719 12768 13728
rect 12716 13685 12725 13719
rect 12725 13685 12759 13719
rect 12759 13685 12768 13719
rect 12716 13676 12768 13685
rect 13084 13676 13136 13728
rect 13268 13676 13320 13728
rect 18052 13744 18104 13796
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 1768 13515 1820 13524
rect 1768 13481 1777 13515
rect 1777 13481 1811 13515
rect 1811 13481 1820 13515
rect 1768 13472 1820 13481
rect 5632 13472 5684 13524
rect 5540 13404 5592 13456
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 3240 13379 3292 13388
rect 3240 13345 3249 13379
rect 3249 13345 3283 13379
rect 3283 13345 3292 13379
rect 3240 13336 3292 13345
rect 4068 13336 4120 13388
rect 2412 13268 2464 13320
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 7104 13472 7156 13524
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 9404 13472 9456 13524
rect 9588 13472 9640 13524
rect 9864 13472 9916 13524
rect 12716 13472 12768 13524
rect 12900 13472 12952 13524
rect 13544 13472 13596 13524
rect 9772 13404 9824 13456
rect 14096 13404 14148 13456
rect 14372 13472 14424 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 9128 13336 9180 13388
rect 11612 13336 11664 13388
rect 12072 13336 12124 13388
rect 12716 13336 12768 13388
rect 12900 13336 12952 13388
rect 13360 13379 13412 13388
rect 13360 13345 13369 13379
rect 13369 13345 13403 13379
rect 13403 13345 13412 13379
rect 13360 13336 13412 13345
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 7840 13311 7892 13320
rect 5816 13200 5868 13252
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 8484 13268 8536 13320
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 9312 13268 9364 13320
rect 10968 13268 11020 13320
rect 11152 13268 11204 13320
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 12624 13268 12676 13320
rect 13636 13311 13688 13320
rect 6736 13200 6788 13252
rect 8392 13200 8444 13252
rect 2872 13132 2924 13184
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 9588 13132 9640 13184
rect 13360 13200 13412 13252
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 14188 13200 14240 13252
rect 12716 13132 12768 13184
rect 15752 13132 15804 13184
rect 18604 13132 18656 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 3332 12928 3384 12980
rect 2412 12792 2464 12844
rect 2044 12724 2096 12776
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 2228 12656 2280 12708
rect 3516 12656 3568 12708
rect 4988 12928 5040 12980
rect 3884 12860 3936 12912
rect 9772 12928 9824 12980
rect 13636 12928 13688 12980
rect 15660 12971 15712 12980
rect 15660 12937 15669 12971
rect 15669 12937 15703 12971
rect 15703 12937 15712 12971
rect 15660 12928 15712 12937
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 3976 12767 4028 12776
rect 3976 12733 3985 12767
rect 3985 12733 4019 12767
rect 4019 12733 4028 12767
rect 3976 12724 4028 12733
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7104 12767 7156 12776
rect 7104 12733 7138 12767
rect 7138 12733 7156 12767
rect 7932 12860 7984 12912
rect 9956 12860 10008 12912
rect 15568 12903 15620 12912
rect 7104 12724 7156 12733
rect 6092 12656 6144 12708
rect 2596 12588 2648 12640
rect 6828 12588 6880 12640
rect 8208 12724 8260 12776
rect 10784 12792 10836 12844
rect 15568 12869 15577 12903
rect 15577 12869 15611 12903
rect 15611 12869 15620 12903
rect 15568 12860 15620 12869
rect 15844 12860 15896 12912
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 13820 12792 13872 12844
rect 14004 12792 14056 12844
rect 15292 12792 15344 12844
rect 10692 12724 10744 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 11244 12724 11296 12776
rect 12532 12724 12584 12776
rect 12716 12767 12768 12776
rect 12716 12733 12750 12767
rect 12750 12733 12768 12767
rect 12716 12724 12768 12733
rect 13268 12724 13320 12776
rect 13728 12724 13780 12776
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 14740 12724 14792 12776
rect 15384 12724 15436 12776
rect 16580 12724 16632 12776
rect 8208 12631 8260 12640
rect 8208 12597 8217 12631
rect 8217 12597 8251 12631
rect 8251 12597 8260 12631
rect 8208 12588 8260 12597
rect 9864 12588 9916 12640
rect 10048 12588 10100 12640
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 11612 12656 11664 12708
rect 10232 12588 10284 12597
rect 11704 12588 11756 12640
rect 13728 12588 13780 12640
rect 16304 12588 16356 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 3516 12384 3568 12436
rect 3608 12384 3660 12436
rect 4252 12384 4304 12436
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 6828 12384 6880 12436
rect 7288 12384 7340 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 10232 12384 10284 12436
rect 10784 12384 10836 12436
rect 11428 12384 11480 12436
rect 12992 12384 13044 12436
rect 15200 12384 15252 12436
rect 15752 12427 15804 12436
rect 15752 12393 15761 12427
rect 15761 12393 15795 12427
rect 15795 12393 15804 12427
rect 15752 12384 15804 12393
rect 2044 12291 2096 12300
rect 2044 12257 2053 12291
rect 2053 12257 2087 12291
rect 2087 12257 2096 12291
rect 2044 12248 2096 12257
rect 3056 12248 3108 12300
rect 4252 12248 4304 12300
rect 5264 12180 5316 12232
rect 7196 12316 7248 12368
rect 9772 12316 9824 12368
rect 9956 12359 10008 12368
rect 9956 12325 9990 12359
rect 9990 12325 10008 12359
rect 9956 12316 10008 12325
rect 15568 12316 15620 12368
rect 6184 12248 6236 12300
rect 9496 12248 9548 12300
rect 11152 12291 11204 12300
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 11428 12291 11480 12300
rect 11428 12257 11462 12291
rect 11462 12257 11480 12291
rect 11428 12248 11480 12257
rect 12256 12248 12308 12300
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 13728 12291 13780 12300
rect 13728 12257 13737 12291
rect 13737 12257 13771 12291
rect 13771 12257 13780 12291
rect 13728 12248 13780 12257
rect 14280 12248 14332 12300
rect 8208 12180 8260 12232
rect 12716 12180 12768 12232
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 5080 12044 5132 12096
rect 7012 12087 7064 12096
rect 7012 12053 7021 12087
rect 7021 12053 7055 12087
rect 7055 12053 7064 12087
rect 7012 12044 7064 12053
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 8668 12044 8720 12096
rect 8852 12044 8904 12096
rect 15200 12112 15252 12164
rect 10600 12044 10652 12096
rect 11796 12044 11848 12096
rect 12072 12044 12124 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 16304 12044 16356 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2320 11840 2372 11892
rect 3240 11840 3292 11892
rect 6184 11840 6236 11892
rect 7380 11840 7432 11892
rect 9956 11840 10008 11892
rect 11704 11840 11756 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13084 11840 13136 11892
rect 3976 11772 4028 11824
rect 8392 11772 8444 11824
rect 9036 11772 9088 11824
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 4068 11704 4120 11756
rect 4252 11704 4304 11756
rect 5080 11704 5132 11756
rect 7012 11704 7064 11756
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 8852 11704 8904 11756
rect 9588 11704 9640 11756
rect 11152 11772 11204 11824
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 13728 11772 13780 11824
rect 11796 11704 11848 11756
rect 12532 11704 12584 11756
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 2320 11636 2372 11688
rect 3424 11636 3476 11688
rect 3884 11636 3936 11688
rect 6828 11636 6880 11688
rect 7104 11636 7156 11688
rect 12900 11636 12952 11688
rect 14096 11636 14148 11688
rect 15200 11679 15252 11688
rect 1492 11611 1544 11620
rect 1492 11577 1501 11611
rect 1501 11577 1535 11611
rect 1535 11577 1544 11611
rect 1492 11568 1544 11577
rect 2964 11568 3016 11620
rect 4896 11568 4948 11620
rect 5080 11568 5132 11620
rect 6736 11568 6788 11620
rect 7380 11568 7432 11620
rect 9680 11568 9732 11620
rect 10876 11568 10928 11620
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 4252 11500 4304 11552
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 5448 11543 5500 11552
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5448 11500 5500 11509
rect 7012 11500 7064 11552
rect 9496 11500 9548 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 14188 11568 14240 11620
rect 15200 11645 15234 11679
rect 15234 11645 15252 11679
rect 15200 11636 15252 11645
rect 15292 11568 15344 11620
rect 11704 11500 11756 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 14096 11543 14148 11552
rect 12900 11500 12952 11509
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 14372 11500 14424 11552
rect 15200 11500 15252 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1952 11296 2004 11348
rect 5356 11296 5408 11348
rect 6828 11296 6880 11348
rect 2964 11228 3016 11280
rect 3608 11228 3660 11280
rect 4068 11228 4120 11280
rect 7288 11228 7340 11280
rect 2320 11160 2372 11212
rect 6736 11203 6788 11212
rect 6736 11169 6770 11203
rect 6770 11169 6788 11203
rect 6736 11160 6788 11169
rect 8208 11203 8260 11212
rect 3056 11092 3108 11144
rect 3700 11092 3752 11144
rect 3976 10956 4028 11008
rect 4988 11024 5040 11076
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 6460 11135 6512 11144
rect 5264 11092 5316 11101
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 8208 11169 8242 11203
rect 8242 11169 8260 11203
rect 8208 11160 8260 11169
rect 8668 11296 8720 11348
rect 9220 11228 9272 11280
rect 12900 11296 12952 11348
rect 13912 11296 13964 11348
rect 14096 11296 14148 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 17224 11228 17276 11280
rect 11244 11160 11296 11212
rect 12440 11160 12492 11212
rect 6460 10956 6512 11008
rect 11888 11092 11940 11144
rect 11980 11092 12032 11144
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 13728 11135 13780 11144
rect 12256 11092 12308 11101
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 13912 11092 13964 11101
rect 8944 11024 8996 11076
rect 9220 11024 9272 11076
rect 8300 10956 8352 11008
rect 8576 10956 8628 11008
rect 10416 11024 10468 11076
rect 17500 11160 17552 11212
rect 14740 11135 14792 11144
rect 14740 11101 14749 11135
rect 14749 11101 14783 11135
rect 14783 11101 14792 11135
rect 14740 11092 14792 11101
rect 15568 11092 15620 11144
rect 14280 11067 14332 11076
rect 14280 11033 14289 11067
rect 14289 11033 14323 11067
rect 14323 11033 14332 11067
rect 14280 11024 14332 11033
rect 9496 10956 9548 11008
rect 12624 10956 12676 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 1584 10752 1636 10804
rect 5448 10752 5500 10804
rect 7012 10752 7064 10804
rect 7104 10684 7156 10736
rect 3884 10616 3936 10668
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5264 10616 5316 10668
rect 1860 10548 1912 10600
rect 2596 10548 2648 10600
rect 3608 10548 3660 10600
rect 6736 10616 6788 10668
rect 11704 10752 11756 10804
rect 13728 10752 13780 10804
rect 14740 10752 14792 10804
rect 9588 10684 9640 10736
rect 9404 10616 9456 10668
rect 10600 10616 10652 10668
rect 12256 10616 12308 10668
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 8300 10591 8352 10600
rect 8300 10557 8309 10591
rect 8309 10557 8343 10591
rect 8343 10557 8352 10591
rect 8300 10548 8352 10557
rect 4344 10480 4396 10532
rect 1492 10412 1544 10464
rect 2320 10412 2372 10464
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3884 10412 3936 10464
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 4620 10455 4672 10464
rect 4620 10421 4629 10455
rect 4629 10421 4663 10455
rect 4663 10421 4672 10455
rect 4620 10412 4672 10421
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 8208 10480 8260 10532
rect 10324 10548 10376 10600
rect 10784 10548 10836 10600
rect 11152 10548 11204 10600
rect 8668 10480 8720 10532
rect 9036 10480 9088 10532
rect 10876 10480 10928 10532
rect 6368 10412 6420 10421
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 9772 10412 9824 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10416 10412 10468 10464
rect 10600 10412 10652 10464
rect 11336 10455 11388 10464
rect 11336 10421 11345 10455
rect 11345 10421 11379 10455
rect 11379 10421 11388 10455
rect 11336 10412 11388 10421
rect 11980 10412 12032 10464
rect 12900 10412 12952 10464
rect 14832 10616 14884 10668
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 13912 10480 13964 10532
rect 14372 10480 14424 10532
rect 14648 10480 14700 10532
rect 14740 10480 14792 10532
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 3700 10251 3752 10260
rect 3700 10217 3709 10251
rect 3709 10217 3743 10251
rect 3743 10217 3752 10251
rect 3700 10208 3752 10217
rect 4620 10208 4672 10260
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 2504 10140 2556 10192
rect 4896 10140 4948 10192
rect 9404 10208 9456 10260
rect 9680 10251 9732 10260
rect 9680 10217 9689 10251
rect 9689 10217 9723 10251
rect 9723 10217 9732 10251
rect 9680 10208 9732 10217
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 11336 10208 11388 10260
rect 12256 10208 12308 10260
rect 14372 10251 14424 10260
rect 1768 10072 1820 10124
rect 3056 10072 3108 10124
rect 3976 10072 4028 10124
rect 6828 10140 6880 10192
rect 7104 10140 7156 10192
rect 1860 10004 1912 10056
rect 6368 10004 6420 10056
rect 6644 10004 6696 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 5632 9936 5684 9988
rect 9036 10140 9088 10192
rect 10232 10140 10284 10192
rect 11796 10183 11848 10192
rect 11796 10149 11830 10183
rect 11830 10149 11848 10183
rect 11796 10140 11848 10149
rect 11888 10140 11940 10192
rect 12348 10140 12400 10192
rect 14372 10217 14381 10251
rect 14381 10217 14415 10251
rect 14415 10217 14424 10251
rect 14372 10208 14424 10217
rect 14648 10251 14700 10260
rect 14648 10217 14657 10251
rect 14657 10217 14691 10251
rect 14691 10217 14700 10251
rect 14648 10208 14700 10217
rect 14740 10208 14792 10260
rect 13268 10183 13320 10192
rect 13268 10149 13302 10183
rect 13302 10149 13320 10183
rect 13268 10140 13320 10149
rect 9680 10072 9732 10124
rect 9864 10072 9916 10124
rect 9956 10072 10008 10124
rect 10784 10072 10836 10124
rect 12164 10072 12216 10124
rect 8208 10004 8260 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 10048 10004 10100 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 8760 9979 8812 9988
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 5448 9868 5500 9877
rect 6644 9868 6696 9920
rect 8760 9945 8769 9979
rect 8769 9945 8803 9979
rect 8803 9945 8812 9979
rect 8760 9936 8812 9945
rect 9772 9936 9824 9988
rect 8852 9868 8904 9920
rect 9864 9868 9916 9920
rect 12532 9868 12584 9920
rect 13544 10072 13596 10124
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 4068 9664 4120 9716
rect 8208 9707 8260 9716
rect 3792 9596 3844 9648
rect 5356 9596 5408 9648
rect 6828 9596 6880 9648
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 9496 9664 9548 9716
rect 9680 9664 9732 9716
rect 10968 9664 11020 9716
rect 11796 9664 11848 9716
rect 8484 9596 8536 9648
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 4160 9528 4212 9580
rect 5448 9528 5500 9580
rect 5724 9528 5776 9580
rect 4252 9460 4304 9512
rect 5632 9460 5684 9512
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6460 9392 6512 9444
rect 7196 9392 7248 9444
rect 9956 9528 10008 9580
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 11244 9596 11296 9648
rect 11980 9571 12032 9580
rect 11980 9537 11989 9571
rect 11989 9537 12023 9571
rect 12023 9537 12032 9571
rect 11980 9528 12032 9537
rect 12900 9664 12952 9716
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 12992 9596 13044 9648
rect 13360 9596 13412 9648
rect 9772 9460 9824 9512
rect 11152 9460 11204 9512
rect 13268 9528 13320 9580
rect 15108 9528 15160 9580
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 5816 9324 5868 9376
rect 6184 9324 6236 9376
rect 7656 9324 7708 9376
rect 8208 9324 8260 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9404 9392 9456 9444
rect 9680 9324 9732 9376
rect 10416 9324 10468 9376
rect 11244 9324 11296 9376
rect 13084 9392 13136 9444
rect 16028 9392 16080 9444
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1768 9120 1820 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 7748 9120 7800 9172
rect 8208 9120 8260 9172
rect 9220 9120 9272 9172
rect 9496 9120 9548 9172
rect 10968 9120 11020 9172
rect 11152 9163 11204 9172
rect 11152 9129 11161 9163
rect 11161 9129 11195 9163
rect 11195 9129 11204 9163
rect 11152 9120 11204 9129
rect 11888 9120 11940 9172
rect 12532 9120 12584 9172
rect 12992 9120 13044 9172
rect 4068 9052 4120 9104
rect 2044 8984 2096 9036
rect 3516 8984 3568 9036
rect 5540 8984 5592 9036
rect 5724 8984 5776 9036
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 8484 8984 8536 9036
rect 8944 8984 8996 9036
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 9956 9027 10008 9036
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 5816 8959 5868 8968
rect 1860 8848 1912 8900
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 9956 8993 9990 9027
rect 9990 8993 10008 9027
rect 9956 8984 10008 8993
rect 13820 9052 13872 9104
rect 14740 9052 14792 9104
rect 11152 8984 11204 9036
rect 9680 8959 9732 8968
rect 7196 8891 7248 8900
rect 7196 8857 7205 8891
rect 7205 8857 7239 8891
rect 7239 8857 7248 8891
rect 7196 8848 7248 8857
rect 7104 8780 7156 8832
rect 7840 8780 7892 8832
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 10876 8916 10928 8968
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 10968 8848 11020 8900
rect 11888 8848 11940 8900
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 13636 9027 13688 9036
rect 12440 8984 12492 8993
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 12992 8916 13044 8968
rect 9864 8780 9916 8832
rect 10048 8780 10100 8832
rect 10784 8780 10836 8832
rect 11244 8780 11296 8832
rect 13084 8780 13136 8832
rect 13268 8823 13320 8832
rect 13268 8789 13277 8823
rect 13277 8789 13311 8823
rect 13311 8789 13320 8823
rect 13268 8780 13320 8789
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 5264 8576 5316 8628
rect 5356 8576 5408 8628
rect 4160 8508 4212 8560
rect 6920 8576 6972 8628
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 11244 8576 11296 8628
rect 12440 8576 12492 8628
rect 5908 8508 5960 8560
rect 9404 8508 9456 8560
rect 9496 8508 9548 8560
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 3148 8372 3200 8424
rect 2780 8236 2832 8288
rect 3424 8304 3476 8356
rect 4252 8372 4304 8424
rect 5080 8372 5132 8424
rect 5816 8372 5868 8424
rect 5540 8304 5592 8356
rect 6368 8440 6420 8492
rect 8300 8440 8352 8492
rect 9772 8483 9824 8492
rect 7104 8372 7156 8424
rect 7472 8372 7524 8424
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10416 8440 10468 8492
rect 10600 8508 10652 8560
rect 11152 8508 11204 8560
rect 11888 8508 11940 8560
rect 17224 8576 17276 8628
rect 13452 8508 13504 8560
rect 9496 8372 9548 8424
rect 9864 8372 9916 8424
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 5356 8236 5408 8288
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 8300 8304 8352 8356
rect 8668 8304 8720 8356
rect 9036 8304 9088 8356
rect 7196 8279 7248 8288
rect 7196 8245 7205 8279
rect 7205 8245 7239 8279
rect 7239 8245 7248 8279
rect 7196 8236 7248 8245
rect 8392 8236 8444 8288
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 9128 8236 9180 8288
rect 11980 8440 12032 8492
rect 12440 8483 12492 8492
rect 12440 8449 12449 8483
rect 12449 8449 12483 8483
rect 12483 8449 12492 8483
rect 12440 8440 12492 8449
rect 12808 8440 12860 8492
rect 12992 8440 13044 8492
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 13636 8440 13688 8449
rect 12532 8372 12584 8424
rect 15568 8372 15620 8424
rect 12624 8347 12676 8356
rect 12624 8313 12633 8347
rect 12633 8313 12667 8347
rect 12667 8313 12676 8347
rect 12624 8304 12676 8313
rect 13452 8304 13504 8356
rect 14372 8304 14424 8356
rect 14648 8304 14700 8356
rect 13084 8236 13136 8288
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 15660 8279 15712 8288
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 2504 8032 2556 8084
rect 2688 8032 2740 8084
rect 5448 8032 5500 8084
rect 5540 8032 5592 8084
rect 7288 8032 7340 8084
rect 1860 7964 1912 8016
rect 6092 7964 6144 8016
rect 2780 7896 2832 7948
rect 3148 7760 3200 7812
rect 4068 7896 4120 7948
rect 8300 7964 8352 8016
rect 6460 7896 6512 7948
rect 6920 7896 6972 7948
rect 7472 7896 7524 7948
rect 10784 7964 10836 8016
rect 10876 7964 10928 8016
rect 12992 7964 13044 8016
rect 15016 7964 15068 8016
rect 16764 7964 16816 8016
rect 9680 7896 9732 7948
rect 12532 7896 12584 7948
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 15476 7896 15528 7948
rect 15844 7896 15896 7948
rect 4160 7760 4212 7812
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 5540 7828 5592 7880
rect 6092 7828 6144 7880
rect 6368 7828 6420 7880
rect 6644 7871 6696 7880
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 7656 7828 7708 7880
rect 5724 7760 5776 7812
rect 6552 7760 6604 7812
rect 5080 7692 5132 7744
rect 6368 7692 6420 7744
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7196 7692 7248 7744
rect 8668 7692 8720 7744
rect 9220 7692 9272 7744
rect 9496 7692 9548 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 13912 7692 13964 7744
rect 14372 7828 14424 7880
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 16120 7760 16172 7812
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 3240 7488 3292 7540
rect 4068 7488 4120 7540
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 5264 7488 5316 7540
rect 6460 7488 6512 7540
rect 9128 7488 9180 7540
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 14648 7488 14700 7540
rect 15016 7531 15068 7540
rect 15016 7497 15025 7531
rect 15025 7497 15059 7531
rect 15059 7497 15068 7531
rect 15016 7488 15068 7497
rect 3332 7420 3384 7472
rect 8760 7420 8812 7472
rect 3148 7352 3200 7404
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6736 7352 6788 7404
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 11888 7420 11940 7472
rect 14740 7420 14792 7472
rect 10324 7352 10376 7404
rect 12348 7352 12400 7404
rect 12716 7352 12768 7404
rect 13084 7352 13136 7404
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 5908 7284 5960 7336
rect 7012 7284 7064 7336
rect 2412 7148 2464 7200
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 5172 7216 5224 7268
rect 3884 7148 3936 7157
rect 5264 7148 5316 7200
rect 6460 7216 6512 7268
rect 11244 7284 11296 7336
rect 11612 7284 11664 7336
rect 13268 7284 13320 7336
rect 15568 7327 15620 7336
rect 15568 7293 15602 7327
rect 15602 7293 15620 7327
rect 7748 7259 7800 7268
rect 7748 7225 7782 7259
rect 7782 7225 7800 7259
rect 7748 7216 7800 7225
rect 11060 7216 11112 7268
rect 8300 7148 8352 7200
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 11612 7148 11664 7200
rect 12348 7216 12400 7268
rect 13912 7216 13964 7268
rect 15568 7284 15620 7293
rect 15476 7216 15528 7268
rect 12532 7148 12584 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 4344 6944 4396 6996
rect 7748 6944 7800 6996
rect 8300 6987 8352 6996
rect 2872 6808 2924 6860
rect 3516 6851 3568 6860
rect 3516 6817 3525 6851
rect 3525 6817 3559 6851
rect 3559 6817 3568 6851
rect 3516 6808 3568 6817
rect 4988 6876 5040 6928
rect 6000 6919 6052 6928
rect 6000 6885 6009 6919
rect 6009 6885 6043 6919
rect 6043 6885 6052 6919
rect 6000 6876 6052 6885
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8392 6944 8444 6996
rect 9772 6944 9824 6996
rect 2780 6740 2832 6792
rect 4896 6808 4948 6860
rect 5080 6808 5132 6860
rect 6736 6851 6788 6860
rect 3976 6740 4028 6792
rect 5356 6740 5408 6792
rect 6736 6817 6770 6851
rect 6770 6817 6788 6851
rect 6736 6808 6788 6817
rect 11612 6944 11664 6996
rect 12348 6944 12400 6996
rect 12440 6944 12492 6996
rect 13820 6987 13872 6996
rect 13820 6953 13829 6987
rect 13829 6953 13863 6987
rect 13863 6953 13872 6987
rect 13820 6944 13872 6953
rect 6460 6783 6512 6792
rect 2044 6715 2096 6724
rect 2044 6681 2053 6715
rect 2053 6681 2087 6715
rect 2087 6681 2096 6715
rect 2044 6672 2096 6681
rect 4896 6672 4948 6724
rect 5908 6672 5960 6724
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 8576 6808 8628 6860
rect 11796 6876 11848 6928
rect 10232 6808 10284 6860
rect 10324 6783 10376 6792
rect 6368 6672 6420 6724
rect 3332 6604 3384 6656
rect 8944 6672 8996 6724
rect 7564 6604 7616 6656
rect 9220 6604 9272 6656
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 11980 6808 12032 6860
rect 14648 6808 14700 6860
rect 17592 6808 17644 6860
rect 14556 6783 14608 6792
rect 10876 6740 10928 6749
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 13084 6672 13136 6724
rect 15200 6672 15252 6724
rect 11980 6604 12032 6656
rect 15752 6604 15804 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 3056 6400 3108 6452
rect 3608 6400 3660 6452
rect 4068 6400 4120 6452
rect 4160 6332 4212 6384
rect 5172 6332 5224 6384
rect 1860 6239 1912 6248
rect 1860 6205 1869 6239
rect 1869 6205 1903 6239
rect 1903 6205 1912 6239
rect 1860 6196 1912 6205
rect 3148 6264 3200 6316
rect 3976 6307 4028 6316
rect 3976 6273 3985 6307
rect 3985 6273 4019 6307
rect 4019 6273 4028 6307
rect 3976 6264 4028 6273
rect 4896 6264 4948 6316
rect 6368 6400 6420 6452
rect 6736 6332 6788 6384
rect 12348 6400 12400 6452
rect 14464 6400 14516 6452
rect 14832 6400 14884 6452
rect 17684 6400 17736 6452
rect 10416 6332 10468 6384
rect 7656 6307 7708 6316
rect 7656 6273 7665 6307
rect 7665 6273 7699 6307
rect 7699 6273 7708 6307
rect 7656 6264 7708 6273
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 4160 6196 4212 6248
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 5356 6196 5408 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 9956 6196 10008 6248
rect 4068 6128 4120 6180
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 7748 6060 7800 6112
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9404 6128 9456 6180
rect 10324 6128 10376 6180
rect 11060 6196 11112 6248
rect 11428 6196 11480 6248
rect 15200 6375 15252 6384
rect 15200 6341 15209 6375
rect 15209 6341 15243 6375
rect 15243 6341 15252 6375
rect 15200 6332 15252 6341
rect 15936 6332 15988 6384
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 10232 6060 10284 6112
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 10968 6060 11020 6112
rect 13084 6128 13136 6180
rect 13912 6196 13964 6248
rect 14464 6196 14516 6248
rect 14648 6196 14700 6248
rect 16028 6196 16080 6248
rect 14188 6128 14240 6180
rect 17408 6128 17460 6180
rect 14280 6060 14332 6112
rect 14556 6060 14608 6112
rect 15292 6103 15344 6112
rect 15292 6069 15301 6103
rect 15301 6069 15335 6103
rect 15335 6069 15344 6103
rect 15292 6060 15344 6069
rect 15384 6060 15436 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3516 5856 3568 5908
rect 4712 5856 4764 5908
rect 4896 5856 4948 5908
rect 5264 5856 5316 5908
rect 5540 5856 5592 5908
rect 5908 5856 5960 5908
rect 6092 5899 6144 5908
rect 6092 5865 6101 5899
rect 6101 5865 6135 5899
rect 6135 5865 6144 5899
rect 6092 5856 6144 5865
rect 7472 5856 7524 5908
rect 8392 5856 8444 5908
rect 8484 5856 8536 5908
rect 10784 5856 10836 5908
rect 10968 5856 11020 5908
rect 14188 5856 14240 5908
rect 14740 5856 14792 5908
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 17684 5856 17736 5908
rect 4068 5788 4120 5840
rect 1860 5720 1912 5772
rect 8208 5788 8260 5840
rect 4712 5763 4764 5772
rect 4712 5729 4721 5763
rect 4721 5729 4755 5763
rect 4755 5729 4764 5763
rect 4712 5720 4764 5729
rect 5264 5720 5316 5772
rect 5356 5720 5408 5772
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 7656 5584 7708 5636
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9680 5788 9732 5840
rect 9947 5831 9999 5840
rect 9947 5797 9979 5831
rect 9979 5797 9999 5831
rect 9947 5788 9999 5797
rect 11888 5788 11940 5840
rect 9772 5720 9824 5772
rect 11152 5720 11204 5772
rect 11244 5720 11296 5772
rect 13084 5788 13136 5840
rect 14556 5763 14608 5772
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9312 5584 9364 5636
rect 11980 5652 12032 5704
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 11428 5584 11480 5636
rect 14372 5584 14424 5636
rect 15476 5652 15528 5704
rect 16028 5695 16080 5704
rect 16028 5661 16037 5695
rect 16037 5661 16071 5695
rect 16071 5661 16080 5695
rect 16028 5652 16080 5661
rect 17040 5584 17092 5636
rect 6736 5516 6788 5568
rect 7104 5516 7156 5568
rect 7748 5516 7800 5568
rect 12440 5516 12492 5568
rect 14004 5559 14056 5568
rect 14004 5525 14013 5559
rect 14013 5525 14047 5559
rect 14047 5525 14056 5559
rect 14004 5516 14056 5525
rect 14648 5516 14700 5568
rect 17500 5559 17552 5568
rect 17500 5525 17509 5559
rect 17509 5525 17543 5559
rect 17543 5525 17552 5559
rect 17500 5516 17552 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 3792 5312 3844 5364
rect 4804 5312 4856 5364
rect 6000 5312 6052 5364
rect 6920 5312 6972 5364
rect 7656 5312 7708 5364
rect 8208 5312 8260 5364
rect 11152 5355 11204 5364
rect 11152 5321 11161 5355
rect 11161 5321 11195 5355
rect 11195 5321 11204 5355
rect 11152 5312 11204 5321
rect 3976 5244 4028 5296
rect 6368 5244 6420 5296
rect 8484 5244 8536 5296
rect 4068 5176 4120 5228
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 6920 5176 6972 5228
rect 10416 5244 10468 5296
rect 11980 5312 12032 5364
rect 14096 5312 14148 5364
rect 14188 5312 14240 5364
rect 17040 5312 17092 5364
rect 17776 5355 17828 5364
rect 17776 5321 17785 5355
rect 17785 5321 17819 5355
rect 17819 5321 17828 5355
rect 17776 5312 17828 5321
rect 9680 5176 9732 5228
rect 18144 5244 18196 5296
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 2688 5108 2740 5160
rect 6644 5108 6696 5160
rect 6736 5108 6788 5160
rect 7288 5108 7340 5160
rect 9404 5108 9456 5160
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 11796 5176 11848 5185
rect 14648 5176 14700 5228
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 16672 5176 16724 5228
rect 13084 5151 13136 5160
rect 2964 5040 3016 5092
rect 3056 4972 3108 5024
rect 3700 4972 3752 5024
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5540 4972 5592 5024
rect 6828 5040 6880 5092
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13176 5108 13228 5160
rect 10416 5040 10468 5092
rect 11060 5040 11112 5092
rect 6276 5015 6328 5024
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6644 4972 6696 5024
rect 6736 4972 6788 5024
rect 8944 4972 8996 5024
rect 9588 4972 9640 5024
rect 10048 4972 10100 5024
rect 11152 4972 11204 5024
rect 11888 4972 11940 5024
rect 12256 5015 12308 5024
rect 12256 4981 12265 5015
rect 12265 4981 12299 5015
rect 12299 4981 12308 5015
rect 12256 4972 12308 4981
rect 13544 4972 13596 5024
rect 13728 5040 13780 5092
rect 15200 5040 15252 5092
rect 15752 5083 15804 5092
rect 15752 5049 15786 5083
rect 15786 5049 15804 5083
rect 15752 5040 15804 5049
rect 16672 5040 16724 5092
rect 17776 5040 17828 5092
rect 19984 5040 20036 5092
rect 14004 4972 14056 5024
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 16948 5015 17000 5024
rect 14556 4972 14608 4981
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17224 4972 17276 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 3424 4811 3476 4820
rect 1676 4700 1728 4752
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 5264 4768 5316 4820
rect 7380 4768 7432 4820
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 11888 4768 11940 4820
rect 13176 4768 13228 4820
rect 13728 4811 13780 4820
rect 13728 4777 13737 4811
rect 13737 4777 13771 4811
rect 13771 4777 13780 4811
rect 13728 4768 13780 4777
rect 3332 4743 3384 4752
rect 3332 4709 3341 4743
rect 3341 4709 3375 4743
rect 3375 4709 3384 4743
rect 3332 4700 3384 4709
rect 15200 4768 15252 4820
rect 15292 4768 15344 4820
rect 1400 4564 1452 4616
rect 3148 4632 3200 4684
rect 2780 4564 2832 4616
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 14556 4700 14608 4752
rect 16948 4768 17000 4820
rect 17500 4768 17552 4820
rect 4712 4632 4764 4684
rect 5448 4632 5500 4684
rect 6920 4632 6972 4684
rect 7656 4675 7708 4684
rect 7656 4641 7665 4675
rect 7665 4641 7699 4675
rect 7699 4641 7708 4675
rect 7656 4632 7708 4641
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 7012 4564 7064 4616
rect 8208 4564 8260 4616
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 8760 4607 8812 4616
rect 8760 4573 8769 4607
rect 8769 4573 8803 4607
rect 8803 4573 8812 4607
rect 8760 4564 8812 4573
rect 10784 4632 10836 4684
rect 11060 4632 11112 4684
rect 6184 4496 6236 4548
rect 9220 4496 9272 4548
rect 4160 4428 4212 4480
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 7012 4428 7064 4480
rect 10416 4607 10468 4616
rect 10416 4573 10425 4607
rect 10425 4573 10459 4607
rect 10459 4573 10468 4607
rect 10416 4564 10468 4573
rect 11980 4632 12032 4684
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 13636 4632 13688 4684
rect 14280 4632 14332 4684
rect 11796 4607 11848 4616
rect 11796 4573 11805 4607
rect 11805 4573 11839 4607
rect 11839 4573 11848 4607
rect 11796 4564 11848 4573
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 12808 4564 12860 4616
rect 13820 4564 13872 4616
rect 14188 4607 14240 4616
rect 14188 4573 14197 4607
rect 14197 4573 14231 4607
rect 14231 4573 14240 4607
rect 14188 4564 14240 4573
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 10140 4428 10192 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 19984 4675 20036 4684
rect 19984 4641 19993 4675
rect 19993 4641 20027 4675
rect 20027 4641 20036 4675
rect 19984 4632 20036 4641
rect 14556 4564 14608 4616
rect 17040 4564 17092 4616
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 12716 4428 12768 4480
rect 12900 4428 12952 4480
rect 15752 4496 15804 4548
rect 15016 4428 15068 4480
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 17132 4428 17184 4480
rect 20812 4428 20864 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2780 4224 2832 4276
rect 4068 4224 4120 4276
rect 6184 4224 6236 4276
rect 6276 4224 6328 4276
rect 4804 4156 4856 4208
rect 5080 4156 5132 4208
rect 5540 4156 5592 4208
rect 6920 4224 6972 4276
rect 8484 4224 8536 4276
rect 10232 4224 10284 4276
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 1860 4063 1912 4072
rect 1860 4029 1869 4063
rect 1869 4029 1903 4063
rect 1903 4029 1912 4063
rect 3332 4063 3384 4072
rect 1860 4020 1912 4029
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 4712 4088 4764 4140
rect 6184 4088 6236 4140
rect 6828 4088 6880 4140
rect 6920 4088 6972 4140
rect 4068 4020 4120 4072
rect 2044 3952 2096 4004
rect 1124 3884 1176 3936
rect 4160 3952 4212 4004
rect 8208 4131 8260 4140
rect 7104 4020 7156 4072
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 8760 4156 8812 4208
rect 9128 4088 9180 4140
rect 10140 4088 10192 4140
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 11060 4156 11112 4208
rect 11796 4156 11848 4208
rect 9404 4020 9456 4072
rect 2504 3884 2556 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6000 3884 6052 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 6552 3884 6604 3936
rect 7472 3884 7524 3936
rect 8576 3952 8628 4004
rect 8484 3884 8536 3936
rect 10048 3952 10100 4004
rect 10140 3952 10192 4004
rect 11980 4020 12032 4072
rect 13636 4224 13688 4276
rect 13820 4224 13872 4276
rect 14372 4224 14424 4276
rect 12256 4156 12308 4208
rect 13268 4156 13320 4208
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 15016 4088 15068 4140
rect 22652 4088 22704 4140
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 8944 3884 8996 3936
rect 10876 3884 10928 3936
rect 12808 3952 12860 4004
rect 13912 3995 13964 4004
rect 13912 3961 13946 3995
rect 13946 3961 13964 3995
rect 13912 3952 13964 3961
rect 14280 3952 14332 4004
rect 17132 4063 17184 4072
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 18052 3952 18104 4004
rect 11888 3884 11940 3936
rect 12256 3884 12308 3936
rect 13820 3884 13872 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 204 3680 256 3732
rect 2780 3680 2832 3732
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 3424 3680 3476 3732
rect 3056 3612 3108 3664
rect 3332 3612 3384 3664
rect 1768 3544 1820 3596
rect 2780 3544 2832 3596
rect 3608 3587 3660 3596
rect 3608 3553 3617 3587
rect 3617 3553 3651 3587
rect 3651 3553 3660 3587
rect 4712 3612 4764 3664
rect 4896 3612 4948 3664
rect 5448 3680 5500 3732
rect 9772 3723 9824 3732
rect 5632 3612 5684 3664
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 10048 3680 10100 3732
rect 10876 3680 10928 3732
rect 3608 3544 3660 3553
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 6736 3544 6788 3596
rect 7472 3612 7524 3664
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 7656 3544 7708 3596
rect 10140 3612 10192 3664
rect 10968 3612 11020 3664
rect 8852 3587 8904 3596
rect 8852 3553 8861 3587
rect 8861 3553 8895 3587
rect 8895 3553 8904 3587
rect 8852 3544 8904 3553
rect 8944 3544 8996 3596
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 2044 3340 2096 3392
rect 6184 3408 6236 3460
rect 6828 3451 6880 3460
rect 6828 3417 6837 3451
rect 6837 3417 6871 3451
rect 6871 3417 6880 3451
rect 6828 3408 6880 3417
rect 6920 3408 6972 3460
rect 6736 3340 6788 3392
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 8760 3476 8812 3528
rect 10048 3476 10100 3528
rect 10140 3408 10192 3460
rect 11428 3544 11480 3596
rect 10324 3476 10376 3528
rect 11704 3476 11756 3528
rect 11796 3476 11848 3528
rect 13084 3680 13136 3732
rect 13636 3680 13688 3732
rect 14188 3680 14240 3732
rect 15568 3612 15620 3664
rect 12523 3587 12575 3596
rect 12523 3553 12532 3587
rect 12532 3553 12566 3587
rect 12566 3553 12575 3587
rect 12523 3544 12575 3553
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 15660 3544 15712 3596
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 13820 3476 13872 3528
rect 13912 3408 13964 3460
rect 16396 3476 16448 3528
rect 8116 3340 8168 3392
rect 9772 3340 9824 3392
rect 11888 3340 11940 3392
rect 13360 3340 13412 3392
rect 14004 3340 14056 3392
rect 14280 3340 14332 3392
rect 20168 3408 20220 3460
rect 18972 3340 19024 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 3608 3179 3660 3188
rect 2780 3136 2832 3145
rect 3608 3145 3617 3179
rect 3617 3145 3651 3179
rect 3651 3145 3660 3179
rect 3608 3136 3660 3145
rect 4896 3136 4948 3188
rect 1676 3068 1728 3120
rect 7104 3136 7156 3188
rect 1584 3000 1636 3052
rect 2688 3000 2740 3052
rect 3056 3000 3108 3052
rect 1492 2932 1544 2984
rect 2596 2864 2648 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 1952 2796 2004 2805
rect 3056 2796 3108 2848
rect 4252 2932 4304 2984
rect 5540 3068 5592 3120
rect 5908 3068 5960 3120
rect 8484 3136 8536 3188
rect 8760 3136 8812 3188
rect 5448 3000 5500 3052
rect 6092 3000 6144 3052
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 5540 2932 5592 2984
rect 5632 2932 5684 2984
rect 7288 3000 7340 3052
rect 7472 2932 7524 2984
rect 8208 2932 8260 2984
rect 9312 3136 9364 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 11796 3136 11848 3188
rect 12532 3136 12584 3188
rect 13820 3179 13872 3188
rect 10048 2932 10100 2984
rect 12072 2932 12124 2984
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 15292 3068 15344 3120
rect 14372 2932 14424 2984
rect 22192 3136 22244 3188
rect 16580 3068 16632 3120
rect 17960 3068 18012 3120
rect 18144 3068 18196 3120
rect 19432 3068 19484 3120
rect 20352 3068 20404 3120
rect 16120 3000 16172 3052
rect 15384 2932 15436 2984
rect 15568 2932 15620 2984
rect 16028 2975 16080 2984
rect 16028 2941 16037 2975
rect 16037 2941 16071 2975
rect 16071 2941 16080 2975
rect 16028 2932 16080 2941
rect 16396 2975 16448 2984
rect 16396 2941 16405 2975
rect 16405 2941 16439 2975
rect 16439 2941 16448 2975
rect 16396 2932 16448 2941
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 17224 2975 17276 2984
rect 17224 2941 17233 2975
rect 17233 2941 17267 2975
rect 17267 2941 17276 2975
rect 17224 2932 17276 2941
rect 17316 2932 17368 2984
rect 17592 2975 17644 2984
rect 17592 2941 17601 2975
rect 17601 2941 17635 2975
rect 17635 2941 17644 2975
rect 17592 2932 17644 2941
rect 17776 2932 17828 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 18144 2932 18196 2984
rect 19064 2975 19116 2984
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 4344 2864 4396 2916
rect 5356 2864 5408 2916
rect 6736 2864 6788 2916
rect 3700 2796 3752 2848
rect 4160 2796 4212 2848
rect 6920 2796 6972 2848
rect 7748 2864 7800 2916
rect 10140 2864 10192 2916
rect 10324 2864 10376 2916
rect 10600 2864 10652 2916
rect 11152 2864 11204 2916
rect 13912 2864 13964 2916
rect 12716 2796 12768 2848
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 14740 2839 14792 2848
rect 12808 2796 12860 2805
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 15200 2796 15252 2848
rect 15660 2796 15712 2848
rect 16120 2796 16172 2848
rect 17040 2864 17092 2916
rect 17500 2796 17552 2848
rect 18144 2796 18196 2848
rect 19892 2864 19944 2916
rect 21272 2796 21324 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 1400 2635 1452 2644
rect 1400 2601 1409 2635
rect 1409 2601 1443 2635
rect 1443 2601 1452 2635
rect 1400 2592 1452 2601
rect 1952 2592 2004 2644
rect 2596 2635 2648 2644
rect 2596 2601 2605 2635
rect 2605 2601 2639 2635
rect 2639 2601 2648 2635
rect 2596 2592 2648 2601
rect 3700 2635 3752 2644
rect 3700 2601 3709 2635
rect 3709 2601 3743 2635
rect 3743 2601 3752 2635
rect 3700 2592 3752 2601
rect 4160 2592 4212 2644
rect 5080 2592 5132 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 6092 2592 6144 2644
rect 8852 2592 8904 2644
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 10416 2592 10468 2644
rect 10600 2592 10652 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 11980 2592 12032 2644
rect 14096 2592 14148 2644
rect 15384 2592 15436 2644
rect 15844 2592 15896 2644
rect 16028 2592 16080 2644
rect 16764 2592 16816 2644
rect 17224 2592 17276 2644
rect 17316 2592 17368 2644
rect 18052 2592 18104 2644
rect 19064 2592 19116 2644
rect 2688 2524 2740 2576
rect 7104 2524 7156 2576
rect 9404 2524 9456 2576
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 4068 2456 4120 2508
rect 5724 2456 5776 2508
rect 6644 2456 6696 2508
rect 10232 2524 10284 2576
rect 12716 2524 12768 2576
rect 9956 2456 10008 2508
rect 12440 2456 12492 2508
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 2872 2320 2924 2372
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 7748 2388 7800 2440
rect 10600 2431 10652 2440
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 5356 2295 5408 2304
rect 5356 2261 5365 2295
rect 5365 2261 5399 2295
rect 5399 2261 5408 2295
rect 5356 2252 5408 2261
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11152 2320 11204 2372
rect 11704 2388 11756 2440
rect 13268 2252 13320 2304
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 14280 2252 14332 2304
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 2044 2048 2096 2100
rect 6644 2048 6696 2100
rect 15752 2048 15804 2100
rect 21732 2048 21784 2100
rect 664 1980 716 2032
rect 6552 1980 6604 2032
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3054 22672 3110 22681
rect 3054 22607 3110 22616
rect 216 16697 244 22200
rect 676 18630 704 22200
rect 1136 18902 1164 22200
rect 1596 21298 1624 22200
rect 1596 21270 1900 21298
rect 1582 21176 1638 21185
rect 1582 21111 1638 21120
rect 1596 20058 1624 21111
rect 1674 20768 1730 20777
rect 1674 20703 1730 20712
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1582 19816 1638 19825
rect 1582 19751 1638 19760
rect 1596 18970 1624 19751
rect 1688 19514 1716 20703
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1676 19508 1728 19514
rect 1676 19450 1728 19456
rect 1780 19378 1808 20334
rect 1768 19372 1820 19378
rect 1768 19314 1820 19320
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1124 18896 1176 18902
rect 1124 18838 1176 18844
rect 1582 18864 1638 18873
rect 1400 18828 1452 18834
rect 1582 18799 1638 18808
rect 1766 18864 1822 18873
rect 1766 18799 1768 18808
rect 1400 18770 1452 18776
rect 664 18624 716 18630
rect 664 18566 716 18572
rect 1412 18086 1440 18770
rect 1596 18426 1624 18799
rect 1820 18799 1822 18808
rect 1768 18770 1820 18776
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1768 18216 1820 18222
rect 1872 18193 1900 21270
rect 1950 20224 2006 20233
rect 1950 20159 2006 20168
rect 1964 20058 1992 20159
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 1964 18970 1992 19207
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2056 18737 2084 22200
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 2148 18902 2176 20334
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2240 19514 2268 19858
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 2516 19394 2544 22200
rect 2870 22128 2926 22137
rect 2870 22063 2926 22072
rect 2778 21720 2834 21729
rect 2778 21655 2834 21664
rect 2792 20602 2820 21655
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2884 20534 2912 22063
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2516 19366 2728 19394
rect 2504 19304 2556 19310
rect 2700 19281 2728 19366
rect 2792 19310 2820 19790
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2884 19378 2912 19722
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2780 19304 2832 19310
rect 2504 19246 2556 19252
rect 2686 19272 2742 19281
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2042 18728 2098 18737
rect 2042 18663 2098 18672
rect 2516 18426 2544 19246
rect 2596 19236 2648 19242
rect 2780 19246 2832 19252
rect 2686 19207 2742 19216
rect 2596 19178 2648 19184
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 1952 18352 2004 18358
rect 1950 18320 1952 18329
rect 2004 18320 2006 18329
rect 2608 18290 2636 19178
rect 2976 19009 3004 22200
rect 2962 19000 3018 19009
rect 2962 18935 3018 18944
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 1950 18255 2006 18264
rect 2596 18284 2648 18290
rect 2596 18226 2648 18232
rect 1768 18158 1820 18164
rect 1858 18184 1914 18193
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 16776 1440 18022
rect 1674 17912 1730 17921
rect 1674 17847 1730 17856
rect 1582 17368 1638 17377
rect 1688 17338 1716 17847
rect 1780 17814 1808 18158
rect 1858 18119 1914 18128
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 2504 17740 2556 17746
rect 2504 17682 2556 17688
rect 1582 17303 1638 17312
rect 1676 17332 1728 17338
rect 1596 16794 1624 17303
rect 1676 17274 1728 17280
rect 1584 16788 1636 16794
rect 1412 16748 1532 16776
rect 202 16688 258 16697
rect 1504 16674 1532 16748
rect 1584 16730 1636 16736
rect 1872 16726 1900 17682
rect 2516 17105 2544 17682
rect 2502 17096 2558 17105
rect 2502 17031 2558 17040
rect 2136 16992 2188 16998
rect 1950 16960 2006 16969
rect 2136 16934 2188 16940
rect 1950 16895 2006 16904
rect 1964 16794 1992 16895
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1860 16720 1912 16726
rect 202 16623 258 16632
rect 1400 16652 1452 16658
rect 1504 16646 1624 16674
rect 1860 16662 1912 16668
rect 2148 16658 2176 16934
rect 1400 16594 1452 16600
rect 1412 16114 1440 16594
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1492 11620 1544 11626
rect 1492 11562 1544 11568
rect 1504 10690 1532 11562
rect 1596 10810 1624 16646
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 1780 15502 1808 16594
rect 1950 16416 2006 16425
rect 1950 16351 2006 16360
rect 1964 16250 1992 16351
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2700 15910 2728 18566
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2792 17814 2820 18090
rect 2780 17808 2832 17814
rect 3068 17762 3096 22607
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 2780 17750 2832 17756
rect 2976 17734 3096 17762
rect 2976 17610 3004 17734
rect 2964 17604 3016 17610
rect 2964 17546 3016 17552
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3068 17202 3096 17546
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 16794 3004 16934
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2778 16008 2834 16017
rect 2778 15943 2834 15952
rect 2872 15972 2924 15978
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2792 15706 2820 15943
rect 2872 15914 2924 15920
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1950 15056 2006 15065
rect 1950 14991 2006 15000
rect 1964 14618 1992 14991
rect 2332 14958 2360 15506
rect 2778 15464 2834 15473
rect 2778 15399 2834 15408
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2792 14618 2820 15399
rect 2884 15026 2912 15914
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 1858 14512 1914 14521
rect 1858 14447 1914 14456
rect 2136 14476 2188 14482
rect 1872 14074 1900 14447
rect 2136 14418 2188 14424
rect 2044 14340 2096 14346
rect 2044 14282 2096 14288
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1504 10662 1624 10690
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1124 3936 1176 3942
rect 1124 3878 1176 3884
rect 204 3732 256 3738
rect 204 3674 256 3680
rect 216 800 244 3674
rect 664 2032 716 2038
rect 664 1974 716 1980
rect 676 800 704 1974
rect 1136 800 1164 3878
rect 1412 2650 1440 4558
rect 1504 3398 1532 10406
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 2990 1532 3334
rect 1596 3058 1624 10662
rect 1688 4758 1716 13806
rect 1766 13560 1822 13569
rect 1766 13495 1768 13504
rect 1820 13495 1822 13504
rect 1768 13466 1820 13472
rect 2056 12782 2084 14282
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 2056 12306 2084 12718
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1964 11354 1992 11494
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1780 9178 1808 10066
rect 1872 10062 1900 10542
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1872 8906 1900 9998
rect 2148 9586 2176 14418
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 13870 2360 14350
rect 2778 14104 2834 14113
rect 2778 14039 2780 14048
rect 2832 14039 2834 14048
rect 2780 14010 2832 14016
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2240 11762 2268 12650
rect 2332 11898 2360 13330
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2424 12850 2452 13262
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 2332 11218 2360 11630
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 10470 2360 11154
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2516 10198 2544 13806
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12646 2636 13262
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 2884 12782 2912 13126
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 10606 2636 12582
rect 2976 11626 3004 13670
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 11762 3096 12242
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8498 1900 8842
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1872 6254 1900 7958
rect 2056 6730 2084 8978
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2516 8090 2544 8910
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2424 7002 2452 7142
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5778 1900 6190
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1872 5166 1900 5714
rect 2700 5166 2728 8026
rect 2792 7954 2820 8230
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2792 6798 2820 7890
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 6866 2912 7686
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2780 6792 2832 6798
rect 2976 6746 3004 11222
rect 3068 11150 3096 11698
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3160 10554 3188 17478
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3252 16726 3280 17138
rect 3436 16998 3464 22200
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 16046 3556 16390
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3896 15858 3924 22200
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3988 18426 4016 18566
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3988 17134 4016 18362
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4080 17134 4108 17274
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16250 4108 17070
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3896 15830 4016 15858
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3344 14074 3372 14758
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3252 11898 3280 13330
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12986 3372 13262
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3436 11694 3464 15506
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14074 3648 14758
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3528 12714 3556 13262
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3528 12442 3556 12650
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3620 11286 3648 12378
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3700 11144 3752 11150
rect 3700 11086 3752 11092
rect 3608 10600 3660 10606
rect 3160 10526 3372 10554
rect 3608 10542 3660 10548
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2780 6734 2832 6740
rect 2884 6718 3004 6746
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1872 4078 1900 5102
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2792 4282 2820 4558
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2778 4176 2834 4185
rect 2778 4111 2834 4120
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1768 3596 1820 3602
rect 1872 3584 1900 4014
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1820 3556 1900 3584
rect 1768 3538 1820 3544
rect 2056 3398 2084 3946
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 1504 2145 1532 2926
rect 1596 2854 1624 2994
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1490 2136 1546 2145
rect 1490 2071 1546 2080
rect 1596 1193 1624 2790
rect 1582 1184 1638 1193
rect 1582 1119 1638 1128
rect 1688 1034 1716 3062
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1964 2650 1992 2790
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2056 2446 2084 3334
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 1596 1006 1716 1034
rect 1596 800 1624 1006
rect 2056 800 2084 2042
rect 2516 800 2544 3878
rect 2792 3738 2820 4111
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2792 3194 2820 3538
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2884 3097 2912 6718
rect 3068 6458 3096 10066
rect 3160 8430 3188 10406
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 7818 3188 8366
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3160 7410 3188 7754
rect 3252 7546 3280 8910
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3344 7478 3372 10526
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3436 8362 3464 8910
rect 3528 8634 3556 8978
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3332 7472 3384 7478
rect 3332 7414 3384 7420
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3344 6746 3372 7414
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3252 6718 3372 6746
rect 3056 6452 3108 6458
rect 3056 6394 3108 6400
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3160 5914 3188 6258
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2870 3088 2926 3097
rect 2688 3052 2740 3058
rect 2870 3023 2926 3032
rect 2688 2994 2740 3000
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2608 2650 2636 2858
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2700 2582 2728 2994
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2884 2378 2912 3023
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2976 800 3004 5034
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3068 3670 3096 4966
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 3738 3188 4626
rect 3252 4604 3280 6718
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3344 4758 3372 6598
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 4826 3464 6054
rect 3528 5914 3556 6802
rect 3620 6610 3648 10542
rect 3712 10266 3740 11086
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3804 9654 3832 14826
rect 3896 14618 3924 14962
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3896 13938 3924 14418
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 3896 13734 3924 13767
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3896 12617 3924 12854
rect 3988 12782 4016 15830
rect 4172 15586 4200 19858
rect 4252 18760 4304 18766
rect 4252 18702 4304 18708
rect 4264 18426 4292 18702
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4356 17882 4384 22200
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4540 20058 4568 20334
rect 4528 20052 4580 20058
rect 4528 19994 4580 20000
rect 4816 19938 4844 22200
rect 4816 19910 5028 19938
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4724 19310 4752 19382
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4618 19136 4674 19145
rect 4618 19071 4674 19080
rect 4632 18970 4660 19071
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4724 18834 4752 19246
rect 4816 19242 4844 19790
rect 4908 19514 4936 19790
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4816 18970 4844 19178
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4816 18193 4844 18362
rect 4908 18290 4936 18566
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4802 18184 4858 18193
rect 4802 18119 4858 18128
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4448 17762 4476 18022
rect 4356 17734 4476 17762
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4264 15706 4292 16594
rect 4356 16130 4384 17734
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 17338 4844 17614
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4816 16590 4844 17070
rect 4908 16794 4936 17274
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4356 16102 4476 16130
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4356 15586 4384 15642
rect 4172 15570 4384 15586
rect 4160 15564 4384 15570
rect 4212 15558 4384 15564
rect 4160 15506 4212 15512
rect 4448 15450 4476 16102
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4632 15502 4660 15914
rect 4264 15422 4476 15450
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 4080 13734 4108 14214
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13394 4108 13670
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3882 12200 3938 12209
rect 3882 12135 3938 12144
rect 3896 11694 3924 12135
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3988 11121 4016 11766
rect 4080 11762 4108 12786
rect 4264 12442 4292 15422
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4252 12300 4304 12306
rect 4172 12260 4252 12288
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4066 11656 4122 11665
rect 4066 11591 4122 11600
rect 4080 11286 4108 11591
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3974 11112 4030 11121
rect 3974 11047 4030 11056
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10713 4016 10950
rect 3974 10704 4030 10713
rect 3884 10668 3936 10674
rect 3974 10639 4030 10648
rect 3884 10610 3936 10616
rect 3896 10470 3924 10610
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3896 8294 3924 10406
rect 3974 10160 4030 10169
rect 3974 10095 3976 10104
rect 4028 10095 4030 10104
rect 3976 10066 4028 10072
rect 4066 9752 4122 9761
rect 4066 9687 4068 9696
rect 4120 9687 4122 9696
rect 4068 9658 4120 9664
rect 4172 9586 4200 12260
rect 4252 12242 4304 12248
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4264 11558 4292 11698
rect 4252 11552 4304 11558
rect 4304 11512 4384 11540
rect 4252 11494 4304 11500
rect 4356 10690 4384 11512
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4356 10662 4476 10690
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4264 9518 4292 10406
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4066 9208 4122 9217
rect 4066 9143 4122 9152
rect 4080 9110 4108 9143
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 4080 7857 4108 7890
rect 4066 7848 4122 7857
rect 4172 7818 4200 8502
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4066 7783 4122 7792
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4080 7313 4108 7482
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3620 6582 3740 6610
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3514 5400 3570 5409
rect 3514 5335 3570 5344
rect 3528 4865 3556 5335
rect 3514 4856 3570 4865
rect 3424 4820 3476 4826
rect 3514 4791 3570 4800
rect 3424 4762 3476 4768
rect 3332 4752 3384 4758
rect 3332 4694 3384 4700
rect 3620 4622 3648 6394
rect 3712 5030 3740 6582
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5370 3832 6054
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3608 4616 3660 4622
rect 3252 4576 3372 4604
rect 3344 4162 3372 4576
rect 3608 4558 3660 4564
rect 3252 4134 3372 4162
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 3068 3058 3096 3606
rect 3252 3505 3280 4134
rect 3332 4072 3384 4078
rect 3712 4049 3740 4966
rect 3332 4014 3384 4020
rect 3698 4040 3754 4049
rect 3344 3670 3372 4014
rect 3698 3975 3754 3984
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3068 2310 3096 2790
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3068 241 3096 2246
rect 3436 800 3464 3674
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3620 3194 3648 3538
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3712 2854 3740 2885
rect 3700 2848 3752 2854
rect 3698 2816 3700 2825
rect 3752 2816 3754 2825
rect 3698 2751 3754 2760
rect 3712 2650 3740 2751
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3896 800 3924 7142
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3988 6322 4016 6734
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4080 6361 4108 6394
rect 4172 6390 4200 7754
rect 4264 7750 4292 8366
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 6384 4212 6390
rect 4066 6352 4122 6361
rect 3976 6316 4028 6322
rect 4160 6326 4212 6332
rect 4066 6287 4122 6296
rect 3976 6258 4028 6264
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 5953 4108 6122
rect 4066 5944 4122 5953
rect 4066 5879 4122 5888
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3988 5001 4016 5238
rect 4080 5234 4108 5782
rect 4172 5574 4200 6190
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 4172 4486 4200 5510
rect 4160 4480 4212 4486
rect 4066 4448 4122 4457
rect 4160 4422 4212 4428
rect 4066 4383 4122 4392
rect 4080 4282 4108 4383
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3505 4108 4014
rect 4172 4010 4200 4422
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 4264 2990 4292 7686
rect 4356 7546 4384 10474
rect 4448 10033 4476 10662
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 10266 4660 10406
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4434 10024 4490 10033
rect 4434 9959 4490 9968
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4356 7002 4384 7482
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4724 5778 4752 5850
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4816 5370 4844 13806
rect 4908 11626 4936 16458
rect 5000 12986 5028 19910
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 5092 19145 5120 19178
rect 5078 19136 5134 19145
rect 5078 19071 5134 19080
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5092 16522 5120 18158
rect 5276 18154 5304 22200
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5552 18290 5580 20198
rect 5736 19145 5764 22200
rect 6196 19904 6224 22200
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6288 19922 6316 20402
rect 6656 20346 6684 22200
rect 7116 20602 7144 22200
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6472 20318 6684 20346
rect 6828 20324 6880 20330
rect 5920 19876 6224 19904
rect 6276 19916 6328 19922
rect 5722 19136 5778 19145
rect 5722 19071 5778 19080
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5736 18290 5764 18838
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5276 17882 5304 18090
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17882 5396 18022
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 5276 16250 5304 16594
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5552 15162 5580 15574
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5736 15094 5764 15982
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13734 5580 14350
rect 5736 13870 5764 15030
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5644 13530 5672 13806
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 4988 12980 5040 12986
rect 5040 12940 5212 12968
rect 4988 12922 5040 12928
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 5092 11762 5120 12038
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 4896 11620 4948 11626
rect 4896 11562 4948 11568
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4908 10198 4936 10610
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4894 10024 4950 10033
rect 4894 9959 4950 9968
rect 4908 6866 4936 9959
rect 5000 6934 5028 11018
rect 5092 8430 5120 11562
rect 5184 9636 5212 12940
rect 5552 12442 5580 13398
rect 5828 13258 5856 13874
rect 5816 13252 5868 13258
rect 5816 13194 5868 13200
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5276 11150 5304 12174
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5368 11354 5396 11494
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5276 10674 5304 11086
rect 5460 10810 5488 11494
rect 5920 10826 5948 19876
rect 6276 19858 6328 19864
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 6196 19310 6224 19722
rect 6288 19514 6316 19858
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6274 19272 6330 19281
rect 6274 19207 6330 19216
rect 5998 19000 6054 19009
rect 5998 18935 6054 18944
rect 6012 18698 6040 18935
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 6288 18154 6316 19207
rect 6380 18902 6408 19654
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6276 18148 6328 18154
rect 6276 18090 6328 18096
rect 6472 17898 6500 20318
rect 6828 20266 6880 20272
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5552 10798 5948 10826
rect 6012 17870 6500 17898
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5356 9648 5408 9654
rect 5184 9608 5356 9636
rect 5356 9590 5408 9596
rect 5460 9586 5488 9862
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5276 8634 5304 9318
rect 5368 8634 5396 9318
rect 5552 9160 5580 10798
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9518 5672 9930
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5736 9178 5764 9522
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5724 9172 5776 9178
rect 5552 9132 5672 9160
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5552 8362 5580 8978
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5356 8288 5408 8294
rect 5262 8256 5318 8265
rect 5356 8230 5408 8236
rect 5262 8191 5318 8200
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 7256 5120 7686
rect 5276 7546 5304 8191
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5172 7268 5224 7274
rect 5092 7228 5172 7256
rect 5172 7210 5224 7216
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4908 6322 4936 6666
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4712 4684 4764 4690
rect 4908 4672 4936 5850
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4764 4644 4936 4672
rect 4712 4626 4764 4632
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4724 3942 4752 4082
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4724 3670 4752 3878
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4816 3074 4844 4150
rect 4908 3670 4936 4644
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 4896 3188 4948 3194
rect 5000 3176 5028 4966
rect 5092 4214 5120 6802
rect 5184 6474 5212 7210
rect 5264 7200 5316 7206
rect 5262 7168 5264 7177
rect 5316 7168 5318 7177
rect 5368 7154 5396 8230
rect 5552 8090 5580 8298
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5460 7970 5488 8026
rect 5460 7942 5580 7970
rect 5552 7886 5580 7942
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5368 7126 5580 7154
rect 5262 7103 5318 7112
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5184 6446 5304 6474
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5078 4040 5134 4049
rect 5078 3975 5134 3984
rect 4948 3148 5028 3176
rect 4896 3130 4948 3136
rect 4816 3046 4936 3074
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4172 2650 4200 2790
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4066 2544 4122 2553
rect 4066 2479 4068 2488
rect 4120 2479 4122 2488
rect 4068 2450 4120 2456
rect 4356 800 4384 2858
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4908 800 4936 3046
rect 5092 2650 5120 3975
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5184 2310 5212 6326
rect 5276 6254 5304 6446
rect 5368 6254 5396 6734
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5276 5914 5304 6190
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5368 5778 5396 6190
rect 5552 5914 5580 7126
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5276 5234 5304 5714
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5276 4826 5304 5170
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5460 3738 5488 4626
rect 5552 4214 5580 4966
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5644 4049 5672 9132
rect 5724 9114 5776 9120
rect 5736 9042 5764 9114
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5828 8974 5856 9318
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5814 8800 5870 8809
rect 5814 8735 5870 8744
rect 5828 8430 5856 8735
rect 5920 8566 5948 9454
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5630 4040 5686 4049
rect 5630 3975 5686 3984
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5460 3058 5488 3674
rect 5552 3126 5580 3878
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5644 2990 5672 3606
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5368 2310 5396 2858
rect 5552 2650 5580 2926
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5736 2514 5764 7754
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5184 1601 5212 2246
rect 5170 1592 5226 1601
rect 5170 1527 5226 1536
rect 5368 800 5396 2246
rect 5828 800 5856 8366
rect 5920 7342 5948 8502
rect 6012 8106 6040 17870
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6472 17202 6500 17682
rect 6564 17678 6592 20198
rect 6840 20058 6868 20266
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 7024 19922 7052 20198
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6932 18834 6960 19314
rect 6920 18828 6972 18834
rect 6920 18770 6972 18776
rect 6932 17762 6960 18770
rect 6840 17734 6960 17762
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14618 6408 14758
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 12714 6132 13806
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 11898 6224 12242
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 11014 6500 11086
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10266 6408 10406
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6274 10160 6330 10169
rect 6274 10095 6330 10104
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 8809 6224 9318
rect 6182 8800 6238 8809
rect 6182 8735 6238 8744
rect 6012 8078 6224 8106
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6104 7886 6132 7958
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 5906 6760 5962 6769
rect 5906 6695 5908 6704
rect 5960 6695 5962 6704
rect 5908 6666 5960 6672
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5920 5250 5948 5850
rect 6012 5370 6040 6870
rect 6104 5914 6132 7822
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6196 5522 6224 8078
rect 6104 5494 6224 5522
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5920 5222 6040 5250
rect 6012 3942 6040 5222
rect 6104 4049 6132 5494
rect 6288 5114 6316 10095
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 8616 6408 9998
rect 6472 9450 6500 10950
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 6380 8588 6500 8616
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6380 7886 6408 8434
rect 6472 7954 6500 8588
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7410 6408 7686
rect 6472 7546 6500 7890
rect 6564 7818 6592 17614
rect 6840 17202 6868 17734
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6656 15162 6684 16934
rect 6748 16522 6776 17002
rect 6932 16794 6960 17070
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6840 16250 6868 16662
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6932 14958 6960 15506
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14346 6960 14894
rect 7024 14822 7052 19858
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19310 7328 19654
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7392 19174 7420 19790
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7392 18902 7420 19110
rect 7380 18896 7432 18902
rect 7380 18838 7432 18844
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 16794 7144 17478
rect 7392 17134 7420 17614
rect 7380 17128 7432 17134
rect 7286 17096 7342 17105
rect 7196 17060 7248 17066
rect 7380 17070 7432 17076
rect 7286 17031 7342 17040
rect 7196 17002 7248 17008
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7208 16454 7236 17002
rect 7300 16726 7328 17031
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 7392 16590 7420 16934
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 16182 7236 16390
rect 7196 16176 7248 16182
rect 7248 16124 7328 16130
rect 7196 16118 7328 16124
rect 7208 16102 7328 16118
rect 7300 15638 7328 16102
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7208 15366 7236 15506
rect 7300 15502 7328 15574
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 15026 7236 15302
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 7024 14278 7052 14758
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 11626 6776 13194
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12646 6868 12718
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12442 6868 12582
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7024 12288 7052 14214
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13530 7144 13670
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6932 12260 7052 12288
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6840 11354 6868 11630
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10674 6776 11154
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6748 10180 6776 10610
rect 6828 10192 6880 10198
rect 6748 10152 6828 10180
rect 6828 10134 6880 10140
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9926 6684 9998
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6656 8294 6684 9862
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7886 6684 8230
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6472 6798 6500 7210
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6380 6458 6408 6666
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6472 5710 6500 6734
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6656 5522 6684 7822
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 6866 6776 7346
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 6390 6776 6802
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6380 5494 6684 5522
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6380 5302 6408 5494
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6748 5166 6776 5510
rect 6644 5160 6696 5166
rect 6288 5086 6408 5114
rect 6644 5102 6696 5108
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6196 4282 6224 4490
rect 6288 4282 6316 4966
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6090 4040 6146 4049
rect 6090 3975 6146 3984
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5920 3126 5948 3878
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6104 3058 6132 3975
rect 6196 3466 6224 4082
rect 6380 4060 6408 5086
rect 6656 5030 6684 5102
rect 6840 5098 6868 9590
rect 6932 8634 6960 12260
rect 7116 12220 7144 12718
rect 7208 12374 7236 13874
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7300 12442 7328 13126
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7024 12192 7144 12220
rect 7024 12102 7052 12192
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7024 11762 7052 12038
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7116 11694 7144 12038
rect 7392 11898 7420 15574
rect 7576 12730 7604 22200
rect 8036 20754 8064 22200
rect 7668 20726 8064 20754
rect 7668 14634 7696 20726
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7760 20058 7788 20538
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8128 19514 8156 19790
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7748 18352 7800 18358
rect 7748 18294 7800 18300
rect 7760 15638 7788 18294
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8128 17066 8156 17138
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8220 16590 8248 17070
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8220 15638 8248 15846
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7668 14606 7788 14634
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7484 12702 7604 12730
rect 7484 12481 7512 12702
rect 7668 12594 7696 14418
rect 7576 12566 7696 12594
rect 7470 12472 7526 12481
rect 7470 12407 7526 12416
rect 7470 12336 7526 12345
rect 7470 12271 7526 12280
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 7024 10810 7052 11494
rect 7288 11280 7340 11286
rect 7288 11222 7340 11228
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 7116 10198 7144 10678
rect 7300 10470 7328 11222
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7102 8936 7158 8945
rect 7208 8906 7236 9386
rect 7102 8871 7158 8880
rect 7196 8900 7248 8906
rect 7116 8838 7144 8871
rect 7196 8842 7248 8848
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7116 8430 7144 8774
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7410 6960 7890
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7024 7342 7052 7686
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7116 5574 7144 8366
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7750 7236 8230
rect 7300 8090 7328 10406
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6932 5234 6960 5306
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6288 4032 6408 4060
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6196 3058 6224 3402
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6104 2650 6132 2994
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6196 2446 6224 2994
rect 6288 2825 6316 4032
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6380 3602 6408 3878
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6274 2816 6330 2825
rect 6274 2751 6330 2760
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6288 800 6316 2751
rect 3054 232 3110 241
rect 3054 167 3110 176
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6380 649 6408 3538
rect 6564 2038 6592 3878
rect 6656 2514 6684 4966
rect 6748 4865 6776 4966
rect 6734 4856 6790 4865
rect 6734 4791 6790 4800
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4486 6960 4626
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7024 4486 7052 4558
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6932 4282 6960 4422
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 7024 4185 7052 4422
rect 7010 4176 7066 4185
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6920 4140 6972 4146
rect 7010 4111 7066 4120
rect 6920 4082 6972 4088
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6748 3398 6776 3538
rect 6840 3466 6868 4082
rect 6932 4026 6960 4082
rect 7104 4072 7156 4078
rect 6932 4020 7104 4026
rect 6932 4014 7156 4020
rect 6932 3998 7144 4014
rect 6828 3460 6880 3466
rect 6828 3402 6880 3408
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 2922 6776 3334
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6656 2106 6684 2450
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6748 800 6776 2858
rect 6932 2854 6960 3402
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 7116 2582 7144 3130
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7208 800 7236 7686
rect 7392 6769 7420 11562
rect 7484 8430 7512 12271
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7484 7954 7512 8366
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7576 7834 7604 12566
rect 7760 12458 7788 14606
rect 8312 13977 8340 19994
rect 8496 19394 8524 22200
rect 8956 20398 8984 22200
rect 8944 20392 8996 20398
rect 8944 20334 8996 20340
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8404 19366 8524 19394
rect 8680 19378 8708 19926
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8668 19372 8720 19378
rect 8298 13968 8354 13977
rect 8298 13903 8354 13912
rect 7840 13864 7892 13870
rect 7838 13832 7840 13841
rect 8024 13864 8076 13870
rect 7892 13832 7894 13841
rect 8076 13824 8248 13852
rect 8024 13806 8076 13812
rect 7838 13767 7894 13776
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7840 13320 7892 13326
rect 7892 13280 7972 13308
rect 7840 13262 7892 13268
rect 7944 12918 7972 13280
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 8220 12782 8248 13824
rect 8298 13832 8354 13841
rect 8298 13767 8354 13776
rect 8312 13530 8340 13767
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13258 8432 19366
rect 8668 19314 8720 19320
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8496 18970 8524 19246
rect 9036 19236 9088 19242
rect 9036 19178 9088 19184
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8482 16688 8538 16697
rect 8482 16623 8538 16632
rect 8496 14822 8524 16623
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8680 15706 8708 15914
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 13326 8524 14758
rect 8680 13530 8708 15438
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8208 12640 8260 12646
rect 8208 12582 8260 12588
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7668 12430 7788 12458
rect 7668 9382 7696 12430
rect 8220 12238 8248 12582
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 8680 12102 8708 13466
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10538 8248 11154
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10606 8340 10950
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7748 10056 7800 10062
rect 8208 10056 8260 10062
rect 7748 9998 7800 10004
rect 7838 10024 7894 10033
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7760 9178 7788 9998
rect 8208 9998 8260 10004
rect 7838 9959 7894 9968
rect 7852 9489 7880 9959
rect 8220 9722 8248 9998
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8220 9178 8248 9318
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8220 9081 8248 9114
rect 8206 9072 8262 9081
rect 8024 9036 8076 9042
rect 8206 9007 8262 9016
rect 8024 8978 8076 8984
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8430 7880 8774
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 8036 8276 8064 8978
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 8362 8340 8434
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8036 8248 8248 8276
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7484 7806 7604 7834
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7378 6760 7434 6769
rect 7378 6695 7434 6704
rect 7484 6225 7512 7806
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7300 3058 7328 5102
rect 7392 4826 7420 6054
rect 7484 5914 7512 6054
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3670 7512 3878
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7472 2984 7524 2990
rect 7576 2972 7604 6598
rect 7668 6322 7696 7822
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7760 7002 7788 7210
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 8220 6882 8248 8248
rect 8312 8022 8340 8298
rect 8404 8294 8432 11766
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 11354 8708 11698
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8482 10568 8538 10577
rect 8482 10503 8538 10512
rect 8496 9654 8524 10503
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8484 9376 8536 9382
rect 8588 9364 8616 10950
rect 8680 10538 8708 11290
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8666 10432 8722 10441
rect 8666 10367 8722 10376
rect 8536 9336 8616 9364
rect 8484 9318 8536 9324
rect 8496 9042 8524 9318
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8673 8524 8774
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8680 8480 8708 10367
rect 8772 9994 8800 18770
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8864 17814 8892 18022
rect 8852 17808 8904 17814
rect 8852 17750 8904 17756
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8864 15910 8892 16186
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8864 13172 8892 15846
rect 8956 15162 8984 18566
rect 9048 15706 9076 19178
rect 9324 19174 9352 19858
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9324 18766 9352 19110
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17882 9260 18022
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 16794 9168 17682
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9048 15502 9076 15642
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 9220 15088 9272 15094
rect 9220 15030 9272 15036
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9036 14952 9088 14958
rect 9036 14894 9088 14900
rect 9048 14618 9076 14894
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8956 13326 8984 13874
rect 9140 13512 9168 14962
rect 9232 14890 9260 15030
rect 9220 14884 9272 14890
rect 9220 14826 9272 14832
rect 9416 14482 9444 22200
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9600 20058 9628 20198
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9692 18970 9720 19654
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 17134 9628 17478
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9692 16794 9720 18022
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9784 17338 9812 17682
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9876 16250 9904 22200
rect 10336 19802 10364 22200
rect 10796 20602 10824 22200
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10060 19774 10364 19802
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9968 17746 9996 18226
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 17338 9996 17682
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10060 16658 10088 19774
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10336 19310 10364 19654
rect 11072 19514 11100 19858
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10414 18864 10470 18873
rect 10414 18799 10470 18808
rect 10876 18828 10928 18834
rect 10428 18766 10456 18799
rect 10876 18770 10928 18776
rect 10416 18760 10468 18766
rect 10322 18728 10378 18737
rect 10416 18702 10468 18708
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10322 18663 10378 18672
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9048 13484 9168 13512
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8864 13144 8984 13172
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11762 8892 12038
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8956 11642 8984 13144
rect 9048 12442 9076 13484
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9048 11830 9076 12378
rect 9036 11824 9088 11830
rect 9036 11766 9088 11772
rect 8864 11614 8984 11642
rect 8864 10441 8892 11614
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8850 10432 8906 10441
rect 8850 10367 8906 10376
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8496 8452 8708 8480
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8312 7290 8340 7958
rect 8312 7262 8432 7290
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 7002 8340 7142
rect 8404 7002 8432 7262
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8220 6854 8340 6882
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 5642 7696 6258
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5681 7788 6054
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 7746 5672 7802 5681
rect 7656 5636 7708 5642
rect 7746 5607 7802 5616
rect 7656 5578 7708 5584
rect 7668 5370 7696 5578
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7668 3602 7696 4626
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7760 3482 7788 5510
rect 8220 5370 8248 5782
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8220 4622 8248 5306
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7524 2944 7604 2972
rect 7668 3454 7788 3482
rect 7472 2926 7524 2932
rect 7668 800 7696 3454
rect 8128 3398 8156 3606
rect 8220 3534 8248 4082
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8220 2990 8248 3470
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 7760 2446 7788 2858
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8312 2632 8340 6854
rect 8496 6202 8524 8452
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8680 7750 8708 8298
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8864 8242 8892 9862
rect 8956 9042 8984 11018
rect 9048 10538 9076 11766
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 10198 9076 10474
rect 9036 10192 9088 10198
rect 9036 10134 9088 10140
rect 9140 9160 9168 13330
rect 9232 11286 9260 14418
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9324 13326 9352 14010
rect 9508 13802 9536 14962
rect 9876 14958 9904 15098
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9416 13172 9444 13466
rect 9324 13144 9444 13172
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9232 11082 9260 11222
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 9178 9260 9998
rect 9048 9132 9168 9160
rect 9220 9172 9272 9178
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 9048 8362 9076 9132
rect 9220 9114 9272 9120
rect 9128 9036 9180 9042
rect 9180 8996 9260 9024
rect 9128 8978 9180 8984
rect 9232 8634 9260 8996
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9128 8288 9180 8294
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8574 6896 8630 6905
rect 8574 6831 8576 6840
rect 8628 6831 8630 6840
rect 8576 6802 8628 6808
rect 8404 6174 8524 6202
rect 8404 5914 8432 6174
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8496 5914 8524 6054
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8404 5794 8432 5850
rect 8404 5766 8524 5794
rect 8392 5704 8444 5710
rect 8390 5672 8392 5681
rect 8444 5672 8446 5681
rect 8390 5607 8446 5616
rect 8496 5302 8524 5766
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8496 4282 8524 4626
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8588 4010 8616 4558
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8484 3936 8536 3942
rect 8680 3890 8708 7686
rect 8772 7478 8800 8230
rect 8864 8214 9076 8242
rect 9128 8230 9180 8236
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6322 8984 6666
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8772 4214 8800 4558
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8484 3878 8536 3884
rect 8496 3194 8524 3878
rect 8588 3862 8708 3890
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8128 2604 8340 2632
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8128 800 8156 2604
rect 8588 800 8616 3862
rect 8772 3534 8800 4150
rect 8956 3942 8984 4966
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8942 3632 8998 3641
rect 8852 3596 8904 3602
rect 8942 3567 8944 3576
rect 8852 3538 8904 3544
rect 8996 3567 8998 3576
rect 8944 3538 8996 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 3194 8800 3470
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8864 2650 8892 3538
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 9048 800 9076 8214
rect 9140 7546 9168 8230
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9140 4146 9168 7482
rect 9232 6662 9260 7686
rect 9324 7562 9352 13144
rect 9508 12306 9536 13738
rect 9692 13546 9720 14554
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 9876 13870 9904 14418
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9692 13530 9904 13546
rect 9588 13524 9640 13530
rect 9692 13524 9916 13530
rect 9692 13518 9864 13524
rect 9692 13512 9720 13518
rect 9640 13484 9720 13512
rect 9588 13466 9640 13472
rect 9864 13466 9916 13472
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9586 13288 9642 13297
rect 9586 13223 9642 13232
rect 9600 13190 9628 13223
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9784 12986 9812 13398
rect 9968 13002 9996 15574
rect 10060 13716 10088 16594
rect 10152 15638 10180 18362
rect 10336 17218 10364 18663
rect 10704 18222 10732 18702
rect 10888 18426 10916 18770
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10692 17808 10744 17814
rect 10692 17750 10744 17756
rect 10336 17190 10456 17218
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10244 14278 10272 16594
rect 10336 16590 10364 17070
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10428 15586 10456 17190
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10612 16590 10640 16730
rect 10704 16590 10732 17750
rect 10600 16584 10652 16590
rect 10598 16552 10600 16561
rect 10692 16584 10744 16590
rect 10652 16552 10654 16561
rect 10692 16526 10744 16532
rect 10598 16487 10654 16496
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10336 15558 10456 15586
rect 10336 14793 10364 15558
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14958 10456 15438
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10322 14784 10378 14793
rect 10322 14719 10378 14728
rect 10336 14482 10364 14719
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10244 13870 10272 14214
rect 10520 13977 10548 16390
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10704 15638 10732 16526
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10796 15042 10824 18090
rect 11072 17746 11100 19450
rect 11256 18714 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11440 18766 11468 19178
rect 11716 18952 11744 22200
rect 12176 20040 12204 22200
rect 12636 20058 12664 22200
rect 13096 20058 13124 22200
rect 13268 20324 13320 20330
rect 13268 20266 13320 20272
rect 13280 20058 13308 20266
rect 12624 20052 12676 20058
rect 12176 20012 12296 20040
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11716 18924 11928 18952
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11164 18686 11284 18714
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11164 16522 11192 18686
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11256 18222 11284 18566
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11716 18290 11744 18770
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11808 18222 11836 18566
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 15484 10916 16390
rect 11164 15994 11192 16458
rect 11256 16454 11284 17682
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11900 16998 11928 18924
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11348 16794 11376 16934
rect 11532 16794 11560 16934
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11992 16250 12020 19926
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 12176 19514 12204 19858
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12176 18358 12204 19450
rect 12268 18970 12296 20012
rect 12624 19994 12676 20000
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12452 18902 12480 19654
rect 12636 19378 12664 19858
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12440 18896 12492 18902
rect 12268 18844 12440 18850
rect 12268 18838 12492 18844
rect 12268 18822 12480 18838
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 12084 17202 12112 17750
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12084 16590 12112 17138
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 10980 15966 11192 15994
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 10980 15706 11008 15966
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11072 15706 11100 15846
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11060 15496 11112 15502
rect 10888 15456 11060 15484
rect 11060 15438 11112 15444
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10612 15014 10824 15042
rect 10876 15020 10928 15026
rect 10612 14482 10640 15014
rect 10876 14962 10928 14968
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10506 13968 10562 13977
rect 10506 13903 10562 13912
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10704 13802 10732 14826
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14550 10824 14758
rect 10888 14618 10916 14962
rect 10980 14890 11008 15302
rect 11072 15162 11100 15438
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10784 14544 10836 14550
rect 10980 14498 11008 14554
rect 10784 14486 10836 14492
rect 10888 14482 11008 14498
rect 10876 14476 11008 14482
rect 10928 14470 11008 14476
rect 10876 14418 10928 14424
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 13938 10824 14214
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10060 13688 10364 13716
rect 9772 12980 9824 12986
rect 9968 12974 10088 13002
rect 9772 12922 9824 12928
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9772 12368 9824 12374
rect 9876 12322 9904 12582
rect 9968 12374 9996 12854
rect 10060 12646 10088 12974
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10244 12481 10272 12582
rect 10230 12472 10286 12481
rect 10230 12407 10232 12416
rect 10284 12407 10286 12416
rect 10232 12378 10284 12384
rect 9824 12316 9904 12322
rect 9772 12310 9904 12316
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9496 12300 9548 12306
rect 9784 12294 9904 12310
rect 9496 12242 9548 12248
rect 9508 11558 9536 12242
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9416 10266 9444 10610
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9508 9722 9536 10950
rect 9600 10742 9628 11698
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9692 10266 9720 11562
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9692 9722 9720 10066
rect 9784 9994 9812 10406
rect 9876 10130 9904 12294
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9968 10130 9996 11834
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 10577 10088 11494
rect 10336 10690 10364 13688
rect 10796 13682 10824 13738
rect 10612 13654 10824 13682
rect 10612 12102 10640 13654
rect 10980 13326 11008 14470
rect 11072 13938 11100 14758
rect 11164 14074 11192 15846
rect 11256 15162 11284 15982
rect 11440 15638 11468 16050
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11716 15076 11744 15574
rect 11348 15048 11744 15076
rect 11348 14906 11376 15048
rect 11256 14878 11376 14906
rect 11256 14822 11284 14878
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14550 11376 14758
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11716 14482 11744 15048
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 11256 13818 11284 14282
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11072 13790 11284 13818
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10152 10662 10364 10690
rect 10046 10568 10102 10577
rect 10046 10503 10102 10512
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10266 10088 10406
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9784 9518 9812 9930
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9416 8566 9444 9386
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9508 9081 9536 9114
rect 9494 9072 9550 9081
rect 9494 9007 9550 9016
rect 9692 8974 9720 9318
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9586 8800 9642 8809
rect 9586 8735 9642 8744
rect 9404 8560 9456 8566
rect 9496 8560 9548 8566
rect 9404 8502 9456 8508
rect 9494 8528 9496 8537
rect 9548 8528 9550 8537
rect 9494 8463 9550 8472
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9508 7750 9536 8366
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9324 7534 9536 7562
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 4554 9260 6598
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5642 9352 6190
rect 9416 6186 9444 7142
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9324 3194 9352 5578
rect 9416 5166 9444 5646
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9416 2582 9444 4014
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9508 898 9536 7534
rect 9600 5030 9628 8735
rect 9692 7954 9720 8910
rect 9784 8498 9812 9454
rect 9876 8838 9904 9862
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9042 9996 9522
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 10060 8838 10088 9998
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9862 8664 9918 8673
rect 9862 8599 9918 8608
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9876 8430 9904 8599
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9784 7002 9812 7142
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9770 5944 9826 5953
rect 9770 5879 9826 5888
rect 9680 5840 9732 5846
rect 9678 5808 9680 5817
rect 9732 5808 9734 5817
rect 9784 5778 9812 5879
rect 9968 5846 9996 6190
rect 9947 5840 9999 5846
rect 9947 5782 9999 5788
rect 9678 5743 9734 5752
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9692 3097 9720 5170
rect 10152 5114 10180 10662
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10244 9654 10272 10134
rect 10336 10062 10364 10542
rect 10428 10470 10456 11018
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 10470 10640 10610
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10598 10160 10654 10169
rect 10598 10095 10654 10104
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10428 8498 10456 9318
rect 10612 8673 10640 10095
rect 10598 8664 10654 8673
rect 10598 8599 10654 8608
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10244 6118 10272 6802
rect 10336 6798 10364 7346
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 6186 10364 6734
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10232 6112 10284 6118
rect 10428 6066 10456 6326
rect 10232 6054 10284 6060
rect 9968 5086 10180 5114
rect 10336 6038 10456 6066
rect 9772 3732 9824 3738
rect 9968 3720 9996 5086
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4185 10088 4966
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10046 4176 10102 4185
rect 10152 4146 10180 4422
rect 10244 4282 10272 4626
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10336 4162 10364 6038
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 10428 5098 10456 5238
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10046 4111 10102 4120
rect 10140 4140 10192 4146
rect 10060 4010 10088 4111
rect 10140 4082 10192 4088
rect 10244 4134 10364 4162
rect 10152 4010 10180 4082
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 9824 3692 9996 3720
rect 10048 3732 10100 3738
rect 9772 3674 9824 3680
rect 10048 3674 10100 3680
rect 9784 3505 9812 3674
rect 10060 3618 10088 3674
rect 10140 3664 10192 3670
rect 9968 3590 10088 3618
rect 10138 3632 10140 3641
rect 10192 3632 10194 3641
rect 9770 3496 9826 3505
rect 9770 3431 9826 3440
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9784 3233 9812 3334
rect 9770 3224 9826 3233
rect 9770 3159 9826 3168
rect 9678 3088 9734 3097
rect 9678 3023 9734 3032
rect 9968 2514 9996 3590
rect 10138 3567 10194 3576
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10060 3369 10088 3470
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 10046 3360 10102 3369
rect 10046 3295 10102 3304
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 9508 870 9628 898
rect 9600 800 9628 870
rect 10060 800 10088 2926
rect 10152 2922 10180 3402
rect 10140 2916 10192 2922
rect 10140 2858 10192 2864
rect 10244 2582 10272 4134
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10336 3369 10364 3470
rect 10322 3360 10378 3369
rect 10322 3295 10378 3304
rect 10428 3194 10456 4558
rect 10612 4146 10640 8502
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10336 2650 10364 2858
rect 10428 2650 10456 3130
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10612 2650 10640 2858
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10612 2446 10640 2586
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 1442 10732 12718
rect 10796 12442 10824 12786
rect 10980 12782 11008 13262
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10796 11762 10824 12378
rect 10980 11778 11008 12718
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10888 11750 11008 11778
rect 10888 11626 10916 11750
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 10130 10824 10542
rect 10876 10532 10928 10538
rect 10876 10474 10928 10480
rect 10888 10266 10916 10474
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9722 11008 9998
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10784 8832 10836 8838
rect 10888 8809 10916 8910
rect 10980 8906 11008 9114
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10784 8774 10836 8780
rect 10874 8800 10930 8809
rect 10796 8022 10824 8774
rect 10874 8735 10930 8744
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10888 6798 10916 7958
rect 11072 7274 11100 13790
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13326 11560 13670
rect 11610 13424 11666 13433
rect 11610 13359 11612 13368
rect 11664 13359 11666 13368
rect 11612 13330 11664 13336
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11164 12764 11192 13262
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11244 12776 11296 12782
rect 11164 12736 11244 12764
rect 11164 12306 11192 12736
rect 11244 12718 11296 12724
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11440 12306 11468 12378
rect 11624 12345 11652 12650
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11610 12336 11666 12345
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 11428 12300 11480 12306
rect 11610 12271 11666 12280
rect 11428 12242 11480 12248
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11898 11744 12582
rect 11808 12102 11836 16186
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11900 12481 11928 14826
rect 11992 14414 12020 14962
rect 11980 14408 12032 14414
rect 11978 14376 11980 14385
rect 12032 14376 12034 14385
rect 11978 14311 12034 14320
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11886 12472 11942 12481
rect 11886 12407 11942 12416
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11900 11898 11928 12407
rect 11992 12186 12020 14214
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12850 12112 13330
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12268 12458 12296 18822
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12360 18426 12388 18702
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12452 18358 12480 18634
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12452 17746 12480 18158
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12544 17542 12572 18090
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12544 16590 12572 17478
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16046 12572 16390
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12544 15570 12572 15982
rect 12636 15706 12664 16050
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12544 14482 12572 14962
rect 12622 14512 12678 14521
rect 12532 14476 12584 14482
rect 12622 14447 12678 14456
rect 12532 14418 12584 14424
rect 12636 14278 12664 14447
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12728 13818 12756 19246
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12820 18630 12848 18906
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12912 17134 12940 19654
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12820 13954 12848 14486
rect 12912 14074 12940 17070
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12820 13926 12940 13954
rect 12636 13790 12756 13818
rect 12808 13796 12860 13802
rect 12636 13410 12664 13790
rect 12808 13738 12860 13744
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13530 12756 13670
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12636 13394 12756 13410
rect 12636 13388 12768 13394
rect 12636 13382 12716 13388
rect 12716 13330 12768 13336
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12268 12430 12388 12458
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 11992 12158 12204 12186
rect 12072 12096 12124 12102
rect 11992 12044 12072 12050
rect 11992 12038 12124 12044
rect 11992 12022 12112 12038
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11164 10606 11192 11766
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11256 9654 11284 11154
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11716 10810 11744 11494
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11702 10704 11758 10713
rect 11702 10639 11758 10648
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11348 10266 11376 10406
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11164 9178 11192 9454
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11152 9036 11204 9042
rect 11256 9024 11284 9318
rect 11204 8996 11284 9024
rect 11152 8978 11204 8984
rect 11164 8566 11192 8978
rect 11242 8936 11298 8945
rect 11242 8871 11298 8880
rect 11256 8838 11284 8871
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11256 7342 11284 8570
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11624 7206 11652 7278
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11624 7002 11652 7142
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 10784 6112 10836 6118
rect 10968 6112 11020 6118
rect 10784 6054 10836 6060
rect 10888 6060 10968 6066
rect 10888 6054 11020 6060
rect 10796 5914 10824 6054
rect 10888 6038 11008 6054
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5794 10916 6038
rect 10966 5944 11022 5953
rect 10966 5879 10968 5888
rect 11020 5879 11022 5888
rect 10968 5850 11020 5856
rect 10796 5766 10916 5794
rect 10796 4690 10824 5766
rect 11072 5098 11100 6190
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11164 5370 11192 5714
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 10796 2650 10824 4626
rect 11072 4486 11100 4626
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4214 11100 4422
rect 11164 4282 11192 4966
rect 11256 4826 11284 5714
rect 11440 5642 11468 6190
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11716 4706 11744 10639
rect 11808 10198 11836 11698
rect 11992 11150 12020 12022
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11900 10198 11928 11086
rect 11992 10470 12020 11086
rect 12176 10690 12204 12158
rect 12268 11150 12296 12242
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12084 10662 12204 10690
rect 12268 10674 12296 11086
rect 12256 10668 12308 10674
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11992 10146 12020 10406
rect 12084 10305 12112 10662
rect 12256 10610 12308 10616
rect 12360 10554 12388 12430
rect 12544 12102 12572 12718
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11762 12572 12038
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 12176 10526 12388 10554
rect 12070 10296 12126 10305
rect 12070 10231 12126 10240
rect 11808 9722 11836 10134
rect 11992 10118 12112 10146
rect 12176 10130 12204 10526
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11808 8974 11836 9658
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8566 11928 8842
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11992 8498 12020 9522
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11808 6934 11836 7686
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11808 5234 11836 6870
rect 11900 5846 11928 7414
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11992 6769 12020 6802
rect 11978 6760 12034 6769
rect 11978 6695 12034 6704
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11992 5710 12020 6598
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5370 12020 5646
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11256 4678 11744 4706
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10888 3738 10916 3878
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10980 2650 11008 3606
rect 11072 3233 11100 4150
rect 11058 3224 11114 3233
rect 11058 3159 11114 3168
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11164 2378 11192 2858
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11256 1442 11284 4678
rect 11808 4622 11836 5170
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4826 11928 4966
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11808 4214 11836 4558
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11900 3942 11928 4762
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11992 4078 12020 4626
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11440 3505 11468 3538
rect 11704 3528 11756 3534
rect 11426 3496 11482 3505
rect 11704 3470 11756 3476
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11426 3431 11482 3440
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11716 2446 11744 3470
rect 11808 3194 11836 3470
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 10704 1414 11008 1442
rect 11256 1414 11468 1442
rect 10506 912 10562 921
rect 10506 847 10562 856
rect 10520 800 10548 847
rect 10980 800 11008 1414
rect 11440 800 11468 1414
rect 11900 800 11928 3334
rect 11992 2650 12020 4014
rect 12084 2990 12112 10118
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12176 4842 12204 10066
rect 12268 7546 12296 10202
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12268 7290 12296 7482
rect 12360 7410 12388 10134
rect 12452 9654 12480 11154
rect 12636 11014 12664 13262
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12782 12756 13126
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12714 12336 12770 12345
rect 12714 12271 12770 12280
rect 12728 12238 12756 12271
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12544 9178 12572 9862
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12452 8634 12480 8978
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12268 7274 12388 7290
rect 12268 7268 12400 7274
rect 12268 7262 12348 7268
rect 12348 7210 12400 7216
rect 12452 7002 12480 8434
rect 12544 8430 12572 9114
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12544 7954 12572 8366
rect 12636 8362 12664 10950
rect 12820 8498 12848 13738
rect 12912 13530 12940 13926
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12912 11694 12940 13330
rect 13004 12442 13032 19246
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13372 17202 13400 17682
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13464 17082 13492 19178
rect 13556 19174 13584 22200
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13740 20058 13768 20198
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13372 17054 13492 17082
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13280 15570 13308 15642
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13188 14822 13216 15098
rect 13280 15026 13308 15506
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13096 14618 13124 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13188 14346 13216 14554
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13096 13734 13124 14214
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12992 12300 13044 12306
rect 13044 12260 13124 12288
rect 12992 12242 13044 12248
rect 13096 11898 13124 12260
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13188 11778 13216 14010
rect 13268 13864 13320 13870
rect 13372 13852 13400 17054
rect 13464 15014 13860 15042
rect 13464 14890 13492 15014
rect 13832 14958 13860 15014
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13452 14544 13504 14550
rect 13450 14512 13452 14521
rect 13504 14512 13506 14521
rect 13450 14447 13506 14456
rect 13556 14074 13584 14894
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14618 13768 14826
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13728 14408 13780 14414
rect 13648 14385 13728 14396
rect 13634 14376 13728 14385
rect 13690 14368 13728 14376
rect 13728 14350 13780 14356
rect 13634 14311 13690 14320
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13450 13968 13506 13977
rect 13450 13903 13452 13912
rect 13504 13903 13506 13912
rect 13452 13874 13504 13880
rect 13320 13824 13400 13852
rect 13268 13806 13320 13812
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13280 13433 13308 13670
rect 13266 13424 13322 13433
rect 13266 13359 13322 13368
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 13258 13400 13330
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13280 12238 13308 12718
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13096 11750 13216 11778
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11354 12940 11494
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 9722 12940 10406
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12992 9648 13044 9654
rect 13096 9625 13124 11750
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13280 10198 13308 10610
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 12992 9590 13044 9596
rect 13082 9616 13138 9625
rect 13004 9178 13032 9590
rect 13280 9586 13308 10134
rect 13372 9654 13400 13194
rect 13464 10169 13492 13874
rect 13648 13870 13676 14311
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13556 13530 13584 13806
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13648 13326 13676 13806
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13648 12986 13676 13262
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13740 12646 13768 12718
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13740 12306 13768 12582
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 11830 13768 12242
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10810 13768 11086
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13450 10160 13506 10169
rect 13556 10130 13584 10542
rect 13450 10095 13506 10104
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13082 9551 13138 9560
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13358 9480 13414 9489
rect 13084 9444 13136 9450
rect 13358 9415 13414 9424
rect 13084 9386 13136 9392
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8498 13032 8910
rect 13096 8838 13124 9386
rect 13372 9330 13400 9415
rect 13452 9376 13504 9382
rect 13372 9324 13452 9330
rect 13372 9318 13504 9324
rect 13372 9302 13492 9318
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 13004 8022 13032 8434
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12360 6458 12388 6938
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12544 6338 12572 7142
rect 12268 6310 12572 6338
rect 12268 5030 12296 6310
rect 12622 6216 12678 6225
rect 12622 6151 12678 6160
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12176 4814 12388 4842
rect 12256 4208 12308 4214
rect 12254 4176 12256 4185
rect 12308 4176 12310 4185
rect 12254 4111 12310 4120
rect 12254 4040 12310 4049
rect 12254 3975 12310 3984
rect 12268 3942 12296 3975
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12360 800 12388 4814
rect 12452 2514 12480 5510
rect 12523 3596 12575 3602
rect 12523 3538 12575 3544
rect 12544 3194 12572 3538
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12636 2394 12664 6151
rect 12728 4706 12756 7346
rect 13004 7290 13032 7958
rect 13096 7410 13124 8230
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13280 7342 13308 8774
rect 13268 7336 13320 7342
rect 13004 7262 13124 7290
rect 13268 7278 13320 7284
rect 13096 6730 13124 7262
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13096 6322 13124 6666
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 13096 5846 13124 6122
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13096 5166 13124 5782
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 12728 4678 12940 4706
rect 12728 4622 12756 4678
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12728 3890 12756 4422
rect 12820 4146 12848 4558
rect 12912 4486 12940 4678
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12820 4010 12848 4082
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12728 3862 12848 3890
rect 12820 2854 12848 3862
rect 13096 3738 13124 5102
rect 13188 4826 13216 5102
rect 13176 4820 13228 4826
rect 13176 4762 13228 4768
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4214 13308 4626
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13372 3398 13400 9302
rect 13832 9194 13860 12786
rect 13924 11354 13952 18770
rect 14016 17882 14044 22200
rect 14186 19408 14242 19417
rect 14242 19366 14320 19394
rect 14186 19343 14242 19352
rect 14292 19310 14320 19366
rect 14280 19304 14332 19310
rect 14476 19258 14504 22200
rect 14936 20346 14964 22200
rect 14752 20318 14964 20346
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14568 19553 14596 19654
rect 14554 19544 14610 19553
rect 14752 19530 14780 20318
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 14752 19502 14964 19530
rect 15396 19514 15424 22200
rect 14554 19479 14610 19488
rect 14280 19246 14332 19252
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18426 14136 18566
rect 14096 18420 14148 18426
rect 14096 18362 14148 18368
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 14108 15706 14136 15914
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14200 15434 14228 17070
rect 14188 15428 14240 15434
rect 14188 15370 14240 15376
rect 14004 15360 14056 15366
rect 14004 15302 14056 15308
rect 14016 12850 14044 15302
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14108 13716 14136 14894
rect 14200 14618 14228 15030
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14108 13688 14228 13716
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14108 11694 14136 13398
rect 14200 13258 14228 13688
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 12782 14228 13194
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14292 12424 14320 19246
rect 14384 19242 14504 19258
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14372 19236 14504 19242
rect 14424 19230 14504 19236
rect 14372 19178 14424 19184
rect 14752 18902 14780 19246
rect 14936 19242 14964 19502
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15660 19304 15712 19310
rect 15856 19258 15884 22200
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15660 19246 15712 19252
rect 14924 19236 14976 19242
rect 14924 19178 14976 19184
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14384 13870 14412 14418
rect 14476 14074 14504 18294
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14568 15162 14596 15506
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14660 14958 14688 15846
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14648 14952 14700 14958
rect 14700 14900 14780 14906
rect 14648 14894 14780 14900
rect 14660 14878 14780 14894
rect 14554 14784 14610 14793
rect 14554 14719 14610 14728
rect 14568 14550 14596 14719
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14752 14414 14780 14878
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 15120 13938 15148 14214
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14384 13530 14412 13806
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14200 12396 14320 12424
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14200 11626 14228 12396
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11354 14136 11494
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10538 13952 11086
rect 14292 11082 14320 12242
rect 14752 11762 14780 12718
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15212 12442 15240 18770
rect 15396 18630 15424 19246
rect 15672 18630 15700 19246
rect 15764 19230 15884 19258
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 15764 19174 15792 19230
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15948 18970 15976 19246
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 13938 15332 14758
rect 15396 14521 15424 18566
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15382 14512 15438 14521
rect 15382 14447 15438 14456
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 12850 15332 13874
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14384 10962 14412 11494
rect 14752 11234 14780 11698
rect 15212 11694 15240 12106
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15292 11620 15344 11626
rect 15292 11562 15344 11568
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14752 11206 14872 11234
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14292 10934 14412 10962
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13832 9166 14044 9194
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13464 8362 13492 8502
rect 13648 8498 13676 8978
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13832 7002 13860 9046
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13924 7410 13952 7686
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13924 6254 13952 7210
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14016 5658 14044 9166
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14200 5914 14228 6122
rect 14292 6118 14320 10934
rect 14752 10810 14780 11086
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14844 10674 14872 11206
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14384 10266 14412 10474
rect 14660 10266 14688 10474
rect 14752 10266 14780 10474
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14372 10260 14424 10266
rect 14648 10260 14700 10266
rect 14372 10202 14424 10208
rect 14568 10220 14648 10248
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14384 7886 14412 8298
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14476 6458 14504 7890
rect 14568 6882 14596 10220
rect 14648 10202 14700 10208
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14752 9110 14780 10202
rect 15108 9580 15160 9586
rect 15212 9568 15240 11494
rect 15304 11354 15332 11562
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15396 10713 15424 12718
rect 15382 10704 15438 10713
rect 15382 10639 15438 10648
rect 15160 9540 15240 9568
rect 15108 9522 15160 9528
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14660 7546 14688 8298
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15028 7546 15056 7958
rect 15488 7954 15516 16934
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15580 14074 15608 14554
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15580 13870 15608 14010
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15764 13530 15792 13942
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12986 15700 13330
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15580 12374 15608 12854
rect 15764 12442 15792 13126
rect 15856 12918 15884 13262
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15580 11150 15608 12310
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 16040 9450 16068 19654
rect 16316 19242 16344 22200
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16304 19236 16356 19242
rect 16304 19178 16356 19184
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16316 12646 16344 18566
rect 16592 16561 16620 19858
rect 16776 19174 16804 22200
rect 17236 20058 17264 22200
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16868 18834 16896 19246
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16578 16552 16634 16561
rect 16578 16487 16634 16496
rect 16592 12986 16620 16487
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16592 12782 16620 12922
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12102 16344 12582
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15580 8294 15608 8366
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14752 6882 14780 7414
rect 15580 7342 15608 8230
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14568 6866 14688 6882
rect 14568 6860 14700 6866
rect 14568 6854 14648 6860
rect 14752 6854 14872 6882
rect 14648 6802 14700 6808
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14568 6338 14596 6734
rect 14384 6310 14596 6338
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 13924 5630 14044 5658
rect 14384 5642 14412 6310
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 14372 5636 14424 5642
rect 13542 5264 13598 5273
rect 13542 5199 13598 5208
rect 13556 5030 13584 5199
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13740 4826 13768 5034
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13648 4282 13676 4626
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 4282 13860 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13924 4162 13952 5630
rect 14372 5578 14424 5584
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14016 5030 14044 5510
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13924 4134 14044 4162
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 3738 13676 4014
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13832 3534 13860 3878
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13832 3194 13860 3470
rect 13924 3466 13952 3946
rect 13912 3460 13964 3466
rect 13912 3402 13964 3408
rect 14016 3398 14044 4134
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12728 2582 12756 2790
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 13924 2514 13952 2858
rect 14108 2802 14136 5306
rect 14200 5273 14228 5306
rect 14186 5264 14242 5273
rect 14186 5199 14242 5208
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 3738 14228 4558
rect 14292 4010 14320 4626
rect 14384 4622 14412 5578
rect 14476 5030 14504 6190
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14568 5778 14596 6054
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14660 5574 14688 6190
rect 14752 5914 14780 6734
rect 14844 6458 14872 6854
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15212 6390 15240 6666
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14660 5234 14688 5510
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 15200 5092 15252 5098
rect 15200 5034 15252 5040
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4616 14424 4622
rect 14476 4604 14504 4966
rect 14568 4758 14596 4966
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15212 4826 15240 5034
rect 15304 4826 15332 6054
rect 15396 5817 15424 6054
rect 15382 5808 15438 5817
rect 15382 5743 15438 5752
rect 15488 5710 15516 7210
rect 15476 5704 15528 5710
rect 15382 5672 15438 5681
rect 15476 5646 15528 5652
rect 15382 5607 15438 5616
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14556 4616 14608 4622
rect 14476 4576 14556 4604
rect 14372 4558 14424 4564
rect 14556 4558 14608 4564
rect 14384 4282 14412 4558
rect 15016 4480 15068 4486
rect 15016 4422 15068 4428
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 15028 4146 15056 4422
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3398 14320 3538
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 15304 3126 15332 4422
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15396 2990 15424 5607
rect 15488 5234 15516 5646
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15568 3664 15620 3670
rect 15568 3606 15620 3612
rect 15580 2990 15608 3606
rect 15672 3602 15700 8230
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6322 15792 6598
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15752 5092 15804 5098
rect 15752 5034 15804 5040
rect 15764 4554 15792 5034
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 14384 2802 14412 2926
rect 14108 2774 14412 2802
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14108 2650 14136 2774
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 12636 2366 12848 2394
rect 12820 800 12848 2366
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 13280 800 13308 2246
rect 13740 800 13768 2246
rect 14292 800 14320 2246
rect 14752 800 14780 2790
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15212 800 15240 2790
rect 15396 2650 15424 2926
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15672 800 15700 2790
rect 15856 2650 15884 7890
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15948 6390 15976 7822
rect 16132 7818 16160 8230
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15936 6384 15988 6390
rect 15936 6326 15988 6332
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16040 5710 16068 6190
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 16316 3641 16344 12038
rect 17236 11286 17264 19178
rect 17512 18766 17540 19246
rect 17696 19174 17724 22200
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17512 11218 17540 18702
rect 18064 18630 18092 19246
rect 18156 19174 18184 22200
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18432 18902 18460 19246
rect 18616 19174 18644 22200
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18800 19310 18828 19654
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 5234 16712 7142
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16684 5098 16712 5170
rect 16672 5092 16724 5098
rect 16672 5034 16724 5040
rect 16302 3632 16358 3641
rect 16302 3567 16358 3576
rect 16396 3528 16448 3534
rect 16118 3496 16174 3505
rect 16396 3470 16448 3476
rect 16118 3431 16174 3440
rect 16132 3058 16160 3431
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16408 2990 16436 3470
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16040 2650 16068 2926
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15764 2106 15792 2246
rect 15752 2100 15804 2106
rect 15752 2042 15804 2048
rect 16132 800 16160 2790
rect 16592 800 16620 3062
rect 16776 2990 16804 7958
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 17052 5370 17080 5578
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16960 4826 16988 4966
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17052 4622 17080 5306
rect 17236 5030 17264 8570
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17420 5914 17448 6122
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17144 4078 17172 4422
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17236 2990 17264 4966
rect 17420 4604 17448 5850
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17512 4826 17540 5510
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17500 4616 17552 4622
rect 17420 4576 17500 4604
rect 17500 4558 17552 4564
rect 17604 2990 17632 6802
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17696 5914 17724 6394
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17788 5370 17816 18362
rect 17958 17232 18014 17241
rect 17958 17167 18014 17176
rect 17972 17066 18000 17167
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 18064 13802 18092 18566
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18800 14890 18828 19246
rect 19076 19174 19104 22200
rect 19536 20262 19564 22200
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 19168 19310 19196 19654
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19168 18358 19196 19246
rect 19536 18902 19564 19246
rect 19996 19242 20024 22200
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 20456 19174 20484 22200
rect 20916 19786 20944 22200
rect 21376 19990 21404 22200
rect 21836 20330 21864 22200
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21364 19984 21416 19990
rect 21364 19926 21416 19932
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 19524 18896 19576 18902
rect 19524 18838 19576 18844
rect 22296 18766 22324 22200
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 22756 14618 22784 22200
rect 22744 14612 22796 14618
rect 22744 14554 22796 14560
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18616 5817 18644 13126
rect 18602 5808 18658 5817
rect 18602 5743 18658 5752
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17788 5098 17816 5306
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17788 2990 17816 5034
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 18064 3602 18092 3946
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18156 3126 18184 5238
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19996 4690 20024 5034
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 20812 4480 20864 4486
rect 20812 4422 20864 4428
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 16776 2650 16804 2926
rect 17040 2916 17092 2922
rect 17040 2858 17092 2864
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17052 800 17080 2858
rect 17236 2650 17264 2926
rect 17328 2650 17356 2926
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17512 800 17540 2790
rect 17972 800 18000 3062
rect 18156 2990 18184 3062
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18064 2650 18092 2926
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18156 1442 18184 2790
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1414 18460 1442
rect 18432 800 18460 1414
rect 18984 800 19012 3334
rect 19432 3120 19484 3126
rect 19062 3088 19118 3097
rect 19432 3062 19484 3068
rect 19062 3023 19118 3032
rect 19076 2990 19104 3023
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19076 2650 19104 2926
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19444 800 19472 3062
rect 20180 3058 20208 3402
rect 20352 3120 20404 3126
rect 20352 3062 20404 3068
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 19904 800 19932 2858
rect 20364 800 20392 3062
rect 20824 800 20852 4422
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21284 800 21312 2790
rect 21732 2100 21784 2106
rect 21732 2042 21784 2048
rect 21744 800 21772 2042
rect 22204 800 22232 3130
rect 22664 800 22692 4082
rect 6366 640 6422 649
rect 6366 575 6422 584
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20350 0 20406 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21730 0 21786 800
rect 22190 0 22246 800
rect 22650 0 22706 800
<< via2 >>
rect 3054 22616 3110 22672
rect 1582 21120 1638 21176
rect 1674 20712 1730 20768
rect 1582 19760 1638 19816
rect 1582 18808 1638 18864
rect 1766 18828 1822 18864
rect 1766 18808 1768 18828
rect 1768 18808 1820 18828
rect 1820 18808 1822 18828
rect 1950 20168 2006 20224
rect 1950 19216 2006 19272
rect 2870 22072 2926 22128
rect 2778 21664 2834 21720
rect 2042 18672 2098 18728
rect 2686 19216 2742 19272
rect 1950 18300 1952 18320
rect 1952 18300 2004 18320
rect 2004 18300 2006 18320
rect 1950 18264 2006 18300
rect 2962 18944 3018 19000
rect 1674 17856 1730 17912
rect 1582 17312 1638 17368
rect 1858 18128 1914 18184
rect 202 16632 258 16688
rect 2502 17040 2558 17096
rect 1950 16904 2006 16960
rect 1950 16360 2006 16416
rect 2778 15952 2834 16008
rect 1950 15000 2006 15056
rect 2778 15408 2834 15464
rect 1858 14456 1914 14512
rect 1766 13524 1822 13560
rect 1766 13504 1768 13524
rect 1768 13504 1820 13524
rect 1820 13504 1822 13524
rect 2778 14068 2834 14104
rect 2778 14048 2780 14068
rect 2780 14048 2832 14068
rect 2832 14048 2834 14068
rect 2778 4120 2834 4176
rect 1490 2080 1546 2136
rect 1582 1128 1638 1184
rect 2870 3032 2926 3088
rect 3882 13776 3938 13832
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4618 19080 4674 19136
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4802 18128 4858 18184
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 3882 12552 3938 12608
rect 3882 12144 3938 12200
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4066 11600 4122 11656
rect 3974 11056 4030 11112
rect 3974 10648 4030 10704
rect 3974 10124 4030 10160
rect 3974 10104 3976 10124
rect 3976 10104 4028 10124
rect 4028 10104 4030 10124
rect 4066 9716 4122 9752
rect 4066 9696 4068 9716
rect 4068 9696 4120 9716
rect 4120 9696 4122 9716
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4066 9152 4122 9208
rect 4066 7792 4122 7848
rect 4066 7248 4122 7304
rect 3514 5344 3570 5400
rect 3514 4800 3570 4856
rect 3698 3984 3754 4040
rect 3238 3440 3294 3496
rect 3698 2796 3700 2816
rect 3700 2796 3752 2816
rect 3752 2796 3754 2816
rect 3698 2760 3754 2796
rect 4066 6296 4122 6352
rect 4066 5888 4122 5944
rect 3974 4936 4030 4992
rect 4066 4392 4122 4448
rect 4066 3440 4122 3496
rect 4434 9968 4490 10024
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 5078 19080 5134 19136
rect 5722 19080 5778 19136
rect 4894 9968 4950 10024
rect 6274 19216 6330 19272
rect 5998 18944 6054 19000
rect 5262 8200 5318 8256
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 5262 7148 5264 7168
rect 5264 7148 5316 7168
rect 5316 7148 5318 7168
rect 5262 7112 5318 7148
rect 5078 3984 5134 4040
rect 4066 2508 4122 2544
rect 4066 2488 4068 2508
rect 4068 2488 4120 2508
rect 4120 2488 4122 2508
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5814 8744 5870 8800
rect 5630 3984 5686 4040
rect 5170 1536 5226 1592
rect 6274 10104 6330 10160
rect 6182 8744 6238 8800
rect 5906 6724 5962 6760
rect 5906 6704 5908 6724
rect 5908 6704 5960 6724
rect 5960 6704 5962 6724
rect 7286 17040 7342 17096
rect 6090 3984 6146 4040
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7470 12416 7526 12472
rect 7470 12280 7526 12336
rect 7102 8880 7158 8936
rect 6274 2760 6330 2816
rect 3054 176 3110 232
rect 6734 4800 6790 4856
rect 7010 4120 7066 4176
rect 8298 13912 8354 13968
rect 7838 13812 7840 13832
rect 7840 13812 7892 13832
rect 7892 13812 7894 13832
rect 7838 13776 7894 13812
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 8298 13776 8354 13832
rect 8482 16632 8538 16688
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7838 9968 7894 10024
rect 7838 9424 7894 9480
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8206 9016 8262 9072
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7378 6704 7434 6760
rect 7470 6160 7526 6216
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 8482 10512 8538 10568
rect 8666 10376 8722 10432
rect 8482 8608 8538 8664
rect 10414 18808 10470 18864
rect 10322 18672 10378 18728
rect 8850 10376 8906 10432
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7746 5616 7802 5672
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 8574 6860 8630 6896
rect 8574 6840 8576 6860
rect 8576 6840 8628 6860
rect 8628 6840 8630 6860
rect 8390 5652 8392 5672
rect 8392 5652 8444 5672
rect 8444 5652 8446 5672
rect 8390 5616 8446 5652
rect 8942 3596 8998 3632
rect 8942 3576 8944 3596
rect 8944 3576 8996 3596
rect 8996 3576 8998 3596
rect 9586 13232 9642 13288
rect 10598 16532 10600 16552
rect 10600 16532 10652 16552
rect 10652 16532 10654 16552
rect 10598 16496 10654 16532
rect 10322 14728 10378 14784
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10506 13912 10562 13968
rect 10230 12436 10286 12472
rect 10230 12416 10232 12436
rect 10232 12416 10284 12436
rect 10284 12416 10286 12436
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 10046 10512 10102 10568
rect 9494 9016 9550 9072
rect 9586 8744 9642 8800
rect 9494 8508 9496 8528
rect 9496 8508 9548 8528
rect 9548 8508 9550 8528
rect 9494 8472 9550 8508
rect 9862 8608 9918 8664
rect 9770 5888 9826 5944
rect 9678 5788 9680 5808
rect 9680 5788 9732 5808
rect 9732 5788 9734 5808
rect 9678 5752 9734 5788
rect 10598 10104 10654 10160
rect 10598 8608 10654 8664
rect 10046 4120 10102 4176
rect 10138 3612 10140 3632
rect 10140 3612 10192 3632
rect 10192 3612 10194 3632
rect 9770 3440 9826 3496
rect 9770 3168 9826 3224
rect 9678 3032 9734 3088
rect 10138 3576 10194 3612
rect 10046 3304 10102 3360
rect 10322 3304 10378 3360
rect 10874 8744 10930 8800
rect 11610 13388 11666 13424
rect 11610 13368 11612 13388
rect 11612 13368 11664 13388
rect 11664 13368 11666 13388
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11610 12280 11666 12336
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11978 14356 11980 14376
rect 11980 14356 12032 14376
rect 12032 14356 12034 14376
rect 11978 14320 12034 14356
rect 11886 12416 11942 12472
rect 12622 14456 12678 14512
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11702 10648 11758 10704
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11242 8880 11298 8936
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 10966 5908 11022 5944
rect 10966 5888 10968 5908
rect 10968 5888 11020 5908
rect 11020 5888 11022 5908
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 12070 10240 12126 10296
rect 11978 6704 12034 6760
rect 11058 3168 11114 3224
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11426 3440 11482 3496
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 10506 856 10562 912
rect 12714 12280 12770 12336
rect 13450 14492 13452 14512
rect 13452 14492 13504 14512
rect 13504 14492 13506 14512
rect 13450 14456 13506 14492
rect 13634 14320 13690 14376
rect 13450 13932 13506 13968
rect 13450 13912 13452 13932
rect 13452 13912 13504 13932
rect 13504 13912 13506 13932
rect 13266 13368 13322 13424
rect 13082 9560 13138 9616
rect 13450 10104 13506 10160
rect 13358 9424 13414 9480
rect 12622 6160 12678 6216
rect 12254 4156 12256 4176
rect 12256 4156 12308 4176
rect 12308 4156 12310 4176
rect 12254 4120 12310 4156
rect 12254 3984 12310 4040
rect 14186 19352 14242 19408
rect 14554 19488 14610 19544
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14554 14728 14610 14784
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 15382 14456 15438 14512
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15382 10648 15438 10704
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 16578 16496 16634 16552
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 13542 5208 13598 5264
rect 14186 5208 14242 5264
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 15382 5752 15438 5808
rect 15382 5616 15438 5672
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 16302 3576 16358 3632
rect 16118 3440 16174 3496
rect 17958 17176 18014 17232
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18602 5752 18658 5808
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19062 3032 19118 3088
rect 6366 584 6422 640
<< metal3 >>
rect 0 22674 800 22704
rect 3049 22674 3115 22677
rect 0 22672 3115 22674
rect 0 22616 3054 22672
rect 3110 22616 3115 22672
rect 0 22614 3115 22616
rect 0 22584 800 22614
rect 3049 22611 3115 22614
rect 0 22130 800 22160
rect 2865 22130 2931 22133
rect 0 22128 2931 22130
rect 0 22072 2870 22128
rect 2926 22072 2931 22128
rect 0 22070 2931 22072
rect 0 22040 800 22070
rect 2865 22067 2931 22070
rect 0 21722 800 21752
rect 2773 21722 2839 21725
rect 0 21720 2839 21722
rect 0 21664 2778 21720
rect 2834 21664 2839 21720
rect 0 21662 2839 21664
rect 0 21632 800 21662
rect 2773 21659 2839 21662
rect 0 21178 800 21208
rect 1577 21178 1643 21181
rect 0 21176 1643 21178
rect 0 21120 1582 21176
rect 1638 21120 1643 21176
rect 0 21118 1643 21120
rect 0 21088 800 21118
rect 1577 21115 1643 21118
rect 0 20770 800 20800
rect 1669 20770 1735 20773
rect 0 20768 1735 20770
rect 0 20712 1674 20768
rect 1730 20712 1735 20768
rect 0 20710 1735 20712
rect 0 20680 800 20710
rect 1669 20707 1735 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20226 800 20256
rect 1945 20226 2011 20229
rect 0 20224 2011 20226
rect 0 20168 1950 20224
rect 2006 20168 2011 20224
rect 0 20166 2011 20168
rect 0 20136 800 20166
rect 1945 20163 2011 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 0 19818 800 19848
rect 1577 19818 1643 19821
rect 0 19816 1643 19818
rect 0 19760 1582 19816
rect 1638 19760 1643 19816
rect 0 19758 1643 19760
rect 0 19728 800 19758
rect 1577 19755 1643 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 14549 19546 14615 19549
rect 14046 19544 14615 19546
rect 14046 19488 14554 19544
rect 14610 19488 14615 19544
rect 14046 19486 14615 19488
rect 14046 19410 14106 19486
rect 14549 19483 14615 19486
rect 14181 19410 14247 19413
rect 14046 19408 14247 19410
rect 14046 19352 14186 19408
rect 14242 19352 14247 19408
rect 14046 19350 14247 19352
rect 14181 19347 14247 19350
rect 0 19274 800 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 800 19214
rect 1945 19211 2011 19214
rect 2681 19274 2747 19277
rect 6269 19274 6335 19277
rect 2681 19272 6335 19274
rect 2681 19216 2686 19272
rect 2742 19216 6274 19272
rect 6330 19216 6335 19272
rect 2681 19214 6335 19216
rect 2681 19211 2747 19214
rect 6269 19211 6335 19214
rect 4613 19138 4679 19141
rect 5073 19138 5139 19141
rect 5717 19140 5783 19141
rect 5717 19138 5764 19140
rect 4613 19136 5139 19138
rect 4613 19080 4618 19136
rect 4674 19080 5078 19136
rect 5134 19080 5139 19136
rect 4613 19078 5139 19080
rect 5672 19136 5764 19138
rect 5672 19080 5722 19136
rect 5672 19078 5764 19080
rect 4613 19075 4679 19078
rect 5073 19075 5139 19078
rect 5717 19076 5764 19078
rect 5828 19076 5834 19140
rect 5717 19075 5783 19076
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 2957 19002 3023 19005
rect 5993 19002 6059 19005
rect 2957 19000 6059 19002
rect 2957 18944 2962 19000
rect 3018 18944 5998 19000
rect 6054 18944 6059 19000
rect 2957 18942 6059 18944
rect 2957 18939 3023 18942
rect 5993 18939 6059 18942
rect 0 18866 800 18896
rect 1577 18866 1643 18869
rect 0 18864 1643 18866
rect 0 18808 1582 18864
rect 1638 18808 1643 18864
rect 0 18806 1643 18808
rect 0 18776 800 18806
rect 1577 18803 1643 18806
rect 1761 18866 1827 18869
rect 10409 18866 10475 18869
rect 1761 18864 10475 18866
rect 1761 18808 1766 18864
rect 1822 18808 10414 18864
rect 10470 18808 10475 18864
rect 1761 18806 10475 18808
rect 1761 18803 1827 18806
rect 10409 18803 10475 18806
rect 2037 18730 2103 18733
rect 10317 18730 10383 18733
rect 2037 18728 10383 18730
rect 2037 18672 2042 18728
rect 2098 18672 10322 18728
rect 10378 18672 10383 18728
rect 2037 18670 10383 18672
rect 2037 18667 2103 18670
rect 10317 18667 10383 18670
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 0 18322 800 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 800 18262
rect 1945 18259 2011 18262
rect 1853 18186 1919 18189
rect 4797 18186 4863 18189
rect 1853 18184 4863 18186
rect 1853 18128 1858 18184
rect 1914 18128 4802 18184
rect 4858 18128 4863 18184
rect 1853 18126 4863 18128
rect 1853 18123 1919 18126
rect 4797 18123 4863 18126
rect 7874 17984 8194 17985
rect 0 17914 800 17944
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 1669 17914 1735 17917
rect 0 17912 1735 17914
rect 0 17856 1674 17912
rect 1730 17856 1735 17912
rect 0 17854 1735 17856
rect 0 17824 800 17854
rect 1669 17851 1735 17854
rect 4409 17440 4729 17441
rect 0 17370 800 17400
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 800 17310
rect 1577 17307 1643 17310
rect 17953 17234 18019 17237
rect 22200 17234 23000 17264
rect 17953 17232 23000 17234
rect 17953 17176 17958 17232
rect 18014 17176 23000 17232
rect 17953 17174 23000 17176
rect 17953 17171 18019 17174
rect 22200 17144 23000 17174
rect 2497 17098 2563 17101
rect 7281 17098 7347 17101
rect 2497 17096 7347 17098
rect 2497 17040 2502 17096
rect 2558 17040 7286 17096
rect 7342 17040 7347 17096
rect 2497 17038 7347 17040
rect 2497 17035 2563 17038
rect 7281 17035 7347 17038
rect 0 16962 800 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 800 16902
rect 1945 16899 2011 16902
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 197 16690 263 16693
rect 8477 16690 8543 16693
rect 197 16688 8543 16690
rect 197 16632 202 16688
rect 258 16632 8482 16688
rect 8538 16632 8543 16688
rect 197 16630 8543 16632
rect 197 16627 263 16630
rect 8477 16627 8543 16630
rect 10593 16554 10659 16557
rect 16573 16554 16639 16557
rect 10593 16552 16639 16554
rect 10593 16496 10598 16552
rect 10654 16496 16578 16552
rect 16634 16496 16639 16552
rect 10593 16494 16639 16496
rect 10593 16491 10659 16494
rect 16573 16491 16639 16494
rect 0 16418 800 16448
rect 1945 16418 2011 16421
rect 0 16416 2011 16418
rect 0 16360 1950 16416
rect 2006 16360 2011 16416
rect 0 16358 2011 16360
rect 0 16328 800 16358
rect 1945 16355 2011 16358
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16010 800 16040
rect 2773 16010 2839 16013
rect 0 16008 2839 16010
rect 0 15952 2778 16008
rect 2834 15952 2839 16008
rect 0 15950 2839 15952
rect 0 15920 800 15950
rect 2773 15947 2839 15950
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15466 800 15496
rect 2773 15466 2839 15469
rect 0 15464 2839 15466
rect 0 15408 2778 15464
rect 2834 15408 2839 15464
rect 0 15406 2839 15408
rect 0 15376 800 15406
rect 2773 15403 2839 15406
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 0 15058 800 15088
rect 1945 15058 2011 15061
rect 0 15056 2011 15058
rect 0 15000 1950 15056
rect 2006 15000 2011 15056
rect 0 14998 2011 15000
rect 0 14968 800 14998
rect 1945 14995 2011 14998
rect 10317 14786 10383 14789
rect 14549 14786 14615 14789
rect 10317 14784 14615 14786
rect 10317 14728 10322 14784
rect 10378 14728 14554 14784
rect 14610 14728 14615 14784
rect 10317 14726 14615 14728
rect 10317 14723 10383 14726
rect 14549 14723 14615 14726
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 0 14514 800 14544
rect 1853 14514 1919 14517
rect 0 14512 1919 14514
rect 0 14456 1858 14512
rect 1914 14456 1919 14512
rect 0 14454 1919 14456
rect 0 14424 800 14454
rect 1853 14451 1919 14454
rect 12617 14514 12683 14517
rect 13445 14514 13511 14517
rect 15377 14514 15443 14517
rect 12617 14512 15443 14514
rect 12617 14456 12622 14512
rect 12678 14456 13450 14512
rect 13506 14456 15382 14512
rect 15438 14456 15443 14512
rect 12617 14454 15443 14456
rect 12617 14451 12683 14454
rect 13445 14451 13511 14454
rect 15377 14451 15443 14454
rect 11973 14378 12039 14381
rect 13629 14378 13695 14381
rect 11973 14376 13695 14378
rect 11973 14320 11978 14376
rect 12034 14320 13634 14376
rect 13690 14320 13695 14376
rect 11973 14318 13695 14320
rect 11973 14315 12039 14318
rect 13629 14315 13695 14318
rect 4409 14176 4729 14177
rect 0 14106 800 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 2773 14106 2839 14109
rect 0 14104 2839 14106
rect 0 14048 2778 14104
rect 2834 14048 2839 14104
rect 0 14046 2839 14048
rect 0 14016 800 14046
rect 2773 14043 2839 14046
rect 8293 13970 8359 13973
rect 3880 13968 8359 13970
rect 3880 13912 8298 13968
rect 8354 13912 8359 13968
rect 3880 13910 8359 13912
rect 3880 13837 3940 13910
rect 8293 13907 8359 13910
rect 10501 13970 10567 13973
rect 13445 13970 13511 13973
rect 10501 13968 13511 13970
rect 10501 13912 10506 13968
rect 10562 13912 13450 13968
rect 13506 13912 13511 13968
rect 10501 13910 13511 13912
rect 10501 13907 10567 13910
rect 13445 13907 13511 13910
rect 3877 13832 3943 13837
rect 3877 13776 3882 13832
rect 3938 13776 3943 13832
rect 3877 13771 3943 13776
rect 7833 13834 7899 13837
rect 8293 13834 8359 13837
rect 7833 13832 8359 13834
rect 7833 13776 7838 13832
rect 7894 13776 8298 13832
rect 8354 13776 8359 13832
rect 7833 13774 8359 13776
rect 7833 13771 7899 13774
rect 8293 13771 8359 13774
rect 7874 13632 8194 13633
rect 0 13562 800 13592
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 1761 13562 1827 13565
rect 0 13560 1827 13562
rect 0 13504 1766 13560
rect 1822 13504 1827 13560
rect 0 13502 1827 13504
rect 0 13472 800 13502
rect 1761 13499 1827 13502
rect 11605 13426 11671 13429
rect 13261 13426 13327 13429
rect 11605 13424 13327 13426
rect 11605 13368 11610 13424
rect 11666 13368 13266 13424
rect 13322 13368 13327 13424
rect 11605 13366 13327 13368
rect 11605 13363 11671 13366
rect 13261 13363 13327 13366
rect 9581 13290 9647 13293
rect 4110 13288 9647 13290
rect 4110 13232 9586 13288
rect 9642 13232 9647 13288
rect 4110 13230 9647 13232
rect 0 13154 800 13184
rect 4110 13154 4170 13230
rect 9581 13227 9647 13230
rect 0 13094 4170 13154
rect 0 13064 800 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12610 800 12640
rect 3877 12610 3943 12613
rect 0 12608 3943 12610
rect 0 12552 3882 12608
rect 3938 12552 3943 12608
rect 0 12550 3943 12552
rect 0 12520 800 12550
rect 3877 12547 3943 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 7465 12476 7531 12477
rect 7414 12474 7420 12476
rect 7374 12414 7420 12474
rect 7484 12472 7531 12476
rect 7526 12416 7531 12472
rect 7414 12412 7420 12414
rect 7484 12412 7531 12416
rect 7465 12411 7531 12412
rect 10225 12474 10291 12477
rect 11881 12474 11947 12477
rect 10225 12472 11947 12474
rect 10225 12416 10230 12472
rect 10286 12416 11886 12472
rect 11942 12416 11947 12472
rect 10225 12414 11947 12416
rect 10225 12411 10291 12414
rect 11881 12411 11947 12414
rect 7465 12340 7531 12341
rect 7414 12276 7420 12340
rect 7484 12338 7531 12340
rect 11605 12338 11671 12341
rect 12709 12338 12775 12341
rect 7484 12336 7576 12338
rect 7526 12280 7576 12336
rect 7484 12278 7576 12280
rect 11605 12336 12775 12338
rect 11605 12280 11610 12336
rect 11666 12280 12714 12336
rect 12770 12280 12775 12336
rect 11605 12278 12775 12280
rect 7484 12276 7531 12278
rect 7465 12275 7531 12276
rect 11605 12275 11671 12278
rect 12709 12275 12775 12278
rect 0 12202 800 12232
rect 3877 12202 3943 12205
rect 0 12200 3943 12202
rect 0 12144 3882 12200
rect 3938 12144 3943 12200
rect 0 12142 3943 12144
rect 0 12112 800 12142
rect 3877 12139 3943 12142
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 0 11658 800 11688
rect 4061 11658 4127 11661
rect 0 11656 4127 11658
rect 0 11600 4066 11656
rect 4122 11600 4127 11656
rect 0 11598 4127 11600
rect 0 11568 800 11598
rect 4061 11595 4127 11598
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 0 11114 800 11144
rect 3969 11114 4035 11117
rect 0 11112 4035 11114
rect 0 11056 3974 11112
rect 4030 11056 4035 11112
rect 0 11054 4035 11056
rect 0 11024 800 11054
rect 3969 11051 4035 11054
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 0 10706 800 10736
rect 3969 10706 4035 10709
rect 0 10704 4035 10706
rect 0 10648 3974 10704
rect 4030 10648 4035 10704
rect 0 10646 4035 10648
rect 0 10616 800 10646
rect 3969 10643 4035 10646
rect 11697 10706 11763 10709
rect 15377 10706 15443 10709
rect 11697 10704 15443 10706
rect 11697 10648 11702 10704
rect 11758 10648 15382 10704
rect 15438 10648 15443 10704
rect 11697 10646 15443 10648
rect 11697 10643 11763 10646
rect 15377 10643 15443 10646
rect 8477 10570 8543 10573
rect 10041 10570 10107 10573
rect 8477 10568 10107 10570
rect 8477 10512 8482 10568
rect 8538 10512 10046 10568
rect 10102 10512 10107 10568
rect 8477 10510 10107 10512
rect 8477 10507 8543 10510
rect 10041 10507 10107 10510
rect 8661 10434 8727 10437
rect 8845 10434 8911 10437
rect 8661 10432 8911 10434
rect 8661 10376 8666 10432
rect 8722 10376 8850 10432
rect 8906 10376 8911 10432
rect 8661 10374 8911 10376
rect 8661 10371 8727 10374
rect 8845 10371 8911 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 12065 10298 12131 10301
rect 8526 10296 12131 10298
rect 8526 10240 12070 10296
rect 12126 10240 12131 10296
rect 8526 10238 12131 10240
rect 0 10162 800 10192
rect 3969 10162 4035 10165
rect 0 10160 4035 10162
rect 0 10104 3974 10160
rect 4030 10104 4035 10160
rect 0 10102 4035 10104
rect 0 10072 800 10102
rect 3969 10099 4035 10102
rect 6269 10162 6335 10165
rect 8526 10162 8586 10238
rect 12065 10235 12131 10238
rect 6269 10160 8586 10162
rect 6269 10104 6274 10160
rect 6330 10104 8586 10160
rect 6269 10102 8586 10104
rect 10593 10162 10659 10165
rect 13445 10162 13511 10165
rect 10593 10160 13511 10162
rect 10593 10104 10598 10160
rect 10654 10104 13450 10160
rect 13506 10104 13511 10160
rect 10593 10102 13511 10104
rect 6269 10099 6335 10102
rect 10593 10099 10659 10102
rect 13445 10099 13511 10102
rect 4429 10026 4495 10029
rect 4889 10026 4955 10029
rect 4429 10024 4955 10026
rect 4429 9968 4434 10024
rect 4490 9968 4894 10024
rect 4950 9968 4955 10024
rect 4429 9966 4955 9968
rect 4429 9963 4495 9966
rect 4889 9963 4955 9966
rect 5758 9964 5764 10028
rect 5828 10026 5834 10028
rect 7833 10026 7899 10029
rect 5828 10024 7899 10026
rect 5828 9968 7838 10024
rect 7894 9968 7899 10024
rect 5828 9966 7899 9968
rect 5828 9964 5834 9966
rect 7833 9963 7899 9966
rect 4409 9824 4729 9825
rect 0 9754 800 9784
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 4061 9754 4127 9757
rect 0 9752 4127 9754
rect 0 9696 4066 9752
rect 4122 9696 4127 9752
rect 0 9694 4127 9696
rect 0 9664 800 9694
rect 4061 9691 4127 9694
rect 13077 9618 13143 9621
rect 13077 9616 13186 9618
rect 13077 9560 13082 9616
rect 13138 9560 13186 9616
rect 13077 9555 13186 9560
rect 7598 9420 7604 9484
rect 7668 9482 7674 9484
rect 7833 9482 7899 9485
rect 7668 9480 7899 9482
rect 7668 9424 7838 9480
rect 7894 9424 7899 9480
rect 7668 9422 7899 9424
rect 13126 9482 13186 9555
rect 13353 9482 13419 9485
rect 13126 9480 13419 9482
rect 13126 9424 13358 9480
rect 13414 9424 13419 9480
rect 13126 9422 13419 9424
rect 7668 9420 7674 9422
rect 7833 9419 7899 9422
rect 13353 9419 13419 9422
rect 7874 9280 8194 9281
rect 0 9210 800 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 4061 9210 4127 9213
rect 0 9208 4127 9210
rect 0 9152 4066 9208
rect 4122 9152 4127 9208
rect 0 9150 4127 9152
rect 0 9120 800 9150
rect 4061 9147 4127 9150
rect 8201 9074 8267 9077
rect 9489 9074 9555 9077
rect 8201 9072 9555 9074
rect 8201 9016 8206 9072
rect 8262 9016 9494 9072
rect 9550 9016 9555 9072
rect 8201 9014 9555 9016
rect 8201 9011 8267 9014
rect 9489 9011 9555 9014
rect 7097 8938 7163 8941
rect 11237 8938 11303 8941
rect 7097 8936 11303 8938
rect 7097 8880 7102 8936
rect 7158 8880 11242 8936
rect 11298 8880 11303 8936
rect 7097 8878 11303 8880
rect 7097 8875 7163 8878
rect 11237 8875 11303 8878
rect 0 8802 800 8832
rect 5809 8802 5875 8805
rect 6177 8802 6243 8805
rect 0 8742 4170 8802
rect 0 8712 800 8742
rect 4110 8530 4170 8742
rect 5809 8800 6243 8802
rect 5809 8744 5814 8800
rect 5870 8744 6182 8800
rect 6238 8744 6243 8800
rect 5809 8742 6243 8744
rect 5809 8739 5875 8742
rect 6177 8739 6243 8742
rect 9581 8802 9647 8805
rect 10869 8802 10935 8805
rect 9581 8800 10935 8802
rect 9581 8744 9586 8800
rect 9642 8744 10874 8800
rect 10930 8744 10935 8800
rect 9581 8742 10935 8744
rect 9581 8739 9647 8742
rect 10869 8739 10935 8742
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 8477 8666 8543 8669
rect 9857 8666 9923 8669
rect 10593 8668 10659 8669
rect 10542 8666 10548 8668
rect 8477 8664 9923 8666
rect 8477 8608 8482 8664
rect 8538 8608 9862 8664
rect 9918 8608 9923 8664
rect 8477 8606 9923 8608
rect 10502 8606 10548 8666
rect 10612 8664 10659 8668
rect 10654 8608 10659 8664
rect 8477 8603 8543 8606
rect 9857 8603 9923 8606
rect 10542 8604 10548 8606
rect 10612 8604 10659 8608
rect 10593 8603 10659 8604
rect 9489 8530 9555 8533
rect 4110 8528 9555 8530
rect 4110 8472 9494 8528
rect 9550 8472 9555 8528
rect 4110 8470 9555 8472
rect 9489 8467 9555 8470
rect 0 8258 800 8288
rect 5257 8258 5323 8261
rect 0 8256 5323 8258
rect 0 8200 5262 8256
rect 5318 8200 5323 8256
rect 0 8198 5323 8200
rect 0 8168 800 8198
rect 5257 8195 5323 8198
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 0 7850 800 7880
rect 4061 7850 4127 7853
rect 0 7848 4127 7850
rect 0 7792 4066 7848
rect 4122 7792 4127 7848
rect 0 7790 4127 7792
rect 0 7760 800 7790
rect 4061 7787 4127 7790
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 0 7306 800 7336
rect 4061 7306 4127 7309
rect 0 7304 4127 7306
rect 0 7248 4066 7304
rect 4122 7248 4127 7304
rect 0 7246 4127 7248
rect 0 7216 800 7246
rect 4061 7243 4127 7246
rect 5257 7170 5323 7173
rect 7598 7170 7604 7172
rect 5257 7168 7604 7170
rect 5257 7112 5262 7168
rect 5318 7112 7604 7168
rect 5257 7110 7604 7112
rect 5257 7107 5323 7110
rect 7598 7108 7604 7110
rect 7668 7108 7674 7172
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6898 800 6928
rect 8569 6898 8635 6901
rect 0 6896 8635 6898
rect 0 6840 8574 6896
rect 8630 6840 8635 6896
rect 0 6838 8635 6840
rect 0 6808 800 6838
rect 8569 6835 8635 6838
rect 5901 6762 5967 6765
rect 7373 6762 7439 6765
rect 11973 6762 12039 6765
rect 5901 6760 12039 6762
rect 5901 6704 5906 6760
rect 5962 6704 7378 6760
rect 7434 6704 11978 6760
rect 12034 6704 12039 6760
rect 5901 6702 12039 6704
rect 5901 6699 5967 6702
rect 7373 6699 7439 6702
rect 11973 6699 12039 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6354 800 6384
rect 4061 6354 4127 6357
rect 0 6352 4127 6354
rect 0 6296 4066 6352
rect 4122 6296 4127 6352
rect 0 6294 4127 6296
rect 0 6264 800 6294
rect 4061 6291 4127 6294
rect 7465 6218 7531 6221
rect 12617 6218 12683 6221
rect 7465 6216 12683 6218
rect 7465 6160 7470 6216
rect 7526 6160 12622 6216
rect 12678 6160 12683 6216
rect 7465 6158 12683 6160
rect 7465 6155 7531 6158
rect 12617 6155 12683 6158
rect 7874 6016 8194 6017
rect 0 5946 800 5976
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 4061 5946 4127 5949
rect 0 5944 4127 5946
rect 0 5888 4066 5944
rect 4122 5888 4127 5944
rect 0 5886 4127 5888
rect 0 5856 800 5886
rect 4061 5883 4127 5886
rect 9765 5946 9831 5949
rect 10961 5946 11027 5949
rect 9765 5944 11027 5946
rect 9765 5888 9770 5944
rect 9826 5888 10966 5944
rect 11022 5888 11027 5944
rect 9765 5886 11027 5888
rect 9765 5883 9831 5886
rect 10961 5883 11027 5886
rect 9673 5810 9739 5813
rect 15377 5810 15443 5813
rect 9673 5808 15443 5810
rect 9673 5752 9678 5808
rect 9734 5752 15382 5808
rect 15438 5752 15443 5808
rect 9673 5750 15443 5752
rect 9673 5747 9739 5750
rect 15377 5747 15443 5750
rect 18597 5810 18663 5813
rect 22200 5810 23000 5840
rect 18597 5808 23000 5810
rect 18597 5752 18602 5808
rect 18658 5752 23000 5808
rect 18597 5750 23000 5752
rect 18597 5747 18663 5750
rect 22200 5720 23000 5750
rect 7598 5612 7604 5676
rect 7668 5674 7674 5676
rect 7741 5674 7807 5677
rect 8385 5674 8451 5677
rect 15377 5674 15443 5677
rect 7668 5672 15443 5674
rect 7668 5616 7746 5672
rect 7802 5616 8390 5672
rect 8446 5616 15382 5672
rect 15438 5616 15443 5672
rect 7668 5614 15443 5616
rect 7668 5612 7674 5614
rect 7741 5611 7807 5614
rect 8385 5611 8451 5614
rect 15377 5611 15443 5614
rect 4409 5472 4729 5473
rect 0 5402 800 5432
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 3509 5402 3575 5405
rect 0 5400 3575 5402
rect 0 5344 3514 5400
rect 3570 5344 3575 5400
rect 0 5342 3575 5344
rect 0 5312 800 5342
rect 3509 5339 3575 5342
rect 13537 5266 13603 5269
rect 14181 5266 14247 5269
rect 13537 5264 14247 5266
rect 13537 5208 13542 5264
rect 13598 5208 14186 5264
rect 14242 5208 14247 5264
rect 13537 5206 14247 5208
rect 13537 5203 13603 5206
rect 14181 5203 14247 5206
rect 0 4994 800 5024
rect 3969 4994 4035 4997
rect 0 4992 4035 4994
rect 0 4936 3974 4992
rect 4030 4936 4035 4992
rect 0 4934 4035 4936
rect 0 4904 800 4934
rect 3969 4931 4035 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 3509 4858 3575 4861
rect 6729 4858 6795 4861
rect 3509 4856 6795 4858
rect 3509 4800 3514 4856
rect 3570 4800 6734 4856
rect 6790 4800 6795 4856
rect 3509 4798 6795 4800
rect 3509 4795 3575 4798
rect 6729 4795 6795 4798
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 2773 4178 2839 4181
rect 7005 4178 7071 4181
rect 2773 4176 7071 4178
rect 2773 4120 2778 4176
rect 2834 4120 7010 4176
rect 7066 4120 7071 4176
rect 2773 4118 7071 4120
rect 2773 4115 2839 4118
rect 7005 4115 7071 4118
rect 10041 4178 10107 4181
rect 12249 4178 12315 4181
rect 10041 4176 12315 4178
rect 10041 4120 10046 4176
rect 10102 4120 12254 4176
rect 12310 4120 12315 4176
rect 10041 4118 12315 4120
rect 10041 4115 10107 4118
rect 12249 4115 12315 4118
rect 0 4042 800 4072
rect 3693 4042 3759 4045
rect 0 4040 3759 4042
rect 0 3984 3698 4040
rect 3754 3984 3759 4040
rect 0 3982 3759 3984
rect 0 3952 800 3982
rect 3693 3979 3759 3982
rect 5073 4042 5139 4045
rect 5625 4042 5691 4045
rect 6085 4042 6151 4045
rect 12249 4042 12315 4045
rect 5073 4040 6010 4042
rect 5073 3984 5078 4040
rect 5134 3984 5630 4040
rect 5686 3984 6010 4040
rect 5073 3982 6010 3984
rect 5073 3979 5139 3982
rect 5625 3979 5691 3982
rect 5950 3770 6010 3982
rect 6085 4040 12315 4042
rect 6085 3984 6090 4040
rect 6146 3984 12254 4040
rect 12310 3984 12315 4040
rect 6085 3982 12315 3984
rect 6085 3979 6151 3982
rect 12249 3979 12315 3982
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 5950 3710 6746 3770
rect 6686 3634 6746 3710
rect 8937 3634 9003 3637
rect 6686 3632 9003 3634
rect 6686 3576 8942 3632
rect 8998 3576 9003 3632
rect 6686 3574 9003 3576
rect 8937 3571 9003 3574
rect 10133 3634 10199 3637
rect 16297 3634 16363 3637
rect 10133 3632 16363 3634
rect 10133 3576 10138 3632
rect 10194 3576 16302 3632
rect 16358 3576 16363 3632
rect 10133 3574 16363 3576
rect 10133 3571 10199 3574
rect 16297 3571 16363 3574
rect 0 3498 800 3528
rect 3233 3498 3299 3501
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 3238 3496
rect 3294 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3408 800 3438
rect 3233 3435 3299 3438
rect 4061 3435 4127 3438
rect 9765 3498 9831 3501
rect 11421 3498 11487 3501
rect 16113 3498 16179 3501
rect 9765 3496 16179 3498
rect 9765 3440 9770 3496
rect 9826 3440 11426 3496
rect 11482 3440 16118 3496
rect 16174 3440 16179 3496
rect 9765 3438 16179 3440
rect 9765 3435 9831 3438
rect 11421 3435 11487 3438
rect 16113 3435 16179 3438
rect 10041 3362 10107 3365
rect 10317 3362 10383 3365
rect 10041 3360 10383 3362
rect 10041 3304 10046 3360
rect 10102 3304 10322 3360
rect 10378 3304 10383 3360
rect 10041 3302 10383 3304
rect 10041 3299 10107 3302
rect 10317 3299 10383 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 9765 3226 9831 3229
rect 11053 3226 11119 3229
rect 9765 3224 11119 3226
rect 9765 3168 9770 3224
rect 9826 3168 11058 3224
rect 11114 3168 11119 3224
rect 9765 3166 11119 3168
rect 9765 3163 9831 3166
rect 11053 3163 11119 3166
rect 0 3090 800 3120
rect 2865 3090 2931 3093
rect 0 3088 2931 3090
rect 0 3032 2870 3088
rect 2926 3032 2931 3088
rect 0 3030 2931 3032
rect 0 3000 800 3030
rect 2865 3027 2931 3030
rect 9673 3090 9739 3093
rect 19057 3090 19123 3093
rect 9673 3088 19123 3090
rect 9673 3032 9678 3088
rect 9734 3032 19062 3088
rect 19118 3032 19123 3088
rect 9673 3030 19123 3032
rect 9673 3027 9739 3030
rect 19057 3027 19123 3030
rect 3693 2818 3759 2821
rect 6269 2818 6335 2821
rect 3693 2816 6335 2818
rect 3693 2760 3698 2816
rect 3754 2760 6274 2816
rect 6330 2760 6335 2816
rect 3693 2758 6335 2760
rect 3693 2755 3759 2758
rect 6269 2755 6335 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 4061 2546 4127 2549
rect 0 2544 4127 2546
rect 0 2488 4066 2544
rect 4122 2488 4127 2544
rect 0 2486 4127 2488
rect 0 2456 800 2486
rect 4061 2483 4127 2486
rect 4409 2208 4729 2209
rect 0 2138 800 2168
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 1485 2138 1551 2141
rect 0 2136 1551 2138
rect 0 2080 1490 2136
rect 1546 2080 1551 2136
rect 0 2078 1551 2080
rect 0 2048 800 2078
rect 1485 2075 1551 2078
rect 0 1594 800 1624
rect 5165 1594 5231 1597
rect 0 1592 5231 1594
rect 0 1536 5170 1592
rect 5226 1536 5231 1592
rect 0 1534 5231 1536
rect 0 1504 800 1534
rect 5165 1531 5231 1534
rect 0 1186 800 1216
rect 1577 1186 1643 1189
rect 0 1184 1643 1186
rect 0 1128 1582 1184
rect 1638 1128 1643 1184
rect 0 1126 1643 1128
rect 0 1096 800 1126
rect 1577 1123 1643 1126
rect 10501 916 10567 917
rect 10501 914 10548 916
rect 10456 912 10548 914
rect 10456 856 10506 912
rect 10456 854 10548 856
rect 10501 852 10548 854
rect 10612 852 10618 916
rect 10501 851 10567 852
rect 0 642 800 672
rect 6361 642 6427 645
rect 0 640 6427 642
rect 0 584 6366 640
rect 6422 584 6427 640
rect 0 582 6427 584
rect 0 552 800 582
rect 6361 579 6427 582
rect 0 234 800 264
rect 3049 234 3115 237
rect 0 232 3115 234
rect 0 176 3054 232
rect 3110 176 3115 232
rect 0 174 3115 176
rect 0 144 800 174
rect 3049 171 3115 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 5764 19136 5828 19140
rect 5764 19080 5778 19136
rect 5778 19080 5828 19136
rect 5764 19076 5828 19080
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 7420 12472 7484 12476
rect 7420 12416 7470 12472
rect 7470 12416 7484 12472
rect 7420 12412 7484 12416
rect 7420 12336 7484 12340
rect 7420 12280 7470 12336
rect 7470 12280 7484 12336
rect 7420 12276 7484 12280
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 5764 9964 5828 10028
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7604 9420 7668 9484
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 10548 8664 10612 8668
rect 10548 8608 10598 8664
rect 10598 8608 10612 8664
rect 10548 8604 10612 8608
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7604 7108 7668 7172
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 7604 5612 7668 5676
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
rect 10548 912 10612 916
rect 10548 856 10562 912
rect 10562 856 10612 912
rect 10548 852 10612 856
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 5763 19140 5829 19141
rect 5763 19076 5764 19140
rect 5828 19076 5829 19140
rect 5763 19075 5829 19076
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 5766 10029 5826 19075
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7419 12476 7485 12477
rect 7419 12412 7420 12476
rect 7484 12412 7485 12476
rect 7419 12411 7485 12412
rect 7422 12341 7482 12411
rect 7419 12340 7485 12341
rect 7419 12276 7420 12340
rect 7484 12276 7485 12340
rect 7419 12275 7485 12276
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 5763 10028 5829 10029
rect 5763 9964 5764 10028
rect 5828 9964 5829 10028
rect 5763 9963 5829 9964
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 7603 9484 7669 9485
rect 7603 9420 7604 9484
rect 7668 9420 7669 9484
rect 7603 9419 7669 9420
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 7606 7173 7666 9419
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 10547 8668 10613 8669
rect 10547 8604 10548 8668
rect 10612 8604 10613 8668
rect 10547 8603 10613 8604
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7603 7172 7669 7173
rect 7603 7108 7604 7172
rect 7668 7108 7669 7172
rect 7603 7107 7669 7108
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 7606 5677 7666 7107
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7603 5676 7669 5677
rect 7603 5612 7604 5676
rect 7668 5612 7669 5676
rect 7603 5611 7669 5612
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 10550 917 10610 8603
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
rect 10547 916 10613 917
rect 10547 852 10548 916
rect 10612 852 10613 916
rect 10547 851 10613 852
use sky130_fd_sc_hd__fill_1  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1608910539
transform 1 0 2208 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 1932 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 2760 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _044_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25
timestamp 1608910539
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_38
timestamp 1608910539
transform 1 0 4600 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1608910539
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4692 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4968 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5520 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1608910539
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1608910539
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608910539
transform 1 0 6348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 6992 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7544 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1608910539
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84
timestamp 1608910539
transform 1 0 8832 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 9936 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10488 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143
timestamp 1608910539
transform 1 0 14260 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1608910539
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13984 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13248 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _088_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608910539
transform 1 0 13524 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608910539
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_146
timestamp 1608910539
transform 1 0 14536 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1608910539
transform 1 0 15088 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608910539
transform 1 0 14904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608910539
transform 1 0 14536 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_156
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1608910539
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608910539
transform 1 0 15548 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608910539
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608910539
transform 1 0 15272 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1608910539
transform 1 0 16284 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1608910539
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1608910539
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608910539
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608910539
transform 1 0 16008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_170
timestamp 1608910539
transform 1 0 16744 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1608910539
transform 1 0 17020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1608910539
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608910539
transform 1 0 16744 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_174
timestamp 1608910539
transform 1 0 17112 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_179
timestamp 1608910539
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_175
timestamp 1608910539
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1608910539
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608910539
transform 1 0 17572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608910539
transform 1 0 17204 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1608910539
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1608910539
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_194
timestamp 1608910539
transform 1 0 18952 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1608910539
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1608910539
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608910539
transform 1 0 19044 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608910539
transform 1 0 18584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_205
timestamp 1608910539
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 1608910539
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1608910539
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1608910539
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608910539
transform 1 0 19412 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_195 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 19044 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1608910539
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_213
timestamp 1608910539
transform 1 0 20700 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1608910539
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1608910539
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1608910539
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608910539
transform 1 0 20332 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 1472 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1656 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1608910539
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4508 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6808 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5980 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8464 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1608910539
transform 1 0 9292 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9844 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10672 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_120
timestamp 1608910539
transform 1 0 12144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_116
timestamp 1608910539
transform 1 0 11776 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12236 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608910539
transform 1 0 11500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 13708 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13892 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_164
timestamp 1608910539
transform 1 0 16192 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1608910539
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1608910539
transform 1 0 14720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1608910539
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15456 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_176
timestamp 1608910539
transform 1 0 17296 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608910539
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_200
timestamp 1608910539
transform 1 0 19504 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_188
timestamp 1608910539
transform 1 0 18400 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1608910539
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1608910539
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1608910539
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1840 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_40
timestamp 1608910539
transform 1 0 4784 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3312 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608910539
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1608910539
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1608910539
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1608910539
transform 1 0 7544 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_92
timestamp 1608910539
transform 1 0 9568 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1608910539
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1608910539
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12512 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_128
timestamp 1608910539
transform 1 0 12880 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13616 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_164
timestamp 1608910539
transform 1 0 16192 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1608910539
transform 1 0 15088 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1608910539
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1608910539
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 17112 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1608910539
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1608910539
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1608910539
transform 1 0 21344 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1608910539
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2024 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1608910539
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4600 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_62
timestamp 1608910539
transform 1 0 6808 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_54
timestamp 1608910539
transform 1 0 6072 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8096 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 7268 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_104
timestamp 1608910539
transform 1 0 10672 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1608910539
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_85
timestamp 1608910539
transform 1 0 8924 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_107
timestamp 1608910539
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1608910539
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1608910539
transform 1 0 14720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 14536 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16100 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_181
timestamp 1608910539
transform 1 0 17756 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16928 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_193
timestamp 1608910539
transform 1 0 18860 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608910539
transform 1 0 19964 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1608910539
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1608910539
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_209
timestamp 1608910539
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1608910539
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1840 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_37
timestamp 1608910539
transform 1 0 4508 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4600 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1608910539
transform 1 0 3680 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_47
timestamp 1608910539
transform 1 0 5428 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 5704 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5888 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_68
timestamp 1608910539
transform 1 0 7360 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7452 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1608910539
transform 1 0 9844 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_87
timestamp 1608910539
transform 1 0 9108 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10304 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_123
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp 1608910539
transform 1 0 12972 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13064 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1608910539
transform 1 0 15364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 14536 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15456 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_186
timestamp 1608910539
transform 1 0 18216 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_201
timestamp 1608910539
transform 1 0 19596 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_194
timestamp 1608910539
transform 1 0 18952 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 19044 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1608910539
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_213
timestamp 1608910539
transform 1 0 20700 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1608910539
transform 1 0 1748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1840 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1748 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_24
timestamp 1608910539
transform 1 0 3312 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1608910539
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1608910539
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3404 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608910539
transform 1 0 3588 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_34
timestamp 1608910539
transform 1 0 4232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_35
timestamp 1608910539
transform 1 0 4324 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4140 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4324 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4692 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_44
timestamp 1608910539
transform 1 0 5152 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_55
timestamp 1608910539
transform 1 0 6164 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5244 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6440 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_79
timestamp 1608910539
transform 1 0 8372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1608910539
transform 1 0 8004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6992 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7912 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8464 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9292 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_7_114
timestamp 1608910539
transform 1 0 11592 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10764 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp 1608910539
transform 1 0 12512 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_118
timestamp 1608910539
transform 1 0 11960 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_7_132
timestamp 1608910539
transform 1 0 13248 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14076 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13800 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1608910539
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 15272 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_163
timestamp 1608910539
transform 1 0 16100 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1608910539
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608910539
transform 1 0 15732 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16376 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16008 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1608910539
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_187
timestamp 1608910539
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608910539
transform 1 0 17480 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1608910539
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1608910539
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_199
timestamp 1608910539
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp 1608910539
transform 1 0 21344 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1608910539
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1608910539
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1608910539
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1608910539
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 2024 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1608910539
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_46
timestamp 1608910539
transform 1 0 5336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6440 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_83
timestamp 1608910539
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 7912 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_87
timestamp 1608910539
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608910539
transform 1 0 10488 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_122
timestamp 1608910539
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_105
timestamp 1608910539
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10856 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_134
timestamp 1608910539
transform 1 0 13432 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13708 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13892 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1608910539
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1608910539
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608910539
transform 1 0 14720 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1608910539
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1608910539
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1608910539
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1608910539
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1608910539
transform 1 0 2300 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1608910539
transform 1 0 4876 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_25
timestamp 1608910539
transform 1 0 3404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608910539
transform 1 0 3128 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1608910539
transform 1 0 5796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 1608910539
transform 1 0 5244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5520 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5888 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_66
timestamp 1608910539
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7452 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608910539
transform 1 0 6900 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_99
timestamp 1608910539
transform 1 0 10212 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_85
timestamp 1608910539
transform 1 0 8924 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 9384 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_114
timestamp 1608910539
transform 1 0 11592 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_141
timestamp 1608910539
transform 1 0 14076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1608910539
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_149
timestamp 1608910539
transform 1 0 14812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15272 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1608910539
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_170
timestamp 1608910539
transform 1 0 16744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1608910539
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1608910539
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 1608910539
transform 1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2852 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1608910539
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4416 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_52
timestamp 1608910539
transform 1 0 5888 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1608910539
transform 1 0 8740 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1608910539
transform 1 0 8188 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6992 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1608910539
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10396 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_117
timestamp 1608910539
transform 1 0 11868 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12604 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14076 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_163
timestamp 1608910539
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_150
timestamp 1608910539
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1608910539
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_175
timestamp 1608910539
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_199
timestamp 1608910539
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1608910539
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1608910539
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1608910539
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_37
timestamp 1608910539
transform 1 0 4508 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4876 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 3496 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608910539
transform 1 0 4600 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1608910539
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7636 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1608910539
transform 1 0 10580 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10304 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9200 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1608910539
transform 1 0 10672 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608910539
transform 1 0 10028 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608910539
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_117
timestamp 1608910539
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1608910539
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1608910539
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_139
timestamp 1608910539
transform 1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12788 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14168 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608910539
transform 1 0 13616 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15640 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1608910539
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_167
timestamp 1608910539
transform 1 0 16468 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1608910539
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1608910539
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 1608910539
transform 1 0 21344 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_17
timestamp 1608910539
transform 1 0 2668 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1608910539
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2760 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4324 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5796 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_69
timestamp 1608910539
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7636 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 12236 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608910539
transform 1 0 11960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1608910539
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1608910539
transform 1 0 12696 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1608910539
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1608910539
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1608910539
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1608910539
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1608910539
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1608910539
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_12
timestamp 1608910539
transform 1 0 2208 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608910539
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1932 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1656 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1608910539
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_40
timestamp 1608910539
transform 1 0 4784 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1608910539
transform 1 0 3588 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4876 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 1608910539
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1608910539
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6348 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608910539
transform 1 0 5520 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1608910539
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7268 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1608910539
transform 1 0 8280 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1608910539
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8096 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10212 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10488 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_110
timestamp 1608910539
transform 1 0 11224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1608910539
transform 1 0 11500 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11500 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1608910539
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_145
timestamp 1608910539
transform 1 0 14444 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13616 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 12972 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1608910539
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608910539
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_157
timestamp 1608910539
transform 1 0 15548 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1608910539
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1608910539
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1608910539
transform 1 0 16652 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1608910539
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1608910539
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1608910539
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1608910539
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1608910539
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 1608910539
transform 1 0 21344 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1748 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1608910539
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_23
timestamp 1608910539
transform 1 0 3220 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4232 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5888 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5060 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1608910539
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8280 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608910539
transform 1 0 7636 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_94
timestamp 1608910539
transform 1 0 9752 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_123
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1608910539
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10856 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608910539
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12696 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13524 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_160
timestamp 1608910539
transform 1 0 15824 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1608910539
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1608910539
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1608910539
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1608910539
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1608910539
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_12
timestamp 1608910539
transform 1 0 2208 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1608910539
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1608910539
transform 1 0 2300 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1608910539
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1608910539
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4692 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608910539
transform 1 0 3128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_57
timestamp 1608910539
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_51
timestamp 1608910539
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6440 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608910539
transform 1 0 5520 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_124
timestamp 1608910539
transform 1 0 12512 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1608910539
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 14260 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1608910539
transform 1 0 13248 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_16_157
timestamp 1608910539
transform 1 0 15548 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1608910539
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_181
timestamp 1608910539
transform 1 0 17756 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_169
timestamp 1608910539
transform 1 0 16652 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1608910539
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1608910539
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1608910539
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1608910539
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_38
timestamp 1608910539
transform 1 0 4600 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_23
timestamp 1608910539
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1608910539
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608910539
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1608910539
transform 1 0 7912 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8004 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 1608910539
transform 1 0 9660 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8832 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1608910539
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_138
timestamp 1608910539
transform 1 0 13800 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_132
timestamp 1608910539
transform 1 0 13248 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14076 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1608910539
transform 1 0 16376 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 14904 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1608910539
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_178
timestamp 1608910539
transform 1 0 17480 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1608910539
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1608910539
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1608910539
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1608910539
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2024 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608910539
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_26
timestamp 1608910539
transform 1 0 3496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4140 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5612 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_74
timestamp 1608910539
transform 1 0 7912 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8648 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1608910539
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 12604 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11132 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_134
timestamp 1608910539
transform 1 0 13432 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 13708 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1608910539
transform 1 0 16284 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1608910539
transform 1 0 17388 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1608910539
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_189
timestamp 1608910539
transform 1 0 18492 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1608910539
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1608910539
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608910539
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_18
timestamp 1608910539
transform 1 0 2760 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2852 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2852 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608910539
transform 1 0 1564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1608910539
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_25
timestamp 1608910539
transform 1 0 3404 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3496 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1608910539
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4508 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5980 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1608910539
transform 1 0 7176 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7268 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8280 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8280 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_20_104
timestamp 1608910539
transform 1 0 10672 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1608910539
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp 1608910539
transform 1 0 11408 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1608910539
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11408 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_20_144
timestamp 1608910539
transform 1 0 14352 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_139
timestamp 1608910539
transform 1 0 13892 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1608910539
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1608910539
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14168 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_20_163
timestamp 1608910539
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1608910539
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 15640 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 16376 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1608910539
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1608910539
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1608910539
transform 1 0 16652 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1608910539
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1608910539
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1608910539
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1608910539
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1608910539
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1608910539
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608910539
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1608910539
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608910539
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608910539
transform 1 0 2576 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_36
timestamp 1608910539
transform 1 0 4416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3312 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608910539
transform 1 0 4140 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1608910539
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 5520 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7084 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7912 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_99
timestamp 1608910539
transform 1 0 10212 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10304 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9384 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_111
timestamp 1608910539
transform 1 0 11316 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1608910539
transform 1 0 12512 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 11868 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1608910539
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12696 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_158
timestamp 1608910539
transform 1 0 15640 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_146
timestamp 1608910539
transform 1 0 14536 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1608910539
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_170
timestamp 1608910539
transform 1 0 16744 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1608910539
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1608910539
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1608910539
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2484 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608910539
transform 1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608910539
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5520 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7176 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8188 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1608910539
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10212 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 9016 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10488 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_115
timestamp 1608910539
transform 1 0 11684 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1608910539
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12236 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1608910539
transform 1 0 13064 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608910539
transform 1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1608910539
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1608910539
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1608910539
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_204
timestamp 1608910539
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_192
timestamp 1608910539
transform 1 0 18768 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1608910539
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1608910539
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608910539
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1608910539
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2576 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_31
timestamp 1608910539
transform 1 0 3956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_51
timestamp 1608910539
transform 1 0 5796 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_43
timestamp 1608910539
transform 1 0 5060 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_81
timestamp 1608910539
transform 1 0 8556 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_77
timestamp 1608910539
transform 1 0 8188 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1608910539
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 7912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608910539
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1608910539
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1608910539
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9844 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12512 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11316 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 13340 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 14352 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_160
timestamp 1608910539
transform 1 0 15824 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1608910539
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_180
timestamp 1608910539
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_172
timestamp 1608910539
transform 1 0 16928 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608910539
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1608910539
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1608910539
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1608910539
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1608910539
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_9
timestamp 1608910539
transform 1 0 1932 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608910539
transform 1 0 2576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1608910539
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608910539
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_50
timestamp 1608910539
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_44
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_83
timestamp 1608910539
transform 1 0 8740 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7268 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1608910539
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_87
timestamp 1608910539
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11224 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12696 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1608910539
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608910539
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1608910539
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1608910539
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1608910539
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1608910539
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608910539
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_17
timestamp 1608910539
transform 1 0 2668 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608910539
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3772 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1608910539
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1608910539
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1608910539
transform 1 0 5244 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 6164 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7912 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_87
timestamp 1608910539
transform 1 0 9108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10212 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1608910539
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_117
timestamp 1608910539
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11040 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_131
timestamp 1608910539
transform 1 0 13156 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13432 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_162
timestamp 1608910539
transform 1 0 16008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_150
timestamp 1608910539
transform 1 0 14904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1608910539
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1608910539
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1608910539
transform 1 0 17112 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608910539
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1608910539
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1608910539
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1608910539
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1932 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608910539
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608910539
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_15
timestamp 1608910539
transform 1 0 2484 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_17
timestamp 1608910539
transform 1 0 2668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2576 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_41
timestamp 1608910539
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1608910539
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1608910539
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4876 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 3404 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608910539
transform 1 0 3588 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1608910539
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1608910539
transform 1 0 6624 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608910539
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6716 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5152 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608910539
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_70
timestamp 1608910539
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8648 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8280 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1608910539
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_84
timestamp 1608910539
transform 1 0 8832 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608910539
transform 1 0 10672 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9752 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608910539
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_125
timestamp 1608910539
transform 1 0 12604 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1608910539
transform 1 0 11776 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10948 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608910539
transform 1 0 11224 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_136
timestamp 1608910539
transform 1 0 13616 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_127
timestamp 1608910539
transform 1 0 12788 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_137
timestamp 1608910539
transform 1 0 13708 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13064 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_160
timestamp 1608910539
transform 1 0 15824 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_148
timestamp 1608910539
transform 1 0 14720 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1608910539
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1608910539
transform 1 0 14812 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1608910539
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1608910539
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_172
timestamp 1608910539
transform 1 0 16928 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1608910539
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608910539
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1608910539
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1608910539
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1608910539
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1608910539
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1608910539
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1608910539
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608910539
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1608910539
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608910539
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2484 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1932 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608910539
transform 1 0 1564 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_21
timestamp 1608910539
transform 1 0 3036 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608910539
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_45
timestamp 1608910539
transform 1 0 5244 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1608910539
transform 1 0 6532 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp 1608910539
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1608910539
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8740 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608910539
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_28_125
timestamp 1608910539
transform 1 0 12604 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11132 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_28_139
timestamp 1608910539
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1608910539
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608910539
transform 1 0 13524 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1608910539
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1608910539
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608910539
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608910539
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1608910539
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1608910539
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1608910539
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1608910539
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608910539
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608910539
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1608910539
transform 1 0 2484 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_5
timestamp 1608910539
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1608910539
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608910539
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2576 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608910539
transform 1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608910539
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4232 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1608910539
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_55
timestamp 1608910539
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608910539
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5060 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608910539
transform 1 0 5888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_82
timestamp 1608910539
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_74
timestamp 1608910539
transform 1 0 7912 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_101
timestamp 1608910539
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1608910539
transform 1 0 9660 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8832 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1608910539
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608910539
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10856 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608910539
transform 1 0 11684 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1608910539
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_163
timestamp 1608910539
transform 1 0 16100 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1608910539
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1608910539
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_175
timestamp 1608910539
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608910539
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1608910539
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1608910539
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_220
timestamp 1608910539
transform 1 0 21344 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608910539
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 1608910539
transform 1 0 2760 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1608910539
transform 1 0 2116 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608910539
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2208 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608910539
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608910539
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_41
timestamp 1608910539
transform 1 0 4876 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1608910539
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_26
timestamp 1608910539
transform 1 0 3496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608910539
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608910539
transform 1 0 3588 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_62
timestamp 1608910539
transform 1 0 6808 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1608910539
transform 1 0 6440 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4968 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1608910539
transform 1 0 8372 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6900 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_30_96
timestamp 1608910539
transform 1 0 9936 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608910539
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 10212 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608910539
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1608910539
transform 1 0 11684 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_105
timestamp 1608910539
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10856 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11776 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1608910539
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14076 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_166
timestamp 1608910539
transform 1 0 16376 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_158
timestamp 1608910539
transform 1 0 15640 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1608910539
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1608910539
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608910539
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1608910539
transform 1 0 18032 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1608910539
transform 1 0 17664 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_175
timestamp 1608910539
transform 1 0 17204 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1608910539
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1608910539
transform 1 0 17848 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 16652 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1608910539
transform 1 0 19228 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_188
timestamp 1608910539
transform 1 0 18400 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1608910539
transform 1 0 18492 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 18676 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1608910539
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1608910539
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1608910539
transform 1 0 20332 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608910539
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608910539
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1608910539
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608910539
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1840 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2392 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608910539
transform 1 0 1472 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4692 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3220 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1608910539
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608910539
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8464 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6992 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_103
timestamp 1608910539
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_86
timestamp 1608910539
transform 1 0 9016 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9108 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1608910539
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608910539
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10764 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1608910539
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 12972 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608910539
transform 1 0 14444 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608910539
transform 1 0 13892 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608910539
transform 1 0 13524 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1608910539
transform 1 0 15548 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 16376 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608910539
transform 1 0 16008 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608910539
transform 1 0 15640 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608910539
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608910539
transform 1 0 14812 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1608910539
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608910539
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1608910539
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608910539
transform 1 0 17480 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_204
timestamp 1608910539
transform 1 0 19872 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1608910539
transform 1 0 19504 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1608910539
transform 1 0 19136 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1608910539
transform 1 0 18768 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1608910539
transform 1 0 18400 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1608910539
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_216
timestamp 1608910539
transform 1 0 20976 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608910539
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_18
timestamp 1608910539
transform 1 0 2760 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp 1608910539
transform 1 0 2116 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608910539
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2208 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608910539
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608910539
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_41
timestamp 1608910539
transform 1 0 4876 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1608910539
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_24
timestamp 1608910539
transform 1 0 3312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608910539
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608910539
transform 1 0 3588 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6440 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4968 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7268 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8096 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_32_104
timestamp 1608910539
transform 1 0 10672 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608910539
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1608910539
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1608910539
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10948 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608910539
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1608910539
transform 1 0 14076 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_134
timestamp 1608910539
transform 1 0 13432 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1608910539
transform 1 0 12972 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1608910539
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1608910539
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1608910539
transform 1 0 13064 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1608910539
transform 1 0 13524 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1608910539
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_154
timestamp 1608910539
transform 1 0 15272 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1608910539
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1608910539
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1608910539
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608910539
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1608910539
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608910539
transform 1 0 16284 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_187
timestamp 1608910539
transform 1 0 18308 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_175
timestamp 1608910539
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1608910539
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1608910539
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1608910539
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_196
timestamp 1608910539
transform 1 0 19136 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_192
timestamp 1608910539
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1608910539
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1608910539
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1608910539
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608910539
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608910539
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1608910539
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1608910539
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1608910539
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608910539
transform 1 0 2116 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608910539
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_40
timestamp 1608910539
transform 1 0 4784 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_32
timestamp 1608910539
transform 1 0 4048 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1608910539
transform 1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4876 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608910539
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_60
timestamp 1608910539
transform 1 0 6624 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_43
timestamp 1608910539
transform 1 0 5060 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1608910539
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5612 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_33_78
timestamp 1608910539
transform 1 0 8280 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_75
timestamp 1608910539
transform 1 0 8004 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1608910539
transform 1 0 7636 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_67
timestamp 1608910539
transform 1 0 7268 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_63
timestamp 1608910539
transform 1 0 6900 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608910539
transform 1 0 7360 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1608910539
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_90
timestamp 1608910539
transform 1 0 9384 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1608910539
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1608910539
transform 1 0 12604 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_118
timestamp 1608910539
transform 1 0 11960 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_106
timestamp 1608910539
transform 1 0 10856 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1608910539
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1608910539
transform 1 0 13708 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_156
timestamp 1608910539
transform 1 0 15456 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_149
timestamp 1608910539
transform 1 0 14812 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1608910539
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_187
timestamp 1608910539
transform 1 0 18308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1608910539
transform 1 0 17664 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_168
timestamp 1608910539
transform 1 0 16560 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1608910539
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_199
timestamp 1608910539
transform 1 0 19412 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1608910539
transform 1 0 21528 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1608910539
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_211
timestamp 1608910539
transform 1 0 20516 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1608910539
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1608910539
transform -1 0 21896 0 1 20128
box -38 -48 314 592
<< labels >>
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 0 nsew signal input
rlabel metal2 s 662 0 718 800 6 bottom_left_grid_pin_43_
port 1 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 bottom_left_grid_pin_44_
port 2 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 bottom_left_grid_pin_45_
port 3 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_46_
port 4 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 bottom_left_grid_pin_47_
port 5 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 bottom_left_grid_pin_48_
port 6 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 bottom_left_grid_pin_49_
port 7 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 bottom_right_grid_pin_1_
port 8 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 9 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 10 nsew signal tristate
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[0]
port 11 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[10]
port 12 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[11]
port 13 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[12]
port 14 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[13]
port 15 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[14]
port 16 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 17 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[16]
port 18 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[17]
port 19 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[18]
port 20 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[19]
port 21 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 22 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[2]
port 23 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[3]
port 24 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 chanx_left_in[4]
port 25 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[5]
port 26 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[6]
port 27 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[7]
port 28 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[8]
port 29 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[9]
port 30 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[0]
port 31 nsew signal tristate
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[10]
port 32 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 33 nsew signal tristate
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[12]
port 34 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 35 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[14]
port 36 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 37 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[16]
port 38 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 39 nsew signal tristate
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[18]
port 40 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 41 nsew signal tristate
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[1]
port 42 nsew signal tristate
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[2]
port 43 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 44 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[4]
port 45 nsew signal tristate
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[5]
port 46 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[6]
port 47 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[7]
port 48 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[8]
port 49 nsew signal tristate
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[9]
port 50 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[0]
port 51 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[10]
port 52 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[11]
port 53 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 54 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[13]
port 55 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[14]
port 56 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[15]
port 57 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[16]
port 58 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[17]
port 59 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[18]
port 60 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[19]
port 61 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[1]
port 62 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_in[2]
port 63 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[3]
port 64 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[4]
port 65 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[5]
port 66 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[6]
port 67 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[7]
port 68 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[8]
port 69 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 70 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[0]
port 71 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 chany_bottom_out[10]
port 72 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_out[11]
port 73 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[12]
port 74 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[13]
port 75 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[14]
port 76 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 chany_bottom_out[15]
port 77 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[16]
port 78 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 chany_bottom_out[17]
port 79 nsew signal tristate
rlabel metal2 s 21730 0 21786 800 6 chany_bottom_out[18]
port 80 nsew signal tristate
rlabel metal2 s 22190 0 22246 800 6 chany_bottom_out[19]
port 81 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[1]
port 82 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[2]
port 83 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[3]
port 84 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[4]
port 85 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[5]
port 86 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_out[6]
port 87 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[7]
port 88 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[8]
port 89 nsew signal tristate
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[9]
port 90 nsew signal tristate
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 91 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 92 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 93 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 94 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 95 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 96 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 97 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 98 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 99 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 100 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 101 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 102 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 103 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 104 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 105 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 106 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 107 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 108 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 109 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 110 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 111 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 112 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 113 nsew signal tristate
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 114 nsew signal tristate
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 115 nsew signal tristate
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 116 nsew signal tristate
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 117 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 118 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 119 nsew signal tristate
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 120 nsew signal tristate
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 121 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 122 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 123 nsew signal tristate
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 124 nsew signal tristate
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 125 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 126 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 127 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 128 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 129 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 130 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 131 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 132 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 left_bottom_grid_pin_36_
port 133 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 134 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_38_
port 135 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 136 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_40_
port 137 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 138 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 139 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 140 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 141 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 142 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 143 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 144 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 145 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 146 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 147 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 148 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 149 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 150 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 151 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 152 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 153 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
