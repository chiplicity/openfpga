VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__1_
  CLASS BLOCK ;
  FOREIGN sb_2__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN bottom_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END bottom_left_grid_pin_34_
  PIN bottom_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 2.400 ;
    END
  END bottom_left_grid_pin_35_
  PIN bottom_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END bottom_left_grid_pin_36_
  PIN bottom_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END bottom_left_grid_pin_37_
  PIN bottom_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END bottom_left_grid_pin_38_
  PIN bottom_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 2.400 ;
    END
  END bottom_left_grid_pin_39_
  PIN bottom_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END bottom_left_grid_pin_40_
  PIN bottom_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END bottom_left_grid_pin_41_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.400 ;
    END
  END bottom_right_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 116.320 140.000 116.920 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 2.400 10.160 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 2.400 27.840 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 2.400 89.040 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.400 92.440 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 2.400 95.160 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 2.400 97.880 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 2.400 104.000 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 2.400 72.040 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 2.400 74.760 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 2.400 83.600 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 2.400 86.320 ;
    END
  END chanx_left_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 137.600 52.810 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 137.600 55.570 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 137.600 58.790 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 137.600 61.550 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 137.600 64.310 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 137.600 67.070 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 137.600 73.050 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 137.600 75.810 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 137.600 78.570 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 137.600 27.050 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 137.600 30.270 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 137.600 33.030 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 137.600 35.790 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 137.600 41.310 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 137.600 44.530 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 137.600 47.290 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 137.600 50.050 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 137.600 81.330 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 137.600 109.850 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 137.600 112.610 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 137.600 115.830 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 137.600 118.590 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 137.600 121.350 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 137.600 124.110 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 137.600 130.090 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 137.600 132.850 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 137.600 84.090 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 137.600 90.070 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 137.600 92.830 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 137.600 95.590 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 137.600 98.350 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 137.600 101.570 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 137.600 104.330 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 137.600 107.090 140.000 ;
    END
  END chany_top_out[9]
  PIN left_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.400 118.280 ;
    END
  END left_top_grid_pin_42_
  PIN left_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 2.400 121.000 ;
    END
  END left_top_grid_pin_43_
  PIN left_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 2.400 124.400 ;
    END
  END left_top_grid_pin_44_
  PIN left_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_top_grid_pin_45_
  PIN left_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END left_top_grid_pin_46_
  PIN left_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.400 133.240 ;
    END
  END left_top_grid_pin_47_
  PIN left_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END left_top_grid_pin_48_
  PIN left_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 2.400 138.680 ;
    END
  END left_top_grid_pin_49_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.160 140.000 23.760 ;
    END
  END prog_clk
  PIN top_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_34_
  PIN top_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 137.600 4.510 140.000 ;
    END
  END top_left_grid_pin_35_
  PIN top_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 137.600 7.270 140.000 ;
    END
  END top_left_grid_pin_36_
  PIN top_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 137.600 10.030 140.000 ;
    END
  END top_left_grid_pin_37_
  PIN top_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 137.600 12.790 140.000 ;
    END
  END top_left_grid_pin_38_
  PIN top_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 137.600 16.010 140.000 ;
    END
  END top_left_grid_pin_39_
  PIN top_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 137.600 18.770 140.000 ;
    END
  END top_left_grid_pin_40_
  PIN top_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 137.600 21.530 140.000 ;
    END
  END top_left_grid_pin_41_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 137.600 138.370 140.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 4.210 8.540 138.390 128.080 ;
      LAYER met2 ;
        RECT 0.090 137.320 1.190 138.565 ;
        RECT 2.030 137.320 3.950 138.565 ;
        RECT 4.790 137.320 6.710 138.565 ;
        RECT 7.550 137.320 9.470 138.565 ;
        RECT 10.310 137.320 12.230 138.565 ;
        RECT 13.070 137.320 15.450 138.565 ;
        RECT 16.290 137.320 18.210 138.565 ;
        RECT 19.050 137.320 20.970 138.565 ;
        RECT 21.810 137.320 23.730 138.565 ;
        RECT 24.570 137.320 26.490 138.565 ;
        RECT 27.330 137.320 29.710 138.565 ;
        RECT 30.550 137.320 32.470 138.565 ;
        RECT 33.310 137.320 35.230 138.565 ;
        RECT 36.070 137.320 37.990 138.565 ;
        RECT 38.830 137.320 40.750 138.565 ;
        RECT 41.590 137.320 43.970 138.565 ;
        RECT 44.810 137.320 46.730 138.565 ;
        RECT 47.570 137.320 49.490 138.565 ;
        RECT 50.330 137.320 52.250 138.565 ;
        RECT 53.090 137.320 55.010 138.565 ;
        RECT 55.850 137.320 58.230 138.565 ;
        RECT 59.070 137.320 60.990 138.565 ;
        RECT 61.830 137.320 63.750 138.565 ;
        RECT 64.590 137.320 66.510 138.565 ;
        RECT 67.350 137.320 69.270 138.565 ;
        RECT 70.110 137.320 72.490 138.565 ;
        RECT 73.330 137.320 75.250 138.565 ;
        RECT 76.090 137.320 78.010 138.565 ;
        RECT 78.850 137.320 80.770 138.565 ;
        RECT 81.610 137.320 83.530 138.565 ;
        RECT 84.370 137.320 86.750 138.565 ;
        RECT 87.590 137.320 89.510 138.565 ;
        RECT 90.350 137.320 92.270 138.565 ;
        RECT 93.110 137.320 95.030 138.565 ;
        RECT 95.870 137.320 97.790 138.565 ;
        RECT 98.630 137.320 101.010 138.565 ;
        RECT 101.850 137.320 103.770 138.565 ;
        RECT 104.610 137.320 106.530 138.565 ;
        RECT 107.370 137.320 109.290 138.565 ;
        RECT 110.130 137.320 112.050 138.565 ;
        RECT 112.890 137.320 115.270 138.565 ;
        RECT 116.110 137.320 118.030 138.565 ;
        RECT 118.870 137.320 120.790 138.565 ;
        RECT 121.630 137.320 123.550 138.565 ;
        RECT 124.390 137.320 126.310 138.565 ;
        RECT 127.150 137.320 129.530 138.565 ;
        RECT 130.370 137.320 132.290 138.565 ;
        RECT 133.130 137.320 135.050 138.565 ;
        RECT 135.890 137.320 137.810 138.565 ;
        RECT 0.090 2.680 138.370 137.320 ;
        RECT 0.090 0.155 1.190 2.680 ;
        RECT 2.030 0.155 3.950 2.680 ;
        RECT 4.790 0.155 6.710 2.680 ;
        RECT 7.550 0.155 9.470 2.680 ;
        RECT 10.310 0.155 12.230 2.680 ;
        RECT 13.070 0.155 15.450 2.680 ;
        RECT 16.290 0.155 18.210 2.680 ;
        RECT 19.050 0.155 20.970 2.680 ;
        RECT 21.810 0.155 23.730 2.680 ;
        RECT 24.570 0.155 26.490 2.680 ;
        RECT 27.330 0.155 29.710 2.680 ;
        RECT 30.550 0.155 32.470 2.680 ;
        RECT 33.310 0.155 35.230 2.680 ;
        RECT 36.070 0.155 37.990 2.680 ;
        RECT 38.830 0.155 40.750 2.680 ;
        RECT 41.590 0.155 43.970 2.680 ;
        RECT 44.810 0.155 46.730 2.680 ;
        RECT 47.570 0.155 49.490 2.680 ;
        RECT 50.330 0.155 52.250 2.680 ;
        RECT 53.090 0.155 55.010 2.680 ;
        RECT 55.850 0.155 58.230 2.680 ;
        RECT 59.070 0.155 60.990 2.680 ;
        RECT 61.830 0.155 63.750 2.680 ;
        RECT 64.590 0.155 66.510 2.680 ;
        RECT 67.350 0.155 69.270 2.680 ;
        RECT 70.110 0.155 72.490 2.680 ;
        RECT 73.330 0.155 75.250 2.680 ;
        RECT 76.090 0.155 78.010 2.680 ;
        RECT 78.850 0.155 80.770 2.680 ;
        RECT 81.610 0.155 83.530 2.680 ;
        RECT 84.370 0.155 86.750 2.680 ;
        RECT 87.590 0.155 89.510 2.680 ;
        RECT 90.350 0.155 92.270 2.680 ;
        RECT 93.110 0.155 95.030 2.680 ;
        RECT 95.870 0.155 97.790 2.680 ;
        RECT 98.630 0.155 101.010 2.680 ;
        RECT 101.850 0.155 103.770 2.680 ;
        RECT 104.610 0.155 106.530 2.680 ;
        RECT 107.370 0.155 109.290 2.680 ;
        RECT 110.130 0.155 112.050 2.680 ;
        RECT 112.890 0.155 115.270 2.680 ;
        RECT 116.110 0.155 118.030 2.680 ;
        RECT 118.870 0.155 120.790 2.680 ;
        RECT 121.630 0.155 123.550 2.680 ;
        RECT 124.390 0.155 126.310 2.680 ;
        RECT 127.150 0.155 129.530 2.680 ;
        RECT 130.370 0.155 132.290 2.680 ;
        RECT 133.130 0.155 135.050 2.680 ;
        RECT 135.890 0.155 137.810 2.680 ;
      LAYER met3 ;
        RECT 2.800 137.680 138.395 138.545 ;
        RECT 0.065 136.360 138.395 137.680 ;
        RECT 2.800 134.960 138.395 136.360 ;
        RECT 0.065 133.640 138.395 134.960 ;
        RECT 2.800 132.240 138.395 133.640 ;
        RECT 0.065 130.240 138.395 132.240 ;
        RECT 2.800 128.840 138.395 130.240 ;
        RECT 0.065 127.520 138.395 128.840 ;
        RECT 2.800 126.120 138.395 127.520 ;
        RECT 0.065 124.800 138.395 126.120 ;
        RECT 2.800 123.400 138.395 124.800 ;
        RECT 0.065 121.400 138.395 123.400 ;
        RECT 2.800 120.000 138.395 121.400 ;
        RECT 0.065 118.680 138.395 120.000 ;
        RECT 2.800 117.320 138.395 118.680 ;
        RECT 2.800 117.280 137.200 117.320 ;
        RECT 0.065 115.960 137.200 117.280 ;
        RECT 2.800 115.920 137.200 115.960 ;
        RECT 2.800 114.560 138.395 115.920 ;
        RECT 0.065 113.240 138.395 114.560 ;
        RECT 2.800 111.840 138.395 113.240 ;
        RECT 0.065 109.840 138.395 111.840 ;
        RECT 2.800 108.440 138.395 109.840 ;
        RECT 0.065 107.120 138.395 108.440 ;
        RECT 2.800 105.720 138.395 107.120 ;
        RECT 0.065 104.400 138.395 105.720 ;
        RECT 2.800 103.000 138.395 104.400 ;
        RECT 0.065 101.000 138.395 103.000 ;
        RECT 2.800 99.600 138.395 101.000 ;
        RECT 0.065 98.280 138.395 99.600 ;
        RECT 2.800 96.880 138.395 98.280 ;
        RECT 0.065 95.560 138.395 96.880 ;
        RECT 2.800 94.160 138.395 95.560 ;
        RECT 0.065 92.840 138.395 94.160 ;
        RECT 2.800 91.440 138.395 92.840 ;
        RECT 0.065 89.440 138.395 91.440 ;
        RECT 2.800 88.040 138.395 89.440 ;
        RECT 0.065 86.720 138.395 88.040 ;
        RECT 2.800 85.320 138.395 86.720 ;
        RECT 0.065 84.000 138.395 85.320 ;
        RECT 2.800 82.600 138.395 84.000 ;
        RECT 0.065 80.600 138.395 82.600 ;
        RECT 2.800 79.200 138.395 80.600 ;
        RECT 0.065 77.880 138.395 79.200 ;
        RECT 2.800 76.480 138.395 77.880 ;
        RECT 0.065 75.160 138.395 76.480 ;
        RECT 2.800 73.760 138.395 75.160 ;
        RECT 0.065 72.440 138.395 73.760 ;
        RECT 2.800 71.040 138.395 72.440 ;
        RECT 0.065 70.400 138.395 71.040 ;
        RECT 0.065 69.040 137.200 70.400 ;
        RECT 2.800 69.000 137.200 69.040 ;
        RECT 2.800 67.640 138.395 69.000 ;
        RECT 0.065 66.320 138.395 67.640 ;
        RECT 2.800 64.920 138.395 66.320 ;
        RECT 0.065 63.600 138.395 64.920 ;
        RECT 2.800 62.200 138.395 63.600 ;
        RECT 0.065 60.200 138.395 62.200 ;
        RECT 2.800 58.800 138.395 60.200 ;
        RECT 0.065 57.480 138.395 58.800 ;
        RECT 2.800 56.080 138.395 57.480 ;
        RECT 0.065 54.760 138.395 56.080 ;
        RECT 2.800 53.360 138.395 54.760 ;
        RECT 0.065 51.360 138.395 53.360 ;
        RECT 2.800 49.960 138.395 51.360 ;
        RECT 0.065 48.640 138.395 49.960 ;
        RECT 2.800 47.240 138.395 48.640 ;
        RECT 0.065 45.920 138.395 47.240 ;
        RECT 2.800 44.520 138.395 45.920 ;
        RECT 0.065 43.200 138.395 44.520 ;
        RECT 2.800 41.800 138.395 43.200 ;
        RECT 0.065 39.800 138.395 41.800 ;
        RECT 2.800 38.400 138.395 39.800 ;
        RECT 0.065 37.080 138.395 38.400 ;
        RECT 2.800 35.680 138.395 37.080 ;
        RECT 0.065 34.360 138.395 35.680 ;
        RECT 2.800 32.960 138.395 34.360 ;
        RECT 0.065 30.960 138.395 32.960 ;
        RECT 2.800 29.560 138.395 30.960 ;
        RECT 0.065 28.240 138.395 29.560 ;
        RECT 2.800 26.840 138.395 28.240 ;
        RECT 0.065 25.520 138.395 26.840 ;
        RECT 2.800 24.160 138.395 25.520 ;
        RECT 2.800 24.120 137.200 24.160 ;
        RECT 0.065 22.800 137.200 24.120 ;
        RECT 2.800 22.760 137.200 22.800 ;
        RECT 2.800 21.400 138.395 22.760 ;
        RECT 0.065 19.400 138.395 21.400 ;
        RECT 2.800 18.000 138.395 19.400 ;
        RECT 0.065 16.680 138.395 18.000 ;
        RECT 2.800 15.280 138.395 16.680 ;
        RECT 0.065 13.960 138.395 15.280 ;
        RECT 2.800 12.560 138.395 13.960 ;
        RECT 0.065 10.560 138.395 12.560 ;
        RECT 2.800 9.160 138.395 10.560 ;
        RECT 0.065 7.840 138.395 9.160 ;
        RECT 2.800 6.440 138.395 7.840 ;
        RECT 0.065 5.120 138.395 6.440 ;
        RECT 2.800 3.720 138.395 5.120 ;
        RECT 0.065 2.400 138.395 3.720 ;
        RECT 2.800 1.000 138.395 2.400 ;
        RECT 0.065 0.175 138.395 1.000 ;
      LAYER met4 ;
        RECT 8.150 10.240 27.655 128.080 ;
        RECT 30.055 10.240 50.985 128.080 ;
        RECT 53.385 10.240 132.610 128.080 ;
        RECT 8.150 5.615 132.610 10.240 ;
      LAYER met5 ;
        RECT 7.940 11.100 132.820 60.300 ;
  END
END sb_2__1_
END LIBRARY

